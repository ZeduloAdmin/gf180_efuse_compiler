* eFuse array netlist with word_width=1, nwords=16

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
X0 ZN I VSS VPW nfet_06v0 W=8.2e-07 L=6e-07  
X1 ZN I VDD VNW pfet_06v0 W=1.22e-06 L=5e-07
.ENDS

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
X00 ZN I VSS VPW nfet_06v0 W=8.2e-07 L=6e-07
X01 VSS I ZN VPW nfet_06v0 W=8.2e-07 L=6e-07
X10 ZN I VDD VNW pfet_06v0 W=1.22e-06 L=5e-07
X11 VDD I ZN VNW pfet_06v0 W=1.22e-06 L=5e-07
.ENDS

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
X17 net_1 net_0 VSS VPW nfet_06v0 W=8.2e-07 L=1e-06
X19 VDD net_1 net_0 VNW pfet_06v0 W=1.22e-06 L=1e-06
.ENDS

.subckt efuse_bitcell VSS VDD SELECT ANODE PARAMS: NUM=-1
X0 ANODE CATHODE efuse NUM={NUM}
X1 CATHODE SELECT VSS VSS nfet_06v0 L=0.60u W=30.5u
.ends

.subckt efuse_senseamp VSS VNW VDD PRESET_N OUT SENSE FUSE
X2 net1 PRESET_N VDD VDD pfet_06v0 L=0.5u W=2.44u nf=2
X1 net2 OUT VDD VDD VSS VNW gf180mcu_fd_sc_mcu7t5v0__inv_1
X2 net1 net2 VDD VDD VSS VNW gf180mcu_fd_sc_mcu7t5v0__inv_1
X3 net2 net1 VDD VDD VSS VNW gf180mcu_fd_sc_mcu7t5v0__inv_1
X1 net1 SENSE FUSE VSS nfet_06v0 L=0.60u W=0.82u
.ends


.subckt efuse_bitline VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] COL_PROG_N OUT PARAMS: LNUM=0
X0 VSS VDD BIT_SEL[0] bitline efuse_bitcell NUM={LNUM*1000+0}
X1 VSS VDD BIT_SEL[1] bitline efuse_bitcell NUM={LNUM*1000+1}
X2 VSS VDD BIT_SEL[2] bitline efuse_bitcell NUM={LNUM*1000+2}
X3 VSS VDD BIT_SEL[3] bitline efuse_bitcell NUM={LNUM*1000+3}
X4 VSS VDD BIT_SEL[4] bitline efuse_bitcell NUM={LNUM*1000+4}
X5 VSS VDD BIT_SEL[5] bitline efuse_bitcell NUM={LNUM*1000+5}
X6 VSS VDD BIT_SEL[6] bitline efuse_bitcell NUM={LNUM*1000+6}
X7 VSS VDD BIT_SEL[7] bitline efuse_bitcell NUM={LNUM*1000+7}
X8 VSS VDD BIT_SEL[8] bitline efuse_bitcell NUM={LNUM*1000+8}
X9 VSS VDD BIT_SEL[9] bitline efuse_bitcell NUM={LNUM*1000+9}
X10 VSS VDD BIT_SEL[10] bitline efuse_bitcell NUM={LNUM*1000+10}
X11 VSS VDD BIT_SEL[11] bitline efuse_bitcell NUM={LNUM*1000+11}
X12 VSS VDD BIT_SEL[12] bitline efuse_bitcell NUM={LNUM*1000+12}
X13 VSS VDD BIT_SEL[13] bitline efuse_bitcell NUM={LNUM*1000+13}
X14 VSS VDD BIT_SEL[14] bitline efuse_bitcell NUM={LNUM*1000+14}
X15 VSS VDD BIT_SEL[15] bitline efuse_bitcell NUM={LNUM*1000+15}
X0 bitline COL_PROG_N VDD VDD pfet_06v0 L=0.50u W=76.5u nf=1
X1 bitline COL_PROG_N VDD VDD pfet_06v0 L=0.50u W=76.5u nf=1
Xsense VSS VSS VDD PRESET_N OUT SENSE bitline efuse_senseamp
.ends
    

.subckt efuse_array_16x1 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] COL_PROG_N[0] OUT[0]  
X0 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15]   COL_PROG_N[0] OUT[0]  efuse_bitline LNUM=0

.ends
    
.end
    