* eFuse array netlist with word_width=8, nwords=32
    
.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
X0 ZN I VSS VPW nfet_06v0 W=8.2e-07 L=6e-07  
X1 ZN I VDD VNW pfet_06v0 W=1.22e-06 L=5e-07
.ENDS

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
X00 ZN I VSS VPW nfet_06v0 W=8.2e-07 L=6e-07
X01 VSS I ZN VPW nfet_06v0 W=8.2e-07 L=6e-07
X10 ZN I VDD VNW pfet_06v0 W=1.22e-06 L=5e-07
X11 VDD I ZN VNW pfet_06v0 W=1.22e-06 L=5e-07
.ENDS

.subckt efuse_bitcell VSS SELECT ANODE
X0 ANODE CATHODE efuse
X1 CATHODE SELECT VSS VSS nfet_06v0 L=0.60u W=30.5u
.ends

.subckt efuse_senseamp  VDD PRESET_N OUT SENSE VSS FUSE
X2 net1 PRESET_N VDD VDD pfet_06v0 L=0.5u W=2.44u nf=2
x1 net2 OUT VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x2 net1 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x3 net2 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X1 net1 SENSE FUSE VSS nfet_06v0 L=0.60u W=0.82u
.ends


.subckt efuse_bitline VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] COL_PROG_N OUT
X0 VSS BIT_SEL[0] bitline efuse_bitcell
X1 VSS BIT_SEL[1] bitline efuse_bitcell
X2 VSS BIT_SEL[2] bitline efuse_bitcell
X3 VSS BIT_SEL[3] bitline efuse_bitcell
X4 VSS BIT_SEL[4] bitline efuse_bitcell
X5 VSS BIT_SEL[5] bitline efuse_bitcell
X6 VSS BIT_SEL[6] bitline efuse_bitcell
X7 VSS BIT_SEL[7] bitline efuse_bitcell
X8 VSS BIT_SEL[8] bitline efuse_bitcell
X9 VSS BIT_SEL[9] bitline efuse_bitcell
X10 VSS BIT_SEL[10] bitline efuse_bitcell
X11 VSS BIT_SEL[11] bitline efuse_bitcell
X12 VSS BIT_SEL[12] bitline efuse_bitcell
X13 VSS BIT_SEL[13] bitline efuse_bitcell
X14 VSS BIT_SEL[14] bitline efuse_bitcell
X15 VSS BIT_SEL[15] bitline efuse_bitcell
X16 VSS BIT_SEL[16] bitline efuse_bitcell
X17 VSS BIT_SEL[17] bitline efuse_bitcell
X18 VSS BIT_SEL[18] bitline efuse_bitcell
X19 VSS BIT_SEL[19] bitline efuse_bitcell
X20 VSS BIT_SEL[20] bitline efuse_bitcell
X21 VSS BIT_SEL[21] bitline efuse_bitcell
X22 VSS BIT_SEL[22] bitline efuse_bitcell
X23 VSS BIT_SEL[23] bitline efuse_bitcell
X24 VSS BIT_SEL[24] bitline efuse_bitcell
X25 VSS BIT_SEL[25] bitline efuse_bitcell
X26 VSS BIT_SEL[26] bitline efuse_bitcell
X27 VSS BIT_SEL[27] bitline efuse_bitcell
X28 VSS BIT_SEL[28] bitline efuse_bitcell
X29 VSS BIT_SEL[29] bitline efuse_bitcell
X30 VSS BIT_SEL[30] bitline efuse_bitcell
X31 VSS BIT_SEL[31] bitline efuse_bitcell
X0 bitline COL_PROG_N VDD VDD pfet_06v0 L=0.50u W=76.5u nf=2
X1 bitline COL_PROG_N VDD VDD pfet_06v0 L=0.50u W=76.5u nf=2
Xsense VDD PRESET_N OUT SENSE VSS bitline efuse_senseamp
.ends
    

.subckt efuse_array_32x8 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] COL_PROG_N[0] OUT[0] COL_PROG_N[1] OUT[1] COL_PROG_N[2] OUT[2] COL_PROG_N[3] OUT[3] COL_PROG_N[4] OUT[4] COL_PROG_N[5] OUT[5] COL_PROG_N[6] OUT[6] COL_PROG_N[7] OUT[7] 
X0_0 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31]  COL_PROG_N[0] OUT[0]  efuse_bitline
X0_1 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31]  COL_PROG_N[1] OUT[1]  efuse_bitline
X0_2 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31]  COL_PROG_N[2] OUT[2]  efuse_bitline
X0_3 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31]  COL_PROG_N[3] OUT[3]  efuse_bitline
X0_4 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31]  COL_PROG_N[4] OUT[4]  efuse_bitline
X0_5 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31]  COL_PROG_N[5] OUT[5]  efuse_bitline
X0_6 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31]  COL_PROG_N[6] OUT[6]  efuse_bitline
X0_7 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31]  COL_PROG_N[7] OUT[7]  efuse_bitline

.ends
    
.end
    