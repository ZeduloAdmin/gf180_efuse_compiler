VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_array_64x8
  CLASS BLOCK ;
  FOREIGN efuse_array_64x8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 141.830 BY 315.825 ;
  PIN COL_PROG_N[0]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 136.790 39.430 140.350 39.730 ;
    END
  END COL_PROG_N[0]
  PIN COL_PROG_N[1]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 136.790 78.815 140.350 79.115 ;
    END
  END COL_PROG_N[1]
  PIN COL_PROG_N[2]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 136.790 118.200 140.350 118.500 ;
    END
  END COL_PROG_N[2]
  PIN COL_PROG_N[3]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 136.790 157.585 140.350 157.885 ;
    END
  END COL_PROG_N[3]
  PIN COL_PROG_N[4]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 136.790 196.970 140.350 197.270 ;
    END
  END COL_PROG_N[4]
  PIN COL_PROG_N[5]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 136.790 236.355 140.350 236.655 ;
    END
  END COL_PROG_N[5]
  PIN COL_PROG_N[6]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 136.790 275.740 140.350 276.040 ;
    END
  END COL_PROG_N[6]
  PIN COL_PROG_N[7]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 136.790 315.125 140.350 315.425 ;
    END
  END COL_PROG_N[7]
  PIN PRESET_N
    ANTENNAGATEAREA 9.760000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.010 295.580 1.290 315.825 ;
        RECT 1.010 295.200 1.370 295.580 ;
        RECT 1.010 256.195 1.290 295.200 ;
        RECT 1.010 255.815 1.370 256.195 ;
        RECT 1.010 216.810 1.290 255.815 ;
        RECT 1.010 216.430 1.370 216.810 ;
        RECT 1.010 177.425 1.290 216.430 ;
        RECT 1.010 177.045 1.370 177.425 ;
        RECT 1.010 138.040 1.290 177.045 ;
        RECT 1.010 137.660 1.370 138.040 ;
        RECT 1.010 98.655 1.290 137.660 ;
        RECT 1.010 98.275 1.370 98.655 ;
        RECT 1.010 59.270 1.290 98.275 ;
        RECT 1.010 58.890 1.370 59.270 ;
        RECT 1.010 19.885 1.290 58.890 ;
        RECT 1.010 19.505 1.370 19.885 ;
        RECT 1.010 0.000 1.290 19.505 ;
    END
  END PRESET_N
  PIN SENSE
    ANTENNAGATEAREA 3.936000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.655 294.395 1.935 315.825 ;
        RECT 1.655 294.015 3.080 294.395 ;
        RECT 1.655 255.010 1.935 294.015 ;
        RECT 1.655 254.630 3.080 255.010 ;
        RECT 1.655 215.625 1.935 254.630 ;
        RECT 1.655 215.245 3.080 215.625 ;
        RECT 1.655 176.240 1.935 215.245 ;
        RECT 1.655 175.860 3.080 176.240 ;
        RECT 1.655 136.855 1.935 175.860 ;
        RECT 1.655 136.475 3.080 136.855 ;
        RECT 1.655 97.470 1.935 136.475 ;
        RECT 1.655 97.090 3.080 97.470 ;
        RECT 1.655 58.085 1.935 97.090 ;
        RECT 1.655 57.705 3.080 58.085 ;
        RECT 1.655 18.700 1.935 57.705 ;
        RECT 1.655 18.320 3.080 18.700 ;
        RECT 1.655 0.000 1.935 18.320 ;
    END
  END SENSE
  PIN OUT[0]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 11.030 2.680 11.410 ;
    END
  END OUT[0]
  PIN OUT[1]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 50.415 2.680 50.795 ;
    END
  END OUT[1]
  PIN OUT[2]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 89.800 2.680 90.180 ;
    END
  END OUT[2]
  PIN OUT[3]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 129.185 2.680 129.565 ;
    END
  END OUT[3]
  PIN OUT[4]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 168.570 2.680 168.950 ;
    END
  END OUT[4]
  PIN OUT[5]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 207.955 2.680 208.335 ;
    END
  END OUT[5]
  PIN OUT[6]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 247.340 2.680 247.720 ;
    END
  END OUT[6]
  PIN OUT[7]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 286.725 2.680 287.105 ;
    END
  END OUT[7]
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 104.050 0.000 106.910 315.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.600 0.000 74.460 315.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 39.150 0.000 42.010 315.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3.710 0.000 4.710 315.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 6.700 0.000 9.560 315.825 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 137.340 0.000 141.590 315.825 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.070 0.000 1.070 315.825 ;
    END
  END VDD
  PIN BIT_SEL[48]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 135.090 299.920 135.370 315.200 ;
        RECT 135.050 299.540 135.430 299.920 ;
        RECT 135.090 260.535 135.370 299.540 ;
        RECT 135.050 260.155 135.430 260.535 ;
        RECT 135.090 221.150 135.370 260.155 ;
        RECT 135.050 220.770 135.430 221.150 ;
        RECT 135.090 181.765 135.370 220.770 ;
        RECT 135.050 181.385 135.430 181.765 ;
        RECT 135.090 142.380 135.370 181.385 ;
        RECT 135.050 142.000 135.430 142.380 ;
        RECT 135.090 102.995 135.370 142.000 ;
        RECT 135.050 102.615 135.430 102.995 ;
        RECT 135.090 63.610 135.370 102.615 ;
        RECT 135.050 63.230 135.430 63.610 ;
        RECT 135.090 24.225 135.370 63.230 ;
        RECT 135.050 23.845 135.430 24.225 ;
        RECT 135.090 0.000 135.370 23.845 ;
    END
  END BIT_SEL[48]
  PIN BIT_SEL[49]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 134.450 291.355 134.730 315.200 ;
        RECT 134.410 290.975 134.790 291.355 ;
        RECT 134.450 251.970 134.730 290.975 ;
        RECT 134.410 251.590 134.790 251.970 ;
        RECT 134.450 212.585 134.730 251.590 ;
        RECT 134.410 212.205 134.790 212.585 ;
        RECT 134.450 173.200 134.730 212.205 ;
        RECT 134.410 172.820 134.790 173.200 ;
        RECT 134.450 133.815 134.730 172.820 ;
        RECT 134.410 133.435 134.790 133.815 ;
        RECT 134.450 94.430 134.730 133.435 ;
        RECT 134.410 94.050 134.790 94.430 ;
        RECT 134.450 55.045 134.730 94.050 ;
        RECT 134.410 54.665 134.790 55.045 ;
        RECT 134.450 15.660 134.730 54.665 ;
        RECT 134.410 15.280 134.790 15.660 ;
        RECT 134.450 0.000 134.730 15.280 ;
    END
  END BIT_SEL[49]
  PIN BIT_SEL[50]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 133.810 301.760 134.090 315.200 ;
        RECT 133.770 301.380 134.150 301.760 ;
        RECT 133.810 262.375 134.090 301.380 ;
        RECT 133.770 261.995 134.150 262.375 ;
        RECT 133.810 222.990 134.090 261.995 ;
        RECT 133.770 222.610 134.150 222.990 ;
        RECT 133.810 183.605 134.090 222.610 ;
        RECT 133.770 183.225 134.150 183.605 ;
        RECT 133.810 144.220 134.090 183.225 ;
        RECT 133.770 143.840 134.150 144.220 ;
        RECT 133.810 104.835 134.090 143.840 ;
        RECT 133.770 104.455 134.150 104.835 ;
        RECT 133.810 65.450 134.090 104.455 ;
        RECT 133.770 65.070 134.150 65.450 ;
        RECT 133.810 26.065 134.090 65.070 ;
        RECT 133.770 25.685 134.150 26.065 ;
        RECT 133.810 0.000 134.090 25.685 ;
    END
  END BIT_SEL[50]
  PIN BIT_SEL[51]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 133.170 289.515 133.450 315.200 ;
        RECT 133.130 289.135 133.510 289.515 ;
        RECT 133.170 250.130 133.450 289.135 ;
        RECT 133.130 249.750 133.510 250.130 ;
        RECT 133.170 210.745 133.450 249.750 ;
        RECT 133.130 210.365 133.510 210.745 ;
        RECT 133.170 171.360 133.450 210.365 ;
        RECT 133.130 170.980 133.510 171.360 ;
        RECT 133.170 131.975 133.450 170.980 ;
        RECT 133.130 131.595 133.510 131.975 ;
        RECT 133.170 92.590 133.450 131.595 ;
        RECT 133.130 92.210 133.510 92.590 ;
        RECT 133.170 53.205 133.450 92.210 ;
        RECT 133.130 52.825 133.510 53.205 ;
        RECT 133.170 13.820 133.450 52.825 ;
        RECT 133.130 13.440 133.510 13.820 ;
        RECT 133.170 0.000 133.450 13.440 ;
    END
  END BIT_SEL[51]
  PIN BIT_SEL[52]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 132.530 303.600 132.810 315.200 ;
        RECT 132.490 303.220 132.870 303.600 ;
        RECT 132.530 264.215 132.810 303.220 ;
        RECT 132.490 263.835 132.870 264.215 ;
        RECT 132.530 224.830 132.810 263.835 ;
        RECT 132.490 224.450 132.870 224.830 ;
        RECT 132.530 185.445 132.810 224.450 ;
        RECT 132.490 185.065 132.870 185.445 ;
        RECT 132.530 146.060 132.810 185.065 ;
        RECT 132.490 145.680 132.870 146.060 ;
        RECT 132.530 106.675 132.810 145.680 ;
        RECT 132.490 106.295 132.870 106.675 ;
        RECT 132.530 67.290 132.810 106.295 ;
        RECT 132.490 66.910 132.870 67.290 ;
        RECT 132.530 27.905 132.810 66.910 ;
        RECT 132.490 27.525 132.870 27.905 ;
        RECT 132.530 0.000 132.810 27.525 ;
    END
  END BIT_SEL[52]
  PIN BIT_SEL[53]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 131.890 287.670 132.170 315.200 ;
        RECT 131.850 287.290 132.230 287.670 ;
        RECT 131.890 248.285 132.170 287.290 ;
        RECT 131.850 247.905 132.230 248.285 ;
        RECT 131.890 208.900 132.170 247.905 ;
        RECT 131.850 208.520 132.230 208.900 ;
        RECT 131.890 169.515 132.170 208.520 ;
        RECT 131.850 169.135 132.230 169.515 ;
        RECT 131.890 130.130 132.170 169.135 ;
        RECT 131.850 129.750 132.230 130.130 ;
        RECT 131.890 90.745 132.170 129.750 ;
        RECT 131.850 90.365 132.230 90.745 ;
        RECT 131.890 51.360 132.170 90.365 ;
        RECT 131.850 50.980 132.230 51.360 ;
        RECT 131.890 11.975 132.170 50.980 ;
        RECT 131.850 11.595 132.230 11.975 ;
        RECT 131.890 0.000 132.170 11.595 ;
    END
  END BIT_SEL[53]
  PIN BIT_SEL[54]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 131.250 306.245 131.530 315.200 ;
        RECT 131.210 305.865 131.590 306.245 ;
        RECT 131.250 266.860 131.530 305.865 ;
        RECT 131.210 266.480 131.590 266.860 ;
        RECT 131.250 227.475 131.530 266.480 ;
        RECT 131.210 227.095 131.590 227.475 ;
        RECT 131.250 188.090 131.530 227.095 ;
        RECT 131.210 187.710 131.590 188.090 ;
        RECT 131.250 148.705 131.530 187.710 ;
        RECT 131.210 148.325 131.590 148.705 ;
        RECT 131.250 109.320 131.530 148.325 ;
        RECT 131.210 108.940 131.590 109.320 ;
        RECT 131.250 69.935 131.530 108.940 ;
        RECT 131.210 69.555 131.590 69.935 ;
        RECT 131.250 30.550 131.530 69.555 ;
        RECT 131.210 30.170 131.590 30.550 ;
        RECT 131.250 0.000 131.530 30.170 ;
    END
  END BIT_SEL[54]
  PIN BIT_SEL[55]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 130.610 285.030 130.890 315.200 ;
        RECT 130.570 284.650 130.950 285.030 ;
        RECT 130.610 245.645 130.890 284.650 ;
        RECT 130.570 245.265 130.950 245.645 ;
        RECT 130.610 206.260 130.890 245.265 ;
        RECT 130.570 205.880 130.950 206.260 ;
        RECT 130.610 166.875 130.890 205.880 ;
        RECT 130.570 166.495 130.950 166.875 ;
        RECT 130.610 127.490 130.890 166.495 ;
        RECT 130.570 127.110 130.950 127.490 ;
        RECT 130.610 88.105 130.890 127.110 ;
        RECT 130.570 87.725 130.950 88.105 ;
        RECT 130.610 48.720 130.890 87.725 ;
        RECT 130.570 48.340 130.950 48.720 ;
        RECT 130.610 9.335 130.890 48.340 ;
        RECT 130.570 8.955 130.950 9.335 ;
        RECT 130.610 0.000 130.890 8.955 ;
    END
  END BIT_SEL[55]
  PIN BIT_SEL[56]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 129.970 308.085 130.250 315.200 ;
        RECT 129.930 307.705 130.310 308.085 ;
        RECT 129.970 268.700 130.250 307.705 ;
        RECT 129.930 268.320 130.310 268.700 ;
        RECT 129.970 229.315 130.250 268.320 ;
        RECT 129.930 228.935 130.310 229.315 ;
        RECT 129.970 189.930 130.250 228.935 ;
        RECT 129.930 189.550 130.310 189.930 ;
        RECT 129.970 150.545 130.250 189.550 ;
        RECT 129.930 150.165 130.310 150.545 ;
        RECT 129.970 111.160 130.250 150.165 ;
        RECT 129.930 110.780 130.310 111.160 ;
        RECT 129.970 71.775 130.250 110.780 ;
        RECT 129.930 71.395 130.310 71.775 ;
        RECT 129.970 32.390 130.250 71.395 ;
        RECT 129.930 32.010 130.310 32.390 ;
        RECT 129.970 0.000 130.250 32.010 ;
    END
  END BIT_SEL[56]
  PIN BIT_SEL[57]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 129.330 283.190 129.610 315.200 ;
        RECT 129.290 282.810 129.670 283.190 ;
        RECT 129.330 243.805 129.610 282.810 ;
        RECT 129.290 243.425 129.670 243.805 ;
        RECT 129.330 204.420 129.610 243.425 ;
        RECT 129.290 204.040 129.670 204.420 ;
        RECT 129.330 165.035 129.610 204.040 ;
        RECT 129.290 164.655 129.670 165.035 ;
        RECT 129.330 125.650 129.610 164.655 ;
        RECT 129.290 125.270 129.670 125.650 ;
        RECT 129.330 86.265 129.610 125.270 ;
        RECT 129.290 85.885 129.670 86.265 ;
        RECT 129.330 46.880 129.610 85.885 ;
        RECT 129.290 46.500 129.670 46.880 ;
        RECT 129.330 7.495 129.610 46.500 ;
        RECT 129.290 7.115 129.670 7.495 ;
        RECT 129.330 0.000 129.610 7.115 ;
    END
  END BIT_SEL[57]
  PIN BIT_SEL[58]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 128.690 309.925 128.970 315.200 ;
        RECT 128.650 309.545 129.030 309.925 ;
        RECT 128.690 270.540 128.970 309.545 ;
        RECT 128.650 270.160 129.030 270.540 ;
        RECT 128.690 231.155 128.970 270.160 ;
        RECT 128.650 230.775 129.030 231.155 ;
        RECT 128.690 191.770 128.970 230.775 ;
        RECT 128.650 191.390 129.030 191.770 ;
        RECT 128.690 152.385 128.970 191.390 ;
        RECT 128.650 152.005 129.030 152.385 ;
        RECT 128.690 113.000 128.970 152.005 ;
        RECT 128.650 112.620 129.030 113.000 ;
        RECT 128.690 73.615 128.970 112.620 ;
        RECT 128.650 73.235 129.030 73.615 ;
        RECT 128.690 34.230 128.970 73.235 ;
        RECT 128.650 33.850 129.030 34.230 ;
        RECT 128.690 0.000 128.970 33.850 ;
    END
  END BIT_SEL[58]
  PIN BIT_SEL[59]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 128.050 281.345 128.330 315.200 ;
        RECT 128.010 280.965 128.390 281.345 ;
        RECT 128.050 241.960 128.330 280.965 ;
        RECT 128.010 241.580 128.390 241.960 ;
        RECT 128.050 202.575 128.330 241.580 ;
        RECT 128.010 202.195 128.390 202.575 ;
        RECT 128.050 163.190 128.330 202.195 ;
        RECT 128.010 162.810 128.390 163.190 ;
        RECT 128.050 123.805 128.330 162.810 ;
        RECT 128.010 123.425 128.390 123.805 ;
        RECT 128.050 84.420 128.330 123.425 ;
        RECT 128.010 84.040 128.390 84.420 ;
        RECT 128.050 45.035 128.330 84.040 ;
        RECT 128.010 44.655 128.390 45.035 ;
        RECT 128.050 5.650 128.330 44.655 ;
        RECT 128.010 5.270 128.390 5.650 ;
        RECT 128.050 0.000 128.330 5.270 ;
    END
  END BIT_SEL[59]
  PIN BIT_SEL[60]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 127.410 312.570 127.690 315.200 ;
        RECT 127.370 312.190 127.750 312.570 ;
        RECT 127.410 273.185 127.690 312.190 ;
        RECT 127.370 272.805 127.750 273.185 ;
        RECT 127.410 233.800 127.690 272.805 ;
        RECT 127.370 233.420 127.750 233.800 ;
        RECT 127.410 194.415 127.690 233.420 ;
        RECT 127.370 194.035 127.750 194.415 ;
        RECT 127.410 155.030 127.690 194.035 ;
        RECT 127.370 154.650 127.750 155.030 ;
        RECT 127.410 115.645 127.690 154.650 ;
        RECT 127.370 115.265 127.750 115.645 ;
        RECT 127.410 76.260 127.690 115.265 ;
        RECT 127.370 75.880 127.750 76.260 ;
        RECT 127.410 36.875 127.690 75.880 ;
        RECT 127.370 36.495 127.750 36.875 ;
        RECT 127.410 0.000 127.690 36.495 ;
    END
  END BIT_SEL[60]
  PIN BIT_SEL[61]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 126.770 278.705 127.050 315.200 ;
        RECT 126.730 278.325 127.110 278.705 ;
        RECT 126.770 239.320 127.050 278.325 ;
        RECT 126.730 238.940 127.110 239.320 ;
        RECT 126.770 199.935 127.050 238.940 ;
        RECT 126.730 199.555 127.110 199.935 ;
        RECT 126.770 160.550 127.050 199.555 ;
        RECT 126.730 160.170 127.110 160.550 ;
        RECT 126.770 121.165 127.050 160.170 ;
        RECT 126.730 120.785 127.110 121.165 ;
        RECT 126.770 81.780 127.050 120.785 ;
        RECT 126.730 81.400 127.110 81.780 ;
        RECT 126.770 42.395 127.050 81.400 ;
        RECT 126.730 42.015 127.110 42.395 ;
        RECT 126.770 3.010 127.050 42.015 ;
        RECT 126.730 2.630 127.110 3.010 ;
        RECT 126.770 0.000 127.050 2.630 ;
    END
  END BIT_SEL[61]
  PIN BIT_SEL[62]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 126.130 314.410 126.410 315.200 ;
        RECT 126.090 314.030 126.470 314.410 ;
        RECT 126.130 275.025 126.410 314.030 ;
        RECT 126.090 274.645 126.470 275.025 ;
        RECT 126.130 235.640 126.410 274.645 ;
        RECT 126.090 235.260 126.470 235.640 ;
        RECT 126.130 196.255 126.410 235.260 ;
        RECT 126.090 195.875 126.470 196.255 ;
        RECT 126.130 156.870 126.410 195.875 ;
        RECT 126.090 156.490 126.470 156.870 ;
        RECT 126.130 117.485 126.410 156.490 ;
        RECT 126.090 117.105 126.470 117.485 ;
        RECT 126.130 78.100 126.410 117.105 ;
        RECT 126.090 77.720 126.470 78.100 ;
        RECT 126.130 38.715 126.410 77.720 ;
        RECT 126.090 38.335 126.470 38.715 ;
        RECT 126.130 0.000 126.410 38.335 ;
    END
  END BIT_SEL[62]
  PIN BIT_SEL[63]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 125.490 276.865 125.770 315.200 ;
        RECT 125.450 276.485 125.830 276.865 ;
        RECT 125.490 237.480 125.770 276.485 ;
        RECT 125.450 237.100 125.830 237.480 ;
        RECT 125.490 198.095 125.770 237.100 ;
        RECT 125.450 197.715 125.830 198.095 ;
        RECT 125.490 158.710 125.770 197.715 ;
        RECT 125.450 158.330 125.830 158.710 ;
        RECT 125.490 119.325 125.770 158.330 ;
        RECT 125.450 118.945 125.830 119.325 ;
        RECT 125.490 79.940 125.770 118.945 ;
        RECT 125.450 79.560 125.830 79.940 ;
        RECT 125.490 40.555 125.770 79.560 ;
        RECT 125.450 40.175 125.830 40.555 ;
        RECT 125.490 1.170 125.770 40.175 ;
        RECT 125.450 0.790 125.830 1.170 ;
        RECT 125.490 0.000 125.770 0.790 ;
    END
  END BIT_SEL[63]
  PIN BIT_SEL[46]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 93.680 314.410 93.960 315.200 ;
        RECT 93.640 314.030 94.020 314.410 ;
        RECT 93.680 275.025 93.960 314.030 ;
        RECT 93.640 274.645 94.020 275.025 ;
        RECT 93.680 235.640 93.960 274.645 ;
        RECT 93.640 235.260 94.020 235.640 ;
        RECT 93.680 196.255 93.960 235.260 ;
        RECT 93.640 195.875 94.020 196.255 ;
        RECT 93.680 156.870 93.960 195.875 ;
        RECT 93.640 156.490 94.020 156.870 ;
        RECT 93.680 117.485 93.960 156.490 ;
        RECT 93.640 117.105 94.020 117.485 ;
        RECT 93.680 78.100 93.960 117.105 ;
        RECT 93.640 77.720 94.020 78.100 ;
        RECT 93.680 38.715 93.960 77.720 ;
        RECT 93.640 38.335 94.020 38.715 ;
        RECT 93.680 0.000 93.960 38.335 ;
    END
  END BIT_SEL[46]
  PIN BIT_SEL[47]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 93.040 276.865 93.320 315.200 ;
        RECT 93.000 276.485 93.380 276.865 ;
        RECT 93.040 237.480 93.320 276.485 ;
        RECT 93.000 237.100 93.380 237.480 ;
        RECT 93.040 198.095 93.320 237.100 ;
        RECT 93.000 197.715 93.380 198.095 ;
        RECT 93.040 158.710 93.320 197.715 ;
        RECT 93.000 158.330 93.380 158.710 ;
        RECT 93.040 119.325 93.320 158.330 ;
        RECT 93.000 118.945 93.380 119.325 ;
        RECT 93.040 79.940 93.320 118.945 ;
        RECT 93.000 79.560 93.380 79.940 ;
        RECT 93.040 40.555 93.320 79.560 ;
        RECT 93.000 40.175 93.380 40.555 ;
        RECT 93.040 1.170 93.320 40.175 ;
        RECT 93.000 0.790 93.380 1.170 ;
        RECT 93.040 0.000 93.320 0.790 ;
    END
  END BIT_SEL[47]
  PIN BIT_SEL[16]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 70.190 299.920 70.470 315.200 ;
        RECT 70.150 299.540 70.530 299.920 ;
        RECT 70.190 260.535 70.470 299.540 ;
        RECT 70.150 260.155 70.530 260.535 ;
        RECT 70.190 221.150 70.470 260.155 ;
        RECT 70.150 220.770 70.530 221.150 ;
        RECT 70.190 181.765 70.470 220.770 ;
        RECT 70.150 181.385 70.530 181.765 ;
        RECT 70.190 142.380 70.470 181.385 ;
        RECT 70.150 142.000 70.530 142.380 ;
        RECT 70.190 102.995 70.470 142.000 ;
        RECT 70.150 102.615 70.530 102.995 ;
        RECT 70.190 63.610 70.470 102.615 ;
        RECT 70.150 63.230 70.530 63.610 ;
        RECT 70.190 24.225 70.470 63.230 ;
        RECT 70.150 23.845 70.530 24.225 ;
        RECT 70.190 0.000 70.470 23.845 ;
    END
  END BIT_SEL[16]
  PIN BIT_SEL[32]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 102.640 299.920 102.920 315.200 ;
        RECT 102.600 299.540 102.980 299.920 ;
        RECT 102.640 260.535 102.920 299.540 ;
        RECT 102.600 260.155 102.980 260.535 ;
        RECT 102.640 221.150 102.920 260.155 ;
        RECT 102.600 220.770 102.980 221.150 ;
        RECT 102.640 181.765 102.920 220.770 ;
        RECT 102.600 181.385 102.980 181.765 ;
        RECT 102.640 142.380 102.920 181.385 ;
        RECT 102.600 142.000 102.980 142.380 ;
        RECT 102.640 102.995 102.920 142.000 ;
        RECT 102.600 102.615 102.980 102.995 ;
        RECT 102.640 63.610 102.920 102.615 ;
        RECT 102.600 63.230 102.980 63.610 ;
        RECT 102.640 24.225 102.920 63.230 ;
        RECT 102.600 23.845 102.980 24.225 ;
        RECT 102.640 0.000 102.920 23.845 ;
    END
  END BIT_SEL[32]
  PIN BIT_SEL[33]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 102.000 291.355 102.280 315.200 ;
        RECT 101.960 290.975 102.340 291.355 ;
        RECT 102.000 251.970 102.280 290.975 ;
        RECT 101.960 251.590 102.340 251.970 ;
        RECT 102.000 212.585 102.280 251.590 ;
        RECT 101.960 212.205 102.340 212.585 ;
        RECT 102.000 173.200 102.280 212.205 ;
        RECT 101.960 172.820 102.340 173.200 ;
        RECT 102.000 133.815 102.280 172.820 ;
        RECT 101.960 133.435 102.340 133.815 ;
        RECT 102.000 94.430 102.280 133.435 ;
        RECT 101.960 94.050 102.340 94.430 ;
        RECT 102.000 55.045 102.280 94.050 ;
        RECT 101.960 54.665 102.340 55.045 ;
        RECT 102.000 15.660 102.280 54.665 ;
        RECT 101.960 15.280 102.340 15.660 ;
        RECT 102.000 0.000 102.280 15.280 ;
    END
  END BIT_SEL[33]
  PIN BIT_SEL[34]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 101.360 301.760 101.640 315.200 ;
        RECT 101.320 301.380 101.700 301.760 ;
        RECT 101.360 262.375 101.640 301.380 ;
        RECT 101.320 261.995 101.700 262.375 ;
        RECT 101.360 222.990 101.640 261.995 ;
        RECT 101.320 222.610 101.700 222.990 ;
        RECT 101.360 183.605 101.640 222.610 ;
        RECT 101.320 183.225 101.700 183.605 ;
        RECT 101.360 144.220 101.640 183.225 ;
        RECT 101.320 143.840 101.700 144.220 ;
        RECT 101.360 104.835 101.640 143.840 ;
        RECT 101.320 104.455 101.700 104.835 ;
        RECT 101.360 65.450 101.640 104.455 ;
        RECT 101.320 65.070 101.700 65.450 ;
        RECT 101.360 26.065 101.640 65.070 ;
        RECT 101.320 25.685 101.700 26.065 ;
        RECT 101.360 0.000 101.640 25.685 ;
    END
  END BIT_SEL[34]
  PIN BIT_SEL[35]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 100.720 289.515 101.000 315.200 ;
        RECT 100.680 289.135 101.060 289.515 ;
        RECT 100.720 250.130 101.000 289.135 ;
        RECT 100.680 249.750 101.060 250.130 ;
        RECT 100.720 210.745 101.000 249.750 ;
        RECT 100.680 210.365 101.060 210.745 ;
        RECT 100.720 171.360 101.000 210.365 ;
        RECT 100.680 170.980 101.060 171.360 ;
        RECT 100.720 131.975 101.000 170.980 ;
        RECT 100.680 131.595 101.060 131.975 ;
        RECT 100.720 92.590 101.000 131.595 ;
        RECT 100.680 92.210 101.060 92.590 ;
        RECT 100.720 53.205 101.000 92.210 ;
        RECT 100.680 52.825 101.060 53.205 ;
        RECT 100.720 13.820 101.000 52.825 ;
        RECT 100.680 13.440 101.060 13.820 ;
        RECT 100.720 0.000 101.000 13.440 ;
    END
  END BIT_SEL[35]
  PIN BIT_SEL[36]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 100.080 303.600 100.360 315.200 ;
        RECT 100.040 303.220 100.420 303.600 ;
        RECT 100.080 264.215 100.360 303.220 ;
        RECT 100.040 263.835 100.420 264.215 ;
        RECT 100.080 224.830 100.360 263.835 ;
        RECT 100.040 224.450 100.420 224.830 ;
        RECT 100.080 185.445 100.360 224.450 ;
        RECT 100.040 185.065 100.420 185.445 ;
        RECT 100.080 146.060 100.360 185.065 ;
        RECT 100.040 145.680 100.420 146.060 ;
        RECT 100.080 106.675 100.360 145.680 ;
        RECT 100.040 106.295 100.420 106.675 ;
        RECT 100.080 67.290 100.360 106.295 ;
        RECT 100.040 66.910 100.420 67.290 ;
        RECT 100.080 27.905 100.360 66.910 ;
        RECT 100.040 27.525 100.420 27.905 ;
        RECT 100.080 0.000 100.360 27.525 ;
    END
  END BIT_SEL[36]
  PIN BIT_SEL[37]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 99.440 287.670 99.720 315.200 ;
        RECT 99.400 287.290 99.780 287.670 ;
        RECT 99.440 248.285 99.720 287.290 ;
        RECT 99.400 247.905 99.780 248.285 ;
        RECT 99.440 208.900 99.720 247.905 ;
        RECT 99.400 208.520 99.780 208.900 ;
        RECT 99.440 169.515 99.720 208.520 ;
        RECT 99.400 169.135 99.780 169.515 ;
        RECT 99.440 130.130 99.720 169.135 ;
        RECT 99.400 129.750 99.780 130.130 ;
        RECT 99.440 90.745 99.720 129.750 ;
        RECT 99.400 90.365 99.780 90.745 ;
        RECT 99.440 51.360 99.720 90.365 ;
        RECT 99.400 50.980 99.780 51.360 ;
        RECT 99.440 11.975 99.720 50.980 ;
        RECT 99.400 11.595 99.780 11.975 ;
        RECT 99.440 0.000 99.720 11.595 ;
    END
  END BIT_SEL[37]
  PIN BIT_SEL[38]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 98.800 306.245 99.080 315.200 ;
        RECT 98.760 305.865 99.140 306.245 ;
        RECT 98.800 266.860 99.080 305.865 ;
        RECT 98.760 266.480 99.140 266.860 ;
        RECT 98.800 227.475 99.080 266.480 ;
        RECT 98.760 227.095 99.140 227.475 ;
        RECT 98.800 188.090 99.080 227.095 ;
        RECT 98.760 187.710 99.140 188.090 ;
        RECT 98.800 148.705 99.080 187.710 ;
        RECT 98.760 148.325 99.140 148.705 ;
        RECT 98.800 109.320 99.080 148.325 ;
        RECT 98.760 108.940 99.140 109.320 ;
        RECT 98.800 69.935 99.080 108.940 ;
        RECT 98.760 69.555 99.140 69.935 ;
        RECT 98.800 30.550 99.080 69.555 ;
        RECT 98.760 30.170 99.140 30.550 ;
        RECT 98.800 0.000 99.080 30.170 ;
    END
  END BIT_SEL[38]
  PIN BIT_SEL[39]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 98.160 285.030 98.440 315.200 ;
        RECT 98.120 284.650 98.500 285.030 ;
        RECT 98.160 245.645 98.440 284.650 ;
        RECT 98.120 245.265 98.500 245.645 ;
        RECT 98.160 206.260 98.440 245.265 ;
        RECT 98.120 205.880 98.500 206.260 ;
        RECT 98.160 166.875 98.440 205.880 ;
        RECT 98.120 166.495 98.500 166.875 ;
        RECT 98.160 127.490 98.440 166.495 ;
        RECT 98.120 127.110 98.500 127.490 ;
        RECT 98.160 88.105 98.440 127.110 ;
        RECT 98.120 87.725 98.500 88.105 ;
        RECT 98.160 48.720 98.440 87.725 ;
        RECT 98.120 48.340 98.500 48.720 ;
        RECT 98.160 9.335 98.440 48.340 ;
        RECT 98.120 8.955 98.500 9.335 ;
        RECT 98.160 0.000 98.440 8.955 ;
    END
  END BIT_SEL[39]
  PIN BIT_SEL[40]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 97.520 308.085 97.800 315.200 ;
        RECT 97.480 307.705 97.860 308.085 ;
        RECT 97.520 268.700 97.800 307.705 ;
        RECT 97.480 268.320 97.860 268.700 ;
        RECT 97.520 229.315 97.800 268.320 ;
        RECT 97.480 228.935 97.860 229.315 ;
        RECT 97.520 189.930 97.800 228.935 ;
        RECT 97.480 189.550 97.860 189.930 ;
        RECT 97.520 150.545 97.800 189.550 ;
        RECT 97.480 150.165 97.860 150.545 ;
        RECT 97.520 111.160 97.800 150.165 ;
        RECT 97.480 110.780 97.860 111.160 ;
        RECT 97.520 71.775 97.800 110.780 ;
        RECT 97.480 71.395 97.860 71.775 ;
        RECT 97.520 32.390 97.800 71.395 ;
        RECT 97.480 32.010 97.860 32.390 ;
        RECT 97.520 0.000 97.800 32.010 ;
    END
  END BIT_SEL[40]
  PIN BIT_SEL[41]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 96.880 283.190 97.160 315.200 ;
        RECT 96.840 282.810 97.220 283.190 ;
        RECT 96.880 243.805 97.160 282.810 ;
        RECT 96.840 243.425 97.220 243.805 ;
        RECT 96.880 204.420 97.160 243.425 ;
        RECT 96.840 204.040 97.220 204.420 ;
        RECT 96.880 165.035 97.160 204.040 ;
        RECT 96.840 164.655 97.220 165.035 ;
        RECT 96.880 125.650 97.160 164.655 ;
        RECT 96.840 125.270 97.220 125.650 ;
        RECT 96.880 86.265 97.160 125.270 ;
        RECT 96.840 85.885 97.220 86.265 ;
        RECT 96.880 46.880 97.160 85.885 ;
        RECT 96.840 46.500 97.220 46.880 ;
        RECT 96.880 7.495 97.160 46.500 ;
        RECT 96.840 7.115 97.220 7.495 ;
        RECT 96.880 0.000 97.160 7.115 ;
    END
  END BIT_SEL[41]
  PIN BIT_SEL[42]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 96.240 309.925 96.520 315.200 ;
        RECT 96.200 309.545 96.580 309.925 ;
        RECT 96.240 270.540 96.520 309.545 ;
        RECT 96.200 270.160 96.580 270.540 ;
        RECT 96.240 231.155 96.520 270.160 ;
        RECT 96.200 230.775 96.580 231.155 ;
        RECT 96.240 191.770 96.520 230.775 ;
        RECT 96.200 191.390 96.580 191.770 ;
        RECT 96.240 152.385 96.520 191.390 ;
        RECT 96.200 152.005 96.580 152.385 ;
        RECT 96.240 113.000 96.520 152.005 ;
        RECT 96.200 112.620 96.580 113.000 ;
        RECT 96.240 73.615 96.520 112.620 ;
        RECT 96.200 73.235 96.580 73.615 ;
        RECT 96.240 34.230 96.520 73.235 ;
        RECT 96.200 33.850 96.580 34.230 ;
        RECT 96.240 0.000 96.520 33.850 ;
    END
  END BIT_SEL[42]
  PIN BIT_SEL[43]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 95.600 281.345 95.880 315.200 ;
        RECT 95.560 280.965 95.940 281.345 ;
        RECT 95.600 241.960 95.880 280.965 ;
        RECT 95.560 241.580 95.940 241.960 ;
        RECT 95.600 202.575 95.880 241.580 ;
        RECT 95.560 202.195 95.940 202.575 ;
        RECT 95.600 163.190 95.880 202.195 ;
        RECT 95.560 162.810 95.940 163.190 ;
        RECT 95.600 123.805 95.880 162.810 ;
        RECT 95.560 123.425 95.940 123.805 ;
        RECT 95.600 84.420 95.880 123.425 ;
        RECT 95.560 84.040 95.940 84.420 ;
        RECT 95.600 45.035 95.880 84.040 ;
        RECT 95.560 44.655 95.940 45.035 ;
        RECT 95.600 5.650 95.880 44.655 ;
        RECT 95.560 5.270 95.940 5.650 ;
        RECT 95.600 0.000 95.880 5.270 ;
    END
  END BIT_SEL[43]
  PIN BIT_SEL[44]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 94.960 312.570 95.240 315.200 ;
        RECT 94.920 312.190 95.300 312.570 ;
        RECT 94.960 273.185 95.240 312.190 ;
        RECT 94.920 272.805 95.300 273.185 ;
        RECT 94.960 233.800 95.240 272.805 ;
        RECT 94.920 233.420 95.300 233.800 ;
        RECT 94.960 194.415 95.240 233.420 ;
        RECT 94.920 194.035 95.300 194.415 ;
        RECT 94.960 155.030 95.240 194.035 ;
        RECT 94.920 154.650 95.300 155.030 ;
        RECT 94.960 115.645 95.240 154.650 ;
        RECT 94.920 115.265 95.300 115.645 ;
        RECT 94.960 76.260 95.240 115.265 ;
        RECT 94.920 75.880 95.300 76.260 ;
        RECT 94.960 36.875 95.240 75.880 ;
        RECT 94.920 36.495 95.300 36.875 ;
        RECT 94.960 0.000 95.240 36.495 ;
    END
  END BIT_SEL[44]
  PIN BIT_SEL[45]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 94.320 278.705 94.600 315.200 ;
        RECT 94.280 278.325 94.660 278.705 ;
        RECT 94.320 239.320 94.600 278.325 ;
        RECT 94.280 238.940 94.660 239.320 ;
        RECT 94.320 199.935 94.600 238.940 ;
        RECT 94.280 199.555 94.660 199.935 ;
        RECT 94.320 160.550 94.600 199.555 ;
        RECT 94.280 160.170 94.660 160.550 ;
        RECT 94.320 121.165 94.600 160.170 ;
        RECT 94.280 120.785 94.660 121.165 ;
        RECT 94.320 81.780 94.600 120.785 ;
        RECT 94.280 81.400 94.660 81.780 ;
        RECT 94.320 42.395 94.600 81.400 ;
        RECT 94.280 42.015 94.660 42.395 ;
        RECT 94.320 3.010 94.600 42.015 ;
        RECT 94.280 2.630 94.660 3.010 ;
        RECT 94.320 0.000 94.600 2.630 ;
    END
  END BIT_SEL[45]
  PIN BIT_SEL[0]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 37.740 299.920 38.020 315.200 ;
        RECT 37.700 299.540 38.080 299.920 ;
        RECT 37.740 260.535 38.020 299.540 ;
        RECT 37.700 260.155 38.080 260.535 ;
        RECT 37.740 221.150 38.020 260.155 ;
        RECT 37.700 220.770 38.080 221.150 ;
        RECT 37.740 181.765 38.020 220.770 ;
        RECT 37.700 181.385 38.080 181.765 ;
        RECT 37.740 142.380 38.020 181.385 ;
        RECT 37.700 142.000 38.080 142.380 ;
        RECT 37.740 102.995 38.020 142.000 ;
        RECT 37.700 102.615 38.080 102.995 ;
        RECT 37.740 63.610 38.020 102.615 ;
        RECT 37.700 63.230 38.080 63.610 ;
        RECT 37.740 24.225 38.020 63.230 ;
        RECT 37.700 23.845 38.080 24.225 ;
        RECT 37.740 0.000 38.020 23.845 ;
    END
  END BIT_SEL[0]
  PIN BIT_SEL[1]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 37.100 291.355 37.380 315.200 ;
        RECT 37.060 290.975 37.440 291.355 ;
        RECT 37.100 251.970 37.380 290.975 ;
        RECT 37.060 251.590 37.440 251.970 ;
        RECT 37.100 212.585 37.380 251.590 ;
        RECT 37.060 212.205 37.440 212.585 ;
        RECT 37.100 173.200 37.380 212.205 ;
        RECT 37.060 172.820 37.440 173.200 ;
        RECT 37.100 133.815 37.380 172.820 ;
        RECT 37.060 133.435 37.440 133.815 ;
        RECT 37.100 94.430 37.380 133.435 ;
        RECT 37.060 94.050 37.440 94.430 ;
        RECT 37.100 55.045 37.380 94.050 ;
        RECT 37.060 54.665 37.440 55.045 ;
        RECT 37.100 15.660 37.380 54.665 ;
        RECT 37.060 15.280 37.440 15.660 ;
        RECT 37.100 0.000 37.380 15.280 ;
    END
  END BIT_SEL[1]
  PIN BIT_SEL[2]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 36.460 301.760 36.740 315.200 ;
        RECT 36.420 301.380 36.800 301.760 ;
        RECT 36.460 262.375 36.740 301.380 ;
        RECT 36.420 261.995 36.800 262.375 ;
        RECT 36.460 222.990 36.740 261.995 ;
        RECT 36.420 222.610 36.800 222.990 ;
        RECT 36.460 183.605 36.740 222.610 ;
        RECT 36.420 183.225 36.800 183.605 ;
        RECT 36.460 144.220 36.740 183.225 ;
        RECT 36.420 143.840 36.800 144.220 ;
        RECT 36.460 104.835 36.740 143.840 ;
        RECT 36.420 104.455 36.800 104.835 ;
        RECT 36.460 65.450 36.740 104.455 ;
        RECT 36.420 65.070 36.800 65.450 ;
        RECT 36.460 26.065 36.740 65.070 ;
        RECT 36.420 25.685 36.800 26.065 ;
        RECT 36.460 0.000 36.740 25.685 ;
    END
  END BIT_SEL[2]
  PIN BIT_SEL[3]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 35.820 289.515 36.100 315.200 ;
        RECT 35.780 289.135 36.160 289.515 ;
        RECT 35.820 250.130 36.100 289.135 ;
        RECT 35.780 249.750 36.160 250.130 ;
        RECT 35.820 210.745 36.100 249.750 ;
        RECT 35.780 210.365 36.160 210.745 ;
        RECT 35.820 171.360 36.100 210.365 ;
        RECT 35.780 170.980 36.160 171.360 ;
        RECT 35.820 131.975 36.100 170.980 ;
        RECT 35.780 131.595 36.160 131.975 ;
        RECT 35.820 92.590 36.100 131.595 ;
        RECT 35.780 92.210 36.160 92.590 ;
        RECT 35.820 53.205 36.100 92.210 ;
        RECT 35.780 52.825 36.160 53.205 ;
        RECT 35.820 13.820 36.100 52.825 ;
        RECT 35.780 13.440 36.160 13.820 ;
        RECT 35.820 0.000 36.100 13.440 ;
    END
  END BIT_SEL[3]
  PIN BIT_SEL[4]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 35.180 303.600 35.460 315.200 ;
        RECT 35.140 303.220 35.520 303.600 ;
        RECT 35.180 264.215 35.460 303.220 ;
        RECT 35.140 263.835 35.520 264.215 ;
        RECT 35.180 224.830 35.460 263.835 ;
        RECT 35.140 224.450 35.520 224.830 ;
        RECT 35.180 185.445 35.460 224.450 ;
        RECT 35.140 185.065 35.520 185.445 ;
        RECT 35.180 146.060 35.460 185.065 ;
        RECT 35.140 145.680 35.520 146.060 ;
        RECT 35.180 106.675 35.460 145.680 ;
        RECT 35.140 106.295 35.520 106.675 ;
        RECT 35.180 67.290 35.460 106.295 ;
        RECT 35.140 66.910 35.520 67.290 ;
        RECT 35.180 27.905 35.460 66.910 ;
        RECT 35.140 27.525 35.520 27.905 ;
        RECT 35.180 0.000 35.460 27.525 ;
    END
  END BIT_SEL[4]
  PIN BIT_SEL[17]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 69.550 291.355 69.830 315.200 ;
        RECT 69.510 290.975 69.890 291.355 ;
        RECT 69.550 251.970 69.830 290.975 ;
        RECT 69.510 251.590 69.890 251.970 ;
        RECT 69.550 212.585 69.830 251.590 ;
        RECT 69.510 212.205 69.890 212.585 ;
        RECT 69.550 173.200 69.830 212.205 ;
        RECT 69.510 172.820 69.890 173.200 ;
        RECT 69.550 133.815 69.830 172.820 ;
        RECT 69.510 133.435 69.890 133.815 ;
        RECT 69.550 94.430 69.830 133.435 ;
        RECT 69.510 94.050 69.890 94.430 ;
        RECT 69.550 55.045 69.830 94.050 ;
        RECT 69.510 54.665 69.890 55.045 ;
        RECT 69.550 15.660 69.830 54.665 ;
        RECT 69.510 15.280 69.890 15.660 ;
        RECT 69.550 0.000 69.830 15.280 ;
    END
  END BIT_SEL[17]
  PIN BIT_SEL[18]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 68.910 301.760 69.190 315.200 ;
        RECT 68.870 301.380 69.250 301.760 ;
        RECT 68.910 262.375 69.190 301.380 ;
        RECT 68.870 261.995 69.250 262.375 ;
        RECT 68.910 222.990 69.190 261.995 ;
        RECT 68.870 222.610 69.250 222.990 ;
        RECT 68.910 183.605 69.190 222.610 ;
        RECT 68.870 183.225 69.250 183.605 ;
        RECT 68.910 144.220 69.190 183.225 ;
        RECT 68.870 143.840 69.250 144.220 ;
        RECT 68.910 104.835 69.190 143.840 ;
        RECT 68.870 104.455 69.250 104.835 ;
        RECT 68.910 65.450 69.190 104.455 ;
        RECT 68.870 65.070 69.250 65.450 ;
        RECT 68.910 26.065 69.190 65.070 ;
        RECT 68.870 25.685 69.250 26.065 ;
        RECT 68.910 0.000 69.190 25.685 ;
    END
  END BIT_SEL[18]
  PIN BIT_SEL[19]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 68.270 289.515 68.550 315.200 ;
        RECT 68.230 289.135 68.610 289.515 ;
        RECT 68.270 250.130 68.550 289.135 ;
        RECT 68.230 249.750 68.610 250.130 ;
        RECT 68.270 210.745 68.550 249.750 ;
        RECT 68.230 210.365 68.610 210.745 ;
        RECT 68.270 171.360 68.550 210.365 ;
        RECT 68.230 170.980 68.610 171.360 ;
        RECT 68.270 131.975 68.550 170.980 ;
        RECT 68.230 131.595 68.610 131.975 ;
        RECT 68.270 92.590 68.550 131.595 ;
        RECT 68.230 92.210 68.610 92.590 ;
        RECT 68.270 53.205 68.550 92.210 ;
        RECT 68.230 52.825 68.610 53.205 ;
        RECT 68.270 13.820 68.550 52.825 ;
        RECT 68.230 13.440 68.610 13.820 ;
        RECT 68.270 0.000 68.550 13.440 ;
    END
  END BIT_SEL[19]
  PIN BIT_SEL[20]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 67.630 303.600 67.910 315.200 ;
        RECT 67.590 303.220 67.970 303.600 ;
        RECT 67.630 264.215 67.910 303.220 ;
        RECT 67.590 263.835 67.970 264.215 ;
        RECT 67.630 224.830 67.910 263.835 ;
        RECT 67.590 224.450 67.970 224.830 ;
        RECT 67.630 185.445 67.910 224.450 ;
        RECT 67.590 185.065 67.970 185.445 ;
        RECT 67.630 146.060 67.910 185.065 ;
        RECT 67.590 145.680 67.970 146.060 ;
        RECT 67.630 106.675 67.910 145.680 ;
        RECT 67.590 106.295 67.970 106.675 ;
        RECT 67.630 67.290 67.910 106.295 ;
        RECT 67.590 66.910 67.970 67.290 ;
        RECT 67.630 27.905 67.910 66.910 ;
        RECT 67.590 27.525 67.970 27.905 ;
        RECT 67.630 0.000 67.910 27.525 ;
    END
  END BIT_SEL[20]
  PIN BIT_SEL[21]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 66.990 287.670 67.270 315.200 ;
        RECT 66.950 287.290 67.330 287.670 ;
        RECT 66.990 248.285 67.270 287.290 ;
        RECT 66.950 247.905 67.330 248.285 ;
        RECT 66.990 208.900 67.270 247.905 ;
        RECT 66.950 208.520 67.330 208.900 ;
        RECT 66.990 169.515 67.270 208.520 ;
        RECT 66.950 169.135 67.330 169.515 ;
        RECT 66.990 130.130 67.270 169.135 ;
        RECT 66.950 129.750 67.330 130.130 ;
        RECT 66.990 90.745 67.270 129.750 ;
        RECT 66.950 90.365 67.330 90.745 ;
        RECT 66.990 51.360 67.270 90.365 ;
        RECT 66.950 50.980 67.330 51.360 ;
        RECT 66.990 11.975 67.270 50.980 ;
        RECT 66.950 11.595 67.330 11.975 ;
        RECT 66.990 0.000 67.270 11.595 ;
    END
  END BIT_SEL[21]
  PIN BIT_SEL[22]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 66.350 306.245 66.630 315.200 ;
        RECT 66.310 305.865 66.690 306.245 ;
        RECT 66.350 266.860 66.630 305.865 ;
        RECT 66.310 266.480 66.690 266.860 ;
        RECT 66.350 227.475 66.630 266.480 ;
        RECT 66.310 227.095 66.690 227.475 ;
        RECT 66.350 188.090 66.630 227.095 ;
        RECT 66.310 187.710 66.690 188.090 ;
        RECT 66.350 148.705 66.630 187.710 ;
        RECT 66.310 148.325 66.690 148.705 ;
        RECT 66.350 109.320 66.630 148.325 ;
        RECT 66.310 108.940 66.690 109.320 ;
        RECT 66.350 69.935 66.630 108.940 ;
        RECT 66.310 69.555 66.690 69.935 ;
        RECT 66.350 30.550 66.630 69.555 ;
        RECT 66.310 30.170 66.690 30.550 ;
        RECT 66.350 0.000 66.630 30.170 ;
    END
  END BIT_SEL[22]
  PIN BIT_SEL[23]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 65.710 285.030 65.990 315.200 ;
        RECT 65.670 284.650 66.050 285.030 ;
        RECT 65.710 245.645 65.990 284.650 ;
        RECT 65.670 245.265 66.050 245.645 ;
        RECT 65.710 206.260 65.990 245.265 ;
        RECT 65.670 205.880 66.050 206.260 ;
        RECT 65.710 166.875 65.990 205.880 ;
        RECT 65.670 166.495 66.050 166.875 ;
        RECT 65.710 127.490 65.990 166.495 ;
        RECT 65.670 127.110 66.050 127.490 ;
        RECT 65.710 88.105 65.990 127.110 ;
        RECT 65.670 87.725 66.050 88.105 ;
        RECT 65.710 48.720 65.990 87.725 ;
        RECT 65.670 48.340 66.050 48.720 ;
        RECT 65.710 9.335 65.990 48.340 ;
        RECT 65.670 8.955 66.050 9.335 ;
        RECT 65.710 0.000 65.990 8.955 ;
    END
  END BIT_SEL[23]
  PIN BIT_SEL[24]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 65.070 308.085 65.350 315.200 ;
        RECT 65.030 307.705 65.410 308.085 ;
        RECT 65.070 268.700 65.350 307.705 ;
        RECT 65.030 268.320 65.410 268.700 ;
        RECT 65.070 229.315 65.350 268.320 ;
        RECT 65.030 228.935 65.410 229.315 ;
        RECT 65.070 189.930 65.350 228.935 ;
        RECT 65.030 189.550 65.410 189.930 ;
        RECT 65.070 150.545 65.350 189.550 ;
        RECT 65.030 150.165 65.410 150.545 ;
        RECT 65.070 111.160 65.350 150.165 ;
        RECT 65.030 110.780 65.410 111.160 ;
        RECT 65.070 71.775 65.350 110.780 ;
        RECT 65.030 71.395 65.410 71.775 ;
        RECT 65.070 32.390 65.350 71.395 ;
        RECT 65.030 32.010 65.410 32.390 ;
        RECT 65.070 0.000 65.350 32.010 ;
    END
  END BIT_SEL[24]
  PIN BIT_SEL[25]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 64.430 283.190 64.710 315.200 ;
        RECT 64.390 282.810 64.770 283.190 ;
        RECT 64.430 243.805 64.710 282.810 ;
        RECT 64.390 243.425 64.770 243.805 ;
        RECT 64.430 204.420 64.710 243.425 ;
        RECT 64.390 204.040 64.770 204.420 ;
        RECT 64.430 165.035 64.710 204.040 ;
        RECT 64.390 164.655 64.770 165.035 ;
        RECT 64.430 125.650 64.710 164.655 ;
        RECT 64.390 125.270 64.770 125.650 ;
        RECT 64.430 86.265 64.710 125.270 ;
        RECT 64.390 85.885 64.770 86.265 ;
        RECT 64.430 46.880 64.710 85.885 ;
        RECT 64.390 46.500 64.770 46.880 ;
        RECT 64.430 7.495 64.710 46.500 ;
        RECT 64.390 7.115 64.770 7.495 ;
        RECT 64.430 0.000 64.710 7.115 ;
    END
  END BIT_SEL[25]
  PIN BIT_SEL[26]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 63.790 309.925 64.070 315.200 ;
        RECT 63.750 309.545 64.130 309.925 ;
        RECT 63.790 270.540 64.070 309.545 ;
        RECT 63.750 270.160 64.130 270.540 ;
        RECT 63.790 231.155 64.070 270.160 ;
        RECT 63.750 230.775 64.130 231.155 ;
        RECT 63.790 191.770 64.070 230.775 ;
        RECT 63.750 191.390 64.130 191.770 ;
        RECT 63.790 152.385 64.070 191.390 ;
        RECT 63.750 152.005 64.130 152.385 ;
        RECT 63.790 113.000 64.070 152.005 ;
        RECT 63.750 112.620 64.130 113.000 ;
        RECT 63.790 73.615 64.070 112.620 ;
        RECT 63.750 73.235 64.130 73.615 ;
        RECT 63.790 34.230 64.070 73.235 ;
        RECT 63.750 33.850 64.130 34.230 ;
        RECT 63.790 0.000 64.070 33.850 ;
    END
  END BIT_SEL[26]
  PIN BIT_SEL[27]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 63.150 281.345 63.430 315.200 ;
        RECT 63.110 280.965 63.490 281.345 ;
        RECT 63.150 241.960 63.430 280.965 ;
        RECT 63.110 241.580 63.490 241.960 ;
        RECT 63.150 202.575 63.430 241.580 ;
        RECT 63.110 202.195 63.490 202.575 ;
        RECT 63.150 163.190 63.430 202.195 ;
        RECT 63.110 162.810 63.490 163.190 ;
        RECT 63.150 123.805 63.430 162.810 ;
        RECT 63.110 123.425 63.490 123.805 ;
        RECT 63.150 84.420 63.430 123.425 ;
        RECT 63.110 84.040 63.490 84.420 ;
        RECT 63.150 45.035 63.430 84.040 ;
        RECT 63.110 44.655 63.490 45.035 ;
        RECT 63.150 5.650 63.430 44.655 ;
        RECT 63.110 5.270 63.490 5.650 ;
        RECT 63.150 0.000 63.430 5.270 ;
    END
  END BIT_SEL[27]
  PIN BIT_SEL[28]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 62.510 312.570 62.790 315.200 ;
        RECT 62.470 312.190 62.850 312.570 ;
        RECT 62.510 273.185 62.790 312.190 ;
        RECT 62.470 272.805 62.850 273.185 ;
        RECT 62.510 233.800 62.790 272.805 ;
        RECT 62.470 233.420 62.850 233.800 ;
        RECT 62.510 194.415 62.790 233.420 ;
        RECT 62.470 194.035 62.850 194.415 ;
        RECT 62.510 155.030 62.790 194.035 ;
        RECT 62.470 154.650 62.850 155.030 ;
        RECT 62.510 115.645 62.790 154.650 ;
        RECT 62.470 115.265 62.850 115.645 ;
        RECT 62.510 76.260 62.790 115.265 ;
        RECT 62.470 75.880 62.850 76.260 ;
        RECT 62.510 36.875 62.790 75.880 ;
        RECT 62.470 36.495 62.850 36.875 ;
        RECT 62.510 0.000 62.790 36.495 ;
    END
  END BIT_SEL[28]
  PIN BIT_SEL[29]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 61.870 278.705 62.150 315.200 ;
        RECT 61.830 278.325 62.210 278.705 ;
        RECT 61.870 239.320 62.150 278.325 ;
        RECT 61.830 238.940 62.210 239.320 ;
        RECT 61.870 199.935 62.150 238.940 ;
        RECT 61.830 199.555 62.210 199.935 ;
        RECT 61.870 160.550 62.150 199.555 ;
        RECT 61.830 160.170 62.210 160.550 ;
        RECT 61.870 121.165 62.150 160.170 ;
        RECT 61.830 120.785 62.210 121.165 ;
        RECT 61.870 81.780 62.150 120.785 ;
        RECT 61.830 81.400 62.210 81.780 ;
        RECT 61.870 42.395 62.150 81.400 ;
        RECT 61.830 42.015 62.210 42.395 ;
        RECT 61.870 3.010 62.150 42.015 ;
        RECT 61.830 2.630 62.210 3.010 ;
        RECT 61.870 0.000 62.150 2.630 ;
    END
  END BIT_SEL[29]
  PIN BIT_SEL[30]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 61.230 314.410 61.510 315.200 ;
        RECT 61.190 314.030 61.570 314.410 ;
        RECT 61.230 275.025 61.510 314.030 ;
        RECT 61.190 274.645 61.570 275.025 ;
        RECT 61.230 235.640 61.510 274.645 ;
        RECT 61.190 235.260 61.570 235.640 ;
        RECT 61.230 196.255 61.510 235.260 ;
        RECT 61.190 195.875 61.570 196.255 ;
        RECT 61.230 156.870 61.510 195.875 ;
        RECT 61.190 156.490 61.570 156.870 ;
        RECT 61.230 117.485 61.510 156.490 ;
        RECT 61.190 117.105 61.570 117.485 ;
        RECT 61.230 78.100 61.510 117.105 ;
        RECT 61.190 77.720 61.570 78.100 ;
        RECT 61.230 38.715 61.510 77.720 ;
        RECT 61.190 38.335 61.570 38.715 ;
        RECT 61.230 0.000 61.510 38.335 ;
    END
  END BIT_SEL[30]
  PIN BIT_SEL[31]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 60.590 276.865 60.870 315.200 ;
        RECT 60.550 276.485 60.930 276.865 ;
        RECT 60.590 237.480 60.870 276.485 ;
        RECT 60.550 237.100 60.930 237.480 ;
        RECT 60.590 198.095 60.870 237.100 ;
        RECT 60.550 197.715 60.930 198.095 ;
        RECT 60.590 158.710 60.870 197.715 ;
        RECT 60.550 158.330 60.930 158.710 ;
        RECT 60.590 119.325 60.870 158.330 ;
        RECT 60.550 118.945 60.930 119.325 ;
        RECT 60.590 79.940 60.870 118.945 ;
        RECT 60.550 79.560 60.930 79.940 ;
        RECT 60.590 40.555 60.870 79.560 ;
        RECT 60.550 40.175 60.930 40.555 ;
        RECT 60.590 1.170 60.870 40.175 ;
        RECT 60.550 0.790 60.930 1.170 ;
        RECT 60.590 0.000 60.870 0.790 ;
    END
  END BIT_SEL[31]
  PIN BIT_SEL[5]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 34.540 287.670 34.820 315.200 ;
        RECT 34.500 287.290 34.880 287.670 ;
        RECT 34.540 248.285 34.820 287.290 ;
        RECT 34.500 247.905 34.880 248.285 ;
        RECT 34.540 208.900 34.820 247.905 ;
        RECT 34.500 208.520 34.880 208.900 ;
        RECT 34.540 169.515 34.820 208.520 ;
        RECT 34.500 169.135 34.880 169.515 ;
        RECT 34.540 130.130 34.820 169.135 ;
        RECT 34.500 129.750 34.880 130.130 ;
        RECT 34.540 90.745 34.820 129.750 ;
        RECT 34.500 90.365 34.880 90.745 ;
        RECT 34.540 51.360 34.820 90.365 ;
        RECT 34.500 50.980 34.880 51.360 ;
        RECT 34.540 11.975 34.820 50.980 ;
        RECT 34.500 11.595 34.880 11.975 ;
        RECT 34.540 0.000 34.820 11.595 ;
    END
  END BIT_SEL[5]
  PIN BIT_SEL[6]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 33.900 306.245 34.180 315.200 ;
        RECT 33.860 305.865 34.240 306.245 ;
        RECT 33.900 266.860 34.180 305.865 ;
        RECT 33.860 266.480 34.240 266.860 ;
        RECT 33.900 227.475 34.180 266.480 ;
        RECT 33.860 227.095 34.240 227.475 ;
        RECT 33.900 188.090 34.180 227.095 ;
        RECT 33.860 187.710 34.240 188.090 ;
        RECT 33.900 148.705 34.180 187.710 ;
        RECT 33.860 148.325 34.240 148.705 ;
        RECT 33.900 109.320 34.180 148.325 ;
        RECT 33.860 108.940 34.240 109.320 ;
        RECT 33.900 69.935 34.180 108.940 ;
        RECT 33.860 69.555 34.240 69.935 ;
        RECT 33.900 30.550 34.180 69.555 ;
        RECT 33.860 30.170 34.240 30.550 ;
        RECT 33.900 0.000 34.180 30.170 ;
    END
  END BIT_SEL[6]
  PIN BIT_SEL[7]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 33.260 285.030 33.540 315.200 ;
        RECT 33.220 284.650 33.600 285.030 ;
        RECT 33.260 245.645 33.540 284.650 ;
        RECT 33.220 245.265 33.600 245.645 ;
        RECT 33.260 206.260 33.540 245.265 ;
        RECT 33.220 205.880 33.600 206.260 ;
        RECT 33.260 166.875 33.540 205.880 ;
        RECT 33.220 166.495 33.600 166.875 ;
        RECT 33.260 127.490 33.540 166.495 ;
        RECT 33.220 127.110 33.600 127.490 ;
        RECT 33.260 88.105 33.540 127.110 ;
        RECT 33.220 87.725 33.600 88.105 ;
        RECT 33.260 48.720 33.540 87.725 ;
        RECT 33.220 48.340 33.600 48.720 ;
        RECT 33.260 9.335 33.540 48.340 ;
        RECT 33.220 8.955 33.600 9.335 ;
        RECT 33.260 0.000 33.540 8.955 ;
    END
  END BIT_SEL[7]
  PIN BIT_SEL[8]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 32.620 308.085 32.900 315.200 ;
        RECT 32.580 307.705 32.960 308.085 ;
        RECT 32.620 268.700 32.900 307.705 ;
        RECT 32.580 268.320 32.960 268.700 ;
        RECT 32.620 229.315 32.900 268.320 ;
        RECT 32.580 228.935 32.960 229.315 ;
        RECT 32.620 189.930 32.900 228.935 ;
        RECT 32.580 189.550 32.960 189.930 ;
        RECT 32.620 150.545 32.900 189.550 ;
        RECT 32.580 150.165 32.960 150.545 ;
        RECT 32.620 111.160 32.900 150.165 ;
        RECT 32.580 110.780 32.960 111.160 ;
        RECT 32.620 71.775 32.900 110.780 ;
        RECT 32.580 71.395 32.960 71.775 ;
        RECT 32.620 32.390 32.900 71.395 ;
        RECT 32.580 32.010 32.960 32.390 ;
        RECT 32.620 0.000 32.900 32.010 ;
    END
  END BIT_SEL[8]
  PIN BIT_SEL[9]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 31.980 283.190 32.260 315.200 ;
        RECT 31.940 282.810 32.320 283.190 ;
        RECT 31.980 243.805 32.260 282.810 ;
        RECT 31.940 243.425 32.320 243.805 ;
        RECT 31.980 204.420 32.260 243.425 ;
        RECT 31.940 204.040 32.320 204.420 ;
        RECT 31.980 165.035 32.260 204.040 ;
        RECT 31.940 164.655 32.320 165.035 ;
        RECT 31.980 125.650 32.260 164.655 ;
        RECT 31.940 125.270 32.320 125.650 ;
        RECT 31.980 86.265 32.260 125.270 ;
        RECT 31.940 85.885 32.320 86.265 ;
        RECT 31.980 46.880 32.260 85.885 ;
        RECT 31.940 46.500 32.320 46.880 ;
        RECT 31.980 7.495 32.260 46.500 ;
        RECT 31.940 7.115 32.320 7.495 ;
        RECT 31.980 0.000 32.260 7.115 ;
    END
  END BIT_SEL[9]
  PIN BIT_SEL[10]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 31.340 309.925 31.620 315.200 ;
        RECT 31.300 309.545 31.680 309.925 ;
        RECT 31.340 270.540 31.620 309.545 ;
        RECT 31.300 270.160 31.680 270.540 ;
        RECT 31.340 231.155 31.620 270.160 ;
        RECT 31.300 230.775 31.680 231.155 ;
        RECT 31.340 191.770 31.620 230.775 ;
        RECT 31.300 191.390 31.680 191.770 ;
        RECT 31.340 152.385 31.620 191.390 ;
        RECT 31.300 152.005 31.680 152.385 ;
        RECT 31.340 113.000 31.620 152.005 ;
        RECT 31.300 112.620 31.680 113.000 ;
        RECT 31.340 73.615 31.620 112.620 ;
        RECT 31.300 73.235 31.680 73.615 ;
        RECT 31.340 34.230 31.620 73.235 ;
        RECT 31.300 33.850 31.680 34.230 ;
        RECT 31.340 0.000 31.620 33.850 ;
    END
  END BIT_SEL[10]
  PIN BIT_SEL[11]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 30.700 281.345 30.980 315.200 ;
        RECT 30.660 280.965 31.040 281.345 ;
        RECT 30.700 241.960 30.980 280.965 ;
        RECT 30.660 241.580 31.040 241.960 ;
        RECT 30.700 202.575 30.980 241.580 ;
        RECT 30.660 202.195 31.040 202.575 ;
        RECT 30.700 163.190 30.980 202.195 ;
        RECT 30.660 162.810 31.040 163.190 ;
        RECT 30.700 123.805 30.980 162.810 ;
        RECT 30.660 123.425 31.040 123.805 ;
        RECT 30.700 84.420 30.980 123.425 ;
        RECT 30.660 84.040 31.040 84.420 ;
        RECT 30.700 45.035 30.980 84.040 ;
        RECT 30.660 44.655 31.040 45.035 ;
        RECT 30.700 5.650 30.980 44.655 ;
        RECT 30.660 5.270 31.040 5.650 ;
        RECT 30.700 0.000 30.980 5.270 ;
    END
  END BIT_SEL[11]
  PIN BIT_SEL[12]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 30.060 312.570 30.340 315.200 ;
        RECT 30.020 312.190 30.400 312.570 ;
        RECT 30.060 273.185 30.340 312.190 ;
        RECT 30.020 272.805 30.400 273.185 ;
        RECT 30.060 233.800 30.340 272.805 ;
        RECT 30.020 233.420 30.400 233.800 ;
        RECT 30.060 194.415 30.340 233.420 ;
        RECT 30.020 194.035 30.400 194.415 ;
        RECT 30.060 155.030 30.340 194.035 ;
        RECT 30.020 154.650 30.400 155.030 ;
        RECT 30.060 115.645 30.340 154.650 ;
        RECT 30.020 115.265 30.400 115.645 ;
        RECT 30.060 76.260 30.340 115.265 ;
        RECT 30.020 75.880 30.400 76.260 ;
        RECT 30.060 36.875 30.340 75.880 ;
        RECT 30.020 36.495 30.400 36.875 ;
        RECT 30.060 0.000 30.340 36.495 ;
    END
  END BIT_SEL[12]
  PIN BIT_SEL[13]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 29.420 278.705 29.700 315.200 ;
        RECT 29.380 278.325 29.760 278.705 ;
        RECT 29.420 239.320 29.700 278.325 ;
        RECT 29.380 238.940 29.760 239.320 ;
        RECT 29.420 199.935 29.700 238.940 ;
        RECT 29.380 199.555 29.760 199.935 ;
        RECT 29.420 160.550 29.700 199.555 ;
        RECT 29.380 160.170 29.760 160.550 ;
        RECT 29.420 121.165 29.700 160.170 ;
        RECT 29.380 120.785 29.760 121.165 ;
        RECT 29.420 81.780 29.700 120.785 ;
        RECT 29.380 81.400 29.760 81.780 ;
        RECT 29.420 42.395 29.700 81.400 ;
        RECT 29.380 42.015 29.760 42.395 ;
        RECT 29.420 3.010 29.700 42.015 ;
        RECT 29.380 2.630 29.760 3.010 ;
        RECT 29.420 0.000 29.700 2.630 ;
    END
  END BIT_SEL[13]
  PIN BIT_SEL[14]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 28.780 314.410 29.060 315.200 ;
        RECT 28.740 314.030 29.120 314.410 ;
        RECT 28.780 275.025 29.060 314.030 ;
        RECT 28.740 274.645 29.120 275.025 ;
        RECT 28.780 235.640 29.060 274.645 ;
        RECT 28.740 235.260 29.120 235.640 ;
        RECT 28.780 196.255 29.060 235.260 ;
        RECT 28.740 195.875 29.120 196.255 ;
        RECT 28.780 156.870 29.060 195.875 ;
        RECT 28.740 156.490 29.120 156.870 ;
        RECT 28.780 117.485 29.060 156.490 ;
        RECT 28.740 117.105 29.120 117.485 ;
        RECT 28.780 78.100 29.060 117.105 ;
        RECT 28.740 77.720 29.120 78.100 ;
        RECT 28.780 38.715 29.060 77.720 ;
        RECT 28.740 38.335 29.120 38.715 ;
        RECT 28.780 0.000 29.060 38.335 ;
    END
  END BIT_SEL[14]
  PIN BIT_SEL[15]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 28.140 276.865 28.420 315.200 ;
        RECT 28.100 276.485 28.480 276.865 ;
        RECT 28.140 237.480 28.420 276.485 ;
        RECT 28.100 237.100 28.480 237.480 ;
        RECT 28.140 198.095 28.420 237.100 ;
        RECT 28.100 197.715 28.480 198.095 ;
        RECT 28.140 158.710 28.420 197.715 ;
        RECT 28.100 158.330 28.480 158.710 ;
        RECT 28.140 119.325 28.420 158.330 ;
        RECT 28.100 118.945 28.480 119.325 ;
        RECT 28.140 79.940 28.420 118.945 ;
        RECT 28.100 79.560 28.480 79.940 ;
        RECT 28.140 40.555 28.420 79.560 ;
        RECT 28.100 40.175 28.480 40.555 ;
        RECT 28.140 1.170 28.420 40.175 ;
        RECT 28.100 0.790 28.480 1.170 ;
        RECT 28.140 0.000 28.420 0.790 ;
    END
  END BIT_SEL[15]
  OBS
      LAYER Metal1 ;
        RECT 0.130 314.915 0.730 315.825 ;
        RECT 4.050 314.915 4.650 315.825 ;
        RECT 0.130 314.575 2.430 314.915 ;
        RECT 3.160 314.575 4.650 314.915 ;
        RECT 6.690 314.590 37.210 314.970 ;
        RECT 39.140 314.590 69.660 314.970 ;
        RECT 71.590 314.590 102.110 314.970 ;
        RECT 104.040 314.590 134.560 314.970 ;
        RECT 0.130 313.960 0.730 314.575 ;
        RECT 0.130 313.730 1.860 313.960 ;
        RECT 2.160 313.730 3.820 313.960 ;
        RECT 0.130 311.720 0.730 313.730 ;
        RECT 2.160 312.695 2.390 313.730 ;
        RECT 2.795 312.440 3.025 313.485 ;
        RECT 4.050 312.440 4.650 314.575 ;
        RECT 5.840 314.335 6.460 314.520 ;
        RECT 37.440 314.335 38.060 314.520 ;
        RECT 5.840 314.105 38.060 314.335 ;
        RECT 5.840 313.920 6.460 314.105 ;
        RECT 37.440 313.920 38.060 314.105 ;
        RECT 38.290 314.335 38.910 314.520 ;
        RECT 69.890 314.335 70.510 314.520 ;
        RECT 38.290 314.105 70.510 314.335 ;
        RECT 38.290 313.920 38.910 314.105 ;
        RECT 69.890 313.920 70.510 314.105 ;
        RECT 70.740 314.335 71.360 314.520 ;
        RECT 102.340 314.335 102.960 314.520 ;
        RECT 70.740 314.105 102.960 314.335 ;
        RECT 70.740 313.920 71.360 314.105 ;
        RECT 102.340 313.920 102.960 314.105 ;
        RECT 103.190 314.335 103.810 314.520 ;
        RECT 134.790 314.335 135.410 314.520 ;
        RECT 103.190 314.105 135.410 314.335 ;
        RECT 103.190 313.920 103.810 314.105 ;
        RECT 134.790 313.920 135.410 314.105 ;
        RECT 33.440 313.840 35.060 313.850 ;
        RECT 65.890 313.840 67.510 313.850 ;
        RECT 98.340 313.840 99.960 313.850 ;
        RECT 130.790 313.840 132.410 313.850 ;
        RECT 6.690 313.470 37.210 313.840 ;
        RECT 39.140 313.470 69.660 313.840 ;
        RECT 71.590 313.470 102.110 313.840 ;
        RECT 104.040 313.470 134.560 313.840 ;
        RECT 6.690 312.750 37.210 313.130 ;
        RECT 39.140 312.750 69.660 313.130 ;
        RECT 71.590 312.750 102.110 313.130 ;
        RECT 104.040 312.750 134.560 313.130 ;
        RECT 0.960 312.210 3.025 312.440 ;
        RECT 3.255 312.210 4.650 312.440 ;
        RECT 0.130 311.490 1.860 311.720 ;
        RECT 2.160 311.490 3.820 311.720 ;
        RECT 0.130 309.480 0.730 311.490 ;
        RECT 2.160 310.455 2.390 311.490 ;
        RECT 2.795 310.200 3.025 311.245 ;
        RECT 4.050 310.200 4.650 312.210 ;
        RECT 5.840 312.495 6.460 312.680 ;
        RECT 37.440 312.495 38.060 312.680 ;
        RECT 5.840 312.265 38.060 312.495 ;
        RECT 5.840 312.080 6.460 312.265 ;
        RECT 37.440 312.080 38.060 312.265 ;
        RECT 38.290 312.495 38.910 312.680 ;
        RECT 69.890 312.495 70.510 312.680 ;
        RECT 38.290 312.265 70.510 312.495 ;
        RECT 38.290 312.080 38.910 312.265 ;
        RECT 69.890 312.080 70.510 312.265 ;
        RECT 70.740 312.495 71.360 312.680 ;
        RECT 102.340 312.495 102.960 312.680 ;
        RECT 70.740 312.265 102.960 312.495 ;
        RECT 70.740 312.080 71.360 312.265 ;
        RECT 102.340 312.080 102.960 312.265 ;
        RECT 103.190 312.495 103.810 312.680 ;
        RECT 134.790 312.495 135.410 312.680 ;
        RECT 103.190 312.265 135.410 312.495 ;
        RECT 103.190 312.080 103.810 312.265 ;
        RECT 134.790 312.080 135.410 312.265 ;
        RECT 29.600 312.000 31.220 312.010 ;
        RECT 62.050 312.000 63.670 312.010 ;
        RECT 94.500 312.000 96.120 312.010 ;
        RECT 126.950 312.000 128.570 312.010 ;
        RECT 6.690 311.630 37.210 312.000 ;
        RECT 39.140 311.630 69.660 312.000 ;
        RECT 71.590 311.630 102.110 312.000 ;
        RECT 104.040 311.630 134.560 312.000 ;
        RECT 6.700 310.835 37.200 311.275 ;
        RECT 39.150 310.835 69.650 311.275 ;
        RECT 71.600 310.835 102.100 311.275 ;
        RECT 104.050 310.835 134.550 311.275 ;
        RECT 0.960 309.970 3.025 310.200 ;
        RECT 3.255 309.970 4.650 310.200 ;
        RECT 6.690 310.105 37.210 310.485 ;
        RECT 39.140 310.105 69.660 310.485 ;
        RECT 71.590 310.105 102.110 310.485 ;
        RECT 104.040 310.105 134.560 310.485 ;
        RECT 0.130 309.250 1.860 309.480 ;
        RECT 2.160 309.250 3.820 309.480 ;
        RECT 0.130 307.240 0.730 309.250 ;
        RECT 2.160 308.215 2.390 309.250 ;
        RECT 2.795 307.960 3.025 309.005 ;
        RECT 4.050 307.960 4.650 309.970 ;
        RECT 5.840 309.850 6.460 310.035 ;
        RECT 37.440 309.850 38.060 310.035 ;
        RECT 5.840 309.620 38.060 309.850 ;
        RECT 5.840 309.435 6.460 309.620 ;
        RECT 37.440 309.435 38.060 309.620 ;
        RECT 38.290 309.850 38.910 310.035 ;
        RECT 69.890 309.850 70.510 310.035 ;
        RECT 38.290 309.620 70.510 309.850 ;
        RECT 38.290 309.435 38.910 309.620 ;
        RECT 69.890 309.435 70.510 309.620 ;
        RECT 70.740 309.850 71.360 310.035 ;
        RECT 102.340 309.850 102.960 310.035 ;
        RECT 70.740 309.620 102.960 309.850 ;
        RECT 70.740 309.435 71.360 309.620 ;
        RECT 102.340 309.435 102.960 309.620 ;
        RECT 103.190 309.850 103.810 310.035 ;
        RECT 134.790 309.850 135.410 310.035 ;
        RECT 103.190 309.620 135.410 309.850 ;
        RECT 103.190 309.435 103.810 309.620 ;
        RECT 134.790 309.435 135.410 309.620 ;
        RECT 25.760 309.355 27.380 309.365 ;
        RECT 58.210 309.355 59.830 309.365 ;
        RECT 90.660 309.355 92.280 309.365 ;
        RECT 123.110 309.355 124.730 309.365 ;
        RECT 6.690 308.985 37.210 309.355 ;
        RECT 39.140 308.985 69.660 309.355 ;
        RECT 71.590 308.985 102.110 309.355 ;
        RECT 104.040 308.985 134.560 309.355 ;
        RECT 6.690 308.265 37.210 308.645 ;
        RECT 39.140 308.265 69.660 308.645 ;
        RECT 71.590 308.265 102.110 308.645 ;
        RECT 104.040 308.265 134.560 308.645 ;
        RECT 0.960 307.730 3.025 307.960 ;
        RECT 3.255 307.730 4.650 307.960 ;
        RECT 0.130 307.010 1.860 307.240 ;
        RECT 2.160 307.010 3.820 307.240 ;
        RECT 0.130 305.000 0.730 307.010 ;
        RECT 2.160 305.975 2.390 307.010 ;
        RECT 2.795 305.720 3.025 306.765 ;
        RECT 4.050 305.720 4.650 307.730 ;
        RECT 5.840 308.010 6.460 308.195 ;
        RECT 37.440 308.010 38.060 308.195 ;
        RECT 5.840 307.780 38.060 308.010 ;
        RECT 5.840 307.595 6.460 307.780 ;
        RECT 37.440 307.595 38.060 307.780 ;
        RECT 38.290 308.010 38.910 308.195 ;
        RECT 69.890 308.010 70.510 308.195 ;
        RECT 38.290 307.780 70.510 308.010 ;
        RECT 38.290 307.595 38.910 307.780 ;
        RECT 69.890 307.595 70.510 307.780 ;
        RECT 70.740 308.010 71.360 308.195 ;
        RECT 102.340 308.010 102.960 308.195 ;
        RECT 70.740 307.780 102.960 308.010 ;
        RECT 70.740 307.595 71.360 307.780 ;
        RECT 102.340 307.595 102.960 307.780 ;
        RECT 103.190 308.010 103.810 308.195 ;
        RECT 134.790 308.010 135.410 308.195 ;
        RECT 103.190 307.780 135.410 308.010 ;
        RECT 103.190 307.595 103.810 307.780 ;
        RECT 134.790 307.595 135.410 307.780 ;
        RECT 21.920 307.515 23.540 307.525 ;
        RECT 54.370 307.515 55.990 307.525 ;
        RECT 86.820 307.515 88.440 307.525 ;
        RECT 119.270 307.515 120.890 307.525 ;
        RECT 6.690 307.145 37.210 307.515 ;
        RECT 39.140 307.145 69.660 307.515 ;
        RECT 71.590 307.145 102.110 307.515 ;
        RECT 104.040 307.145 134.560 307.515 ;
        RECT 6.690 306.425 37.210 306.805 ;
        RECT 39.140 306.425 69.660 306.805 ;
        RECT 71.590 306.425 102.110 306.805 ;
        RECT 104.040 306.425 134.560 306.805 ;
        RECT 5.840 306.170 6.460 306.355 ;
        RECT 37.440 306.170 38.060 306.355 ;
        RECT 5.840 305.940 38.060 306.170 ;
        RECT 5.840 305.755 6.460 305.940 ;
        RECT 37.440 305.755 38.060 305.940 ;
        RECT 38.290 306.170 38.910 306.355 ;
        RECT 69.890 306.170 70.510 306.355 ;
        RECT 38.290 305.940 70.510 306.170 ;
        RECT 38.290 305.755 38.910 305.940 ;
        RECT 69.890 305.755 70.510 305.940 ;
        RECT 70.740 306.170 71.360 306.355 ;
        RECT 102.340 306.170 102.960 306.355 ;
        RECT 70.740 305.940 102.960 306.170 ;
        RECT 70.740 305.755 71.360 305.940 ;
        RECT 102.340 305.755 102.960 305.940 ;
        RECT 103.190 306.170 103.810 306.355 ;
        RECT 134.790 306.170 135.410 306.355 ;
        RECT 103.190 305.940 135.410 306.170 ;
        RECT 103.190 305.755 103.810 305.940 ;
        RECT 134.790 305.755 135.410 305.940 ;
        RECT 0.960 305.490 3.025 305.720 ;
        RECT 3.255 305.490 4.650 305.720 ;
        RECT 18.080 305.675 19.700 305.685 ;
        RECT 50.530 305.675 52.150 305.685 ;
        RECT 82.980 305.675 84.600 305.685 ;
        RECT 115.430 305.675 117.050 305.685 ;
        RECT 0.130 304.770 1.860 305.000 ;
        RECT 2.160 304.770 3.820 305.000 ;
        RECT 0.130 302.615 0.730 304.770 ;
        RECT 2.160 303.735 2.390 304.770 ;
        RECT 2.795 303.480 3.025 304.525 ;
        RECT 4.050 303.480 4.650 305.490 ;
        RECT 6.690 305.305 37.210 305.675 ;
        RECT 39.140 305.305 69.660 305.675 ;
        RECT 71.590 305.305 102.110 305.675 ;
        RECT 104.040 305.305 134.560 305.675 ;
        RECT 6.700 304.510 37.200 304.950 ;
        RECT 39.150 304.510 69.650 304.950 ;
        RECT 71.600 304.510 102.100 304.950 ;
        RECT 104.050 304.510 134.550 304.950 ;
        RECT 6.690 303.780 37.210 304.160 ;
        RECT 39.140 303.780 69.660 304.160 ;
        RECT 71.590 303.780 102.110 304.160 ;
        RECT 104.040 303.780 134.560 304.160 ;
        RECT 0.960 303.250 3.025 303.480 ;
        RECT 3.255 303.250 4.650 303.480 ;
        RECT 4.050 302.615 4.650 303.250 ;
        RECT 5.840 303.525 6.460 303.710 ;
        RECT 37.440 303.525 38.060 303.710 ;
        RECT 5.840 303.295 38.060 303.525 ;
        RECT 5.840 303.110 6.460 303.295 ;
        RECT 37.440 303.110 38.060 303.295 ;
        RECT 38.290 303.525 38.910 303.710 ;
        RECT 69.890 303.525 70.510 303.710 ;
        RECT 38.290 303.295 70.510 303.525 ;
        RECT 38.290 303.110 38.910 303.295 ;
        RECT 69.890 303.110 70.510 303.295 ;
        RECT 70.740 303.525 71.360 303.710 ;
        RECT 102.340 303.525 102.960 303.710 ;
        RECT 70.740 303.295 102.960 303.525 ;
        RECT 70.740 303.110 71.360 303.295 ;
        RECT 102.340 303.110 102.960 303.295 ;
        RECT 103.190 303.525 103.810 303.710 ;
        RECT 134.790 303.525 135.410 303.710 ;
        RECT 103.190 303.295 135.410 303.525 ;
        RECT 103.190 303.110 103.810 303.295 ;
        RECT 134.790 303.110 135.410 303.295 ;
        RECT 14.240 303.030 15.860 303.040 ;
        RECT 46.690 303.030 48.310 303.040 ;
        RECT 79.140 303.030 80.760 303.040 ;
        RECT 111.590 303.030 113.210 303.040 ;
        RECT 6.690 302.660 37.210 303.030 ;
        RECT 39.140 302.660 69.660 303.030 ;
        RECT 71.590 302.660 102.110 303.030 ;
        RECT 104.040 302.660 134.560 303.030 ;
        RECT 0.130 302.275 2.420 302.615 ;
        RECT 3.165 302.275 4.650 302.615 ;
        RECT 0.130 301.640 0.730 302.275 ;
        RECT 0.130 301.410 1.860 301.640 ;
        RECT 2.160 301.410 3.820 301.640 ;
        RECT 0.130 299.400 0.730 301.410 ;
        RECT 2.160 300.375 2.390 301.410 ;
        RECT 2.795 300.120 3.025 301.165 ;
        RECT 4.050 300.120 4.650 302.275 ;
        RECT 6.690 301.940 37.210 302.320 ;
        RECT 39.140 301.940 69.660 302.320 ;
        RECT 71.590 301.940 102.110 302.320 ;
        RECT 104.040 301.940 134.560 302.320 ;
        RECT 5.840 301.685 6.460 301.870 ;
        RECT 37.440 301.685 38.060 301.870 ;
        RECT 5.840 301.455 38.060 301.685 ;
        RECT 5.840 301.270 6.460 301.455 ;
        RECT 37.440 301.270 38.060 301.455 ;
        RECT 38.290 301.685 38.910 301.870 ;
        RECT 69.890 301.685 70.510 301.870 ;
        RECT 38.290 301.455 70.510 301.685 ;
        RECT 38.290 301.270 38.910 301.455 ;
        RECT 69.890 301.270 70.510 301.455 ;
        RECT 70.740 301.685 71.360 301.870 ;
        RECT 102.340 301.685 102.960 301.870 ;
        RECT 70.740 301.455 102.960 301.685 ;
        RECT 70.740 301.270 71.360 301.455 ;
        RECT 102.340 301.270 102.960 301.455 ;
        RECT 103.190 301.685 103.810 301.870 ;
        RECT 134.790 301.685 135.410 301.870 ;
        RECT 103.190 301.455 135.410 301.685 ;
        RECT 103.190 301.270 103.810 301.455 ;
        RECT 134.790 301.270 135.410 301.455 ;
        RECT 10.400 301.190 12.020 301.200 ;
        RECT 42.850 301.190 44.470 301.200 ;
        RECT 75.300 301.190 76.920 301.200 ;
        RECT 107.750 301.190 109.370 301.200 ;
        RECT 6.690 300.820 37.210 301.190 ;
        RECT 39.140 300.820 69.660 301.190 ;
        RECT 71.590 300.820 102.110 301.190 ;
        RECT 104.040 300.820 134.560 301.190 ;
        RECT 0.960 299.890 3.025 300.120 ;
        RECT 3.255 299.890 4.650 300.120 ;
        RECT 6.690 300.100 37.210 300.480 ;
        RECT 39.140 300.100 69.660 300.480 ;
        RECT 71.590 300.100 102.110 300.480 ;
        RECT 104.040 300.100 134.560 300.480 ;
        RECT 0.130 299.170 1.860 299.400 ;
        RECT 2.160 299.170 3.820 299.400 ;
        RECT 0.130 297.015 0.730 299.170 ;
        RECT 2.160 298.135 2.390 299.170 ;
        RECT 2.795 297.880 3.025 298.925 ;
        RECT 4.050 297.880 4.650 299.890 ;
        RECT 5.840 299.845 6.460 300.030 ;
        RECT 37.440 299.845 38.060 300.030 ;
        RECT 5.840 299.615 38.060 299.845 ;
        RECT 5.840 299.430 6.460 299.615 ;
        RECT 37.440 299.430 38.060 299.615 ;
        RECT 38.290 299.845 38.910 300.030 ;
        RECT 69.890 299.845 70.510 300.030 ;
        RECT 38.290 299.615 70.510 299.845 ;
        RECT 38.290 299.430 38.910 299.615 ;
        RECT 69.890 299.430 70.510 299.615 ;
        RECT 70.740 299.845 71.360 300.030 ;
        RECT 102.340 299.845 102.960 300.030 ;
        RECT 70.740 299.615 102.960 299.845 ;
        RECT 70.740 299.430 71.360 299.615 ;
        RECT 102.340 299.430 102.960 299.615 ;
        RECT 103.190 299.845 103.810 300.030 ;
        RECT 134.790 299.845 135.410 300.030 ;
        RECT 103.190 299.615 135.410 299.845 ;
        RECT 103.190 299.430 103.810 299.615 ;
        RECT 134.790 299.430 135.410 299.615 ;
        RECT 6.690 298.980 37.210 299.350 ;
        RECT 39.140 298.980 69.660 299.350 ;
        RECT 71.590 298.980 102.110 299.350 ;
        RECT 104.040 298.980 134.560 299.350 ;
        RECT 0.960 297.650 3.025 297.880 ;
        RECT 3.255 297.650 4.650 297.880 ;
        RECT 4.050 297.015 4.650 297.650 ;
        RECT 0.130 296.675 2.420 297.015 ;
        RECT 3.165 296.675 4.650 297.015 ;
        RECT 0.130 296.040 0.730 296.675 ;
        RECT 0.130 295.810 1.710 296.040 ;
        RECT 0.130 293.770 0.730 295.810 ;
        RECT 2.140 295.580 2.500 295.665 ;
        RECT 1.010 295.350 2.500 295.580 ;
        RECT 1.010 295.200 1.370 295.350 ;
        RECT 0.960 294.565 1.910 294.970 ;
        RECT 0.130 293.540 1.420 293.770 ;
        RECT 0.130 292.580 0.730 293.540 ;
        RECT 1.650 293.220 1.910 294.565 ;
        RECT 2.140 293.915 2.500 295.350 ;
        RECT 2.730 294.015 3.080 295.215 ;
        RECT 3.440 294.605 3.820 296.250 ;
        RECT 2.520 293.220 2.870 293.280 ;
        RECT 3.440 293.220 3.780 293.825 ;
        RECT 1.650 292.960 3.780 293.220 ;
        RECT 2.520 292.900 2.870 292.960 ;
        RECT 4.050 292.680 4.650 296.675 ;
        RECT 6.495 296.195 8.245 298.980 ;
        RECT 8.885 296.195 9.695 297.195 ;
        RECT 10.335 296.195 12.085 298.490 ;
        RECT 12.725 296.195 13.535 297.195 ;
        RECT 14.175 296.195 15.925 298.490 ;
        RECT 16.565 296.195 17.375 297.195 ;
        RECT 18.015 296.195 19.765 298.490 ;
        RECT 20.405 296.195 21.215 297.195 ;
        RECT 21.855 296.195 23.605 298.490 ;
        RECT 24.245 296.195 25.055 297.195 ;
        RECT 25.695 296.195 27.445 298.490 ;
        RECT 28.085 296.195 28.895 297.195 ;
        RECT 29.535 296.195 31.285 298.490 ;
        RECT 31.925 296.195 32.735 297.195 ;
        RECT 33.375 296.195 35.125 298.490 ;
        RECT 35.765 296.195 36.575 297.195 ;
        RECT 38.945 296.195 40.695 298.980 ;
        RECT 41.335 296.195 42.145 297.195 ;
        RECT 42.785 296.195 44.535 298.490 ;
        RECT 45.175 296.195 45.985 297.195 ;
        RECT 46.625 296.195 48.375 298.490 ;
        RECT 49.015 296.195 49.825 297.195 ;
        RECT 50.465 296.195 52.215 298.490 ;
        RECT 52.855 296.195 53.665 297.195 ;
        RECT 54.305 296.195 56.055 298.490 ;
        RECT 56.695 296.195 57.505 297.195 ;
        RECT 58.145 296.195 59.895 298.490 ;
        RECT 60.535 296.195 61.345 297.195 ;
        RECT 61.985 296.195 63.735 298.490 ;
        RECT 64.375 296.195 65.185 297.195 ;
        RECT 65.825 296.195 67.575 298.490 ;
        RECT 68.215 296.195 69.025 297.195 ;
        RECT 71.395 296.195 73.145 298.980 ;
        RECT 73.785 296.195 74.595 297.195 ;
        RECT 75.235 296.195 76.985 298.490 ;
        RECT 77.625 296.195 78.435 297.195 ;
        RECT 79.075 296.195 80.825 298.490 ;
        RECT 81.465 296.195 82.275 297.195 ;
        RECT 82.915 296.195 84.665 298.490 ;
        RECT 85.305 296.195 86.115 297.195 ;
        RECT 86.755 296.195 88.505 298.490 ;
        RECT 89.145 296.195 89.955 297.195 ;
        RECT 90.595 296.195 92.345 298.490 ;
        RECT 92.985 296.195 93.795 297.195 ;
        RECT 94.435 296.195 96.185 298.490 ;
        RECT 96.825 296.195 97.635 297.195 ;
        RECT 98.275 296.195 100.025 298.490 ;
        RECT 100.665 296.195 101.475 297.195 ;
        RECT 103.845 296.195 105.595 298.980 ;
        RECT 106.235 296.195 107.045 297.195 ;
        RECT 107.685 296.195 109.435 298.490 ;
        RECT 110.075 296.195 110.885 297.195 ;
        RECT 111.525 296.195 113.275 298.490 ;
        RECT 113.915 296.195 114.725 297.195 ;
        RECT 115.365 296.195 117.115 298.490 ;
        RECT 117.755 296.195 118.565 297.195 ;
        RECT 119.205 296.195 120.955 298.490 ;
        RECT 121.595 296.195 122.405 297.195 ;
        RECT 123.045 296.195 124.795 298.490 ;
        RECT 125.435 296.195 126.245 297.195 ;
        RECT 126.885 296.195 128.635 298.490 ;
        RECT 129.275 296.195 130.085 297.195 ;
        RECT 130.725 296.195 132.475 298.490 ;
        RECT 133.115 296.195 133.925 297.195 ;
        RECT 136.340 296.385 136.710 314.895 ;
        RECT 137.360 311.260 137.730 314.895 ;
        RECT 137.355 310.880 137.735 311.260 ;
        RECT 137.360 308.260 137.730 310.880 ;
        RECT 137.355 307.880 137.735 308.260 ;
        RECT 137.360 305.260 137.730 307.880 ;
        RECT 137.355 304.880 137.735 305.260 ;
        RECT 137.360 302.260 137.730 304.880 ;
        RECT 137.355 301.880 137.735 302.260 ;
        RECT 137.360 299.260 137.730 301.880 ;
        RECT 137.355 298.880 137.735 299.260 ;
        RECT 136.340 296.005 136.720 296.385 ;
        RECT 136.340 294.935 136.710 296.005 ;
        RECT 6.965 293.745 7.775 294.745 ;
        RECT 0.130 292.350 1.820 292.580 ;
        RECT 3.190 292.450 4.650 292.680 ;
        RECT 0.130 290.340 0.730 292.350 ;
        RECT 2.150 291.890 3.150 292.215 ;
        RECT 0.960 291.330 3.820 291.660 ;
        RECT 0.130 290.110 1.820 290.340 ;
        RECT 0.130 288.100 0.730 290.110 ;
        RECT 2.535 289.975 2.800 291.330 ;
        RECT 4.050 290.440 4.650 292.450 ;
        RECT 8.415 291.915 10.165 294.745 ;
        RECT 10.805 293.745 11.615 294.745 ;
        RECT 12.255 292.450 14.005 294.745 ;
        RECT 14.645 293.745 15.455 294.745 ;
        RECT 16.095 292.450 17.845 294.745 ;
        RECT 18.485 293.745 19.295 294.745 ;
        RECT 19.935 292.450 21.685 294.745 ;
        RECT 22.325 293.745 23.135 294.745 ;
        RECT 23.775 292.450 25.525 294.745 ;
        RECT 26.165 293.745 26.975 294.745 ;
        RECT 27.615 292.450 29.365 294.745 ;
        RECT 30.005 293.745 30.815 294.745 ;
        RECT 31.455 292.450 33.205 294.745 ;
        RECT 33.845 293.745 34.655 294.745 ;
        RECT 35.295 292.450 37.045 294.745 ;
        RECT 39.415 293.745 40.225 294.745 ;
        RECT 40.865 291.915 42.615 294.745 ;
        RECT 43.255 293.745 44.065 294.745 ;
        RECT 44.705 292.450 46.455 294.745 ;
        RECT 47.095 293.745 47.905 294.745 ;
        RECT 48.545 292.450 50.295 294.745 ;
        RECT 50.935 293.745 51.745 294.745 ;
        RECT 52.385 292.450 54.135 294.745 ;
        RECT 54.775 293.745 55.585 294.745 ;
        RECT 56.225 292.450 57.975 294.745 ;
        RECT 58.615 293.745 59.425 294.745 ;
        RECT 60.065 292.450 61.815 294.745 ;
        RECT 62.455 293.745 63.265 294.745 ;
        RECT 63.905 292.450 65.655 294.745 ;
        RECT 66.295 293.745 67.105 294.745 ;
        RECT 67.745 292.450 69.495 294.745 ;
        RECT 71.865 293.745 72.675 294.745 ;
        RECT 73.315 291.915 75.065 294.745 ;
        RECT 75.705 293.745 76.515 294.745 ;
        RECT 77.155 292.450 78.905 294.745 ;
        RECT 79.545 293.745 80.355 294.745 ;
        RECT 80.995 292.450 82.745 294.745 ;
        RECT 83.385 293.745 84.195 294.745 ;
        RECT 84.835 292.450 86.585 294.745 ;
        RECT 87.225 293.745 88.035 294.745 ;
        RECT 88.675 292.450 90.425 294.745 ;
        RECT 91.065 293.745 91.875 294.745 ;
        RECT 92.515 292.450 94.265 294.745 ;
        RECT 94.905 293.745 95.715 294.745 ;
        RECT 96.355 292.450 98.105 294.745 ;
        RECT 98.745 293.745 99.555 294.745 ;
        RECT 100.195 292.450 101.945 294.745 ;
        RECT 104.315 293.745 105.125 294.745 ;
        RECT 105.765 291.915 107.515 294.745 ;
        RECT 108.155 293.745 108.965 294.745 ;
        RECT 109.605 292.450 111.355 294.745 ;
        RECT 111.995 293.745 112.805 294.745 ;
        RECT 113.445 292.450 115.195 294.745 ;
        RECT 115.835 293.745 116.645 294.745 ;
        RECT 117.285 292.450 119.035 294.745 ;
        RECT 119.675 293.745 120.485 294.745 ;
        RECT 121.125 292.450 122.875 294.745 ;
        RECT 123.515 293.745 124.325 294.745 ;
        RECT 124.965 292.450 126.715 294.745 ;
        RECT 127.355 293.745 128.165 294.745 ;
        RECT 128.805 292.450 130.555 294.745 ;
        RECT 131.195 293.745 132.005 294.745 ;
        RECT 132.645 292.450 134.395 294.745 ;
        RECT 136.340 294.555 136.720 294.935 ;
        RECT 6.690 291.545 37.210 291.915 ;
        RECT 39.140 291.545 69.660 291.915 ;
        RECT 71.590 291.545 102.110 291.915 ;
        RECT 104.040 291.545 134.560 291.915 ;
        RECT 5.840 291.280 6.460 291.465 ;
        RECT 37.440 291.280 38.060 291.465 ;
        RECT 5.840 291.050 38.060 291.280 ;
        RECT 5.840 290.865 6.460 291.050 ;
        RECT 37.440 290.865 38.060 291.050 ;
        RECT 38.290 291.280 38.910 291.465 ;
        RECT 69.890 291.280 70.510 291.465 ;
        RECT 38.290 291.050 70.510 291.280 ;
        RECT 38.290 290.865 38.910 291.050 ;
        RECT 69.890 290.865 70.510 291.050 ;
        RECT 70.740 291.280 71.360 291.465 ;
        RECT 102.340 291.280 102.960 291.465 ;
        RECT 70.740 291.050 102.960 291.280 ;
        RECT 70.740 290.865 71.360 291.050 ;
        RECT 102.340 290.865 102.960 291.050 ;
        RECT 103.190 291.280 103.810 291.465 ;
        RECT 134.790 291.280 135.410 291.465 ;
        RECT 103.190 291.050 135.410 291.280 ;
        RECT 103.190 290.865 103.810 291.050 ;
        RECT 134.790 290.865 135.410 291.050 ;
        RECT 3.190 290.210 4.650 290.440 ;
        RECT 6.690 290.415 37.210 290.795 ;
        RECT 39.140 290.415 69.660 290.795 ;
        RECT 71.590 290.415 102.110 290.795 ;
        RECT 104.040 290.415 134.560 290.795 ;
        RECT 2.150 289.650 3.150 289.975 ;
        RECT 0.960 289.090 3.820 289.420 ;
        RECT 4.050 288.200 4.650 290.210 ;
        RECT 6.690 289.705 37.210 290.075 ;
        RECT 39.140 289.705 69.660 290.075 ;
        RECT 71.590 289.705 102.110 290.075 ;
        RECT 104.040 289.705 134.560 290.075 ;
        RECT 12.320 289.695 13.940 289.705 ;
        RECT 44.770 289.695 46.390 289.705 ;
        RECT 77.220 289.695 78.840 289.705 ;
        RECT 109.670 289.695 111.290 289.705 ;
        RECT 5.840 289.440 6.460 289.625 ;
        RECT 37.440 289.440 38.060 289.625 ;
        RECT 5.840 289.210 38.060 289.440 ;
        RECT 5.840 289.025 6.460 289.210 ;
        RECT 37.440 289.025 38.060 289.210 ;
        RECT 38.290 289.440 38.910 289.625 ;
        RECT 69.890 289.440 70.510 289.625 ;
        RECT 38.290 289.210 70.510 289.440 ;
        RECT 38.290 289.025 38.910 289.210 ;
        RECT 69.890 289.025 70.510 289.210 ;
        RECT 70.740 289.440 71.360 289.625 ;
        RECT 102.340 289.440 102.960 289.625 ;
        RECT 70.740 289.210 102.960 289.440 ;
        RECT 70.740 289.025 71.360 289.210 ;
        RECT 102.340 289.025 102.960 289.210 ;
        RECT 103.190 289.440 103.810 289.625 ;
        RECT 134.790 289.440 135.410 289.625 ;
        RECT 103.190 289.210 135.410 289.440 ;
        RECT 103.190 289.025 103.810 289.210 ;
        RECT 134.790 289.025 135.410 289.210 ;
        RECT 6.690 288.575 37.210 288.955 ;
        RECT 39.140 288.575 69.660 288.955 ;
        RECT 71.590 288.575 102.110 288.955 ;
        RECT 104.040 288.575 134.560 288.955 ;
        RECT 0.130 287.870 1.820 288.100 ;
        RECT 3.190 287.970 4.650 288.200 ;
        RECT 0.130 285.815 0.730 287.870 ;
        RECT 2.150 287.410 3.150 287.735 ;
        RECT 0.960 286.850 3.820 287.180 ;
        RECT 2.300 286.725 2.680 286.850 ;
        RECT 4.050 285.815 4.650 287.970 ;
        RECT 6.690 287.860 37.210 288.230 ;
        RECT 39.140 287.860 69.660 288.230 ;
        RECT 71.590 287.860 102.110 288.230 ;
        RECT 104.040 287.860 134.560 288.230 ;
        RECT 16.160 287.850 17.780 287.860 ;
        RECT 48.610 287.850 50.230 287.860 ;
        RECT 81.060 287.850 82.680 287.860 ;
        RECT 113.510 287.850 115.130 287.860 ;
        RECT 5.840 287.595 6.460 287.780 ;
        RECT 37.440 287.595 38.060 287.780 ;
        RECT 5.840 287.365 38.060 287.595 ;
        RECT 5.840 287.180 6.460 287.365 ;
        RECT 37.440 287.180 38.060 287.365 ;
        RECT 38.290 287.595 38.910 287.780 ;
        RECT 69.890 287.595 70.510 287.780 ;
        RECT 38.290 287.365 70.510 287.595 ;
        RECT 38.290 287.180 38.910 287.365 ;
        RECT 69.890 287.180 70.510 287.365 ;
        RECT 70.740 287.595 71.360 287.780 ;
        RECT 102.340 287.595 102.960 287.780 ;
        RECT 70.740 287.365 102.960 287.595 ;
        RECT 70.740 287.180 71.360 287.365 ;
        RECT 102.340 287.180 102.960 287.365 ;
        RECT 103.190 287.595 103.810 287.780 ;
        RECT 134.790 287.595 135.410 287.780 ;
        RECT 103.190 287.365 135.410 287.595 ;
        RECT 103.190 287.180 103.810 287.365 ;
        RECT 134.790 287.180 135.410 287.365 ;
        RECT 6.690 286.730 37.210 287.110 ;
        RECT 39.140 286.730 69.660 287.110 ;
        RECT 71.590 286.730 102.110 287.110 ;
        RECT 104.040 286.730 134.560 287.110 ;
        RECT 6.700 285.940 37.200 286.380 ;
        RECT 39.150 285.940 69.650 286.380 ;
        RECT 71.600 285.940 102.100 286.380 ;
        RECT 104.050 285.940 134.550 286.380 ;
        RECT 0.130 285.475 2.420 285.815 ;
        RECT 3.165 285.475 4.650 285.815 ;
        RECT 0.130 284.695 0.730 285.475 ;
        RECT 4.050 284.695 4.650 285.475 ;
        RECT 6.690 285.220 37.210 285.590 ;
        RECT 39.140 285.220 69.660 285.590 ;
        RECT 71.590 285.220 102.110 285.590 ;
        RECT 104.040 285.220 134.560 285.590 ;
        RECT 20.000 285.210 21.620 285.220 ;
        RECT 52.450 285.210 54.070 285.220 ;
        RECT 84.900 285.210 86.520 285.220 ;
        RECT 117.350 285.210 118.970 285.220 ;
        RECT 0.130 284.355 2.420 284.695 ;
        RECT 3.165 284.355 4.650 284.695 ;
        RECT 5.840 284.955 6.460 285.140 ;
        RECT 37.440 284.955 38.060 285.140 ;
        RECT 5.840 284.725 38.060 284.955 ;
        RECT 5.840 284.540 6.460 284.725 ;
        RECT 37.440 284.540 38.060 284.725 ;
        RECT 38.290 284.955 38.910 285.140 ;
        RECT 69.890 284.955 70.510 285.140 ;
        RECT 38.290 284.725 70.510 284.955 ;
        RECT 38.290 284.540 38.910 284.725 ;
        RECT 69.890 284.540 70.510 284.725 ;
        RECT 70.740 284.955 71.360 285.140 ;
        RECT 102.340 284.955 102.960 285.140 ;
        RECT 70.740 284.725 102.960 284.955 ;
        RECT 70.740 284.540 71.360 284.725 ;
        RECT 102.340 284.540 102.960 284.725 ;
        RECT 103.190 284.955 103.810 285.140 ;
        RECT 134.790 284.955 135.410 285.140 ;
        RECT 103.190 284.725 135.410 284.955 ;
        RECT 103.190 284.540 103.810 284.725 ;
        RECT 134.790 284.540 135.410 284.725 ;
        RECT 0.130 283.720 0.730 284.355 ;
        RECT 0.130 283.490 1.860 283.720 ;
        RECT 2.160 283.490 3.820 283.720 ;
        RECT 0.130 281.480 0.730 283.490 ;
        RECT 2.160 282.455 2.390 283.490 ;
        RECT 2.795 282.200 3.025 283.245 ;
        RECT 4.050 282.200 4.650 284.355 ;
        RECT 6.690 284.090 37.210 284.470 ;
        RECT 39.140 284.090 69.660 284.470 ;
        RECT 71.590 284.090 102.110 284.470 ;
        RECT 104.040 284.090 134.560 284.470 ;
        RECT 6.690 283.380 37.210 283.750 ;
        RECT 39.140 283.380 69.660 283.750 ;
        RECT 71.590 283.380 102.110 283.750 ;
        RECT 104.040 283.380 134.560 283.750 ;
        RECT 23.840 283.370 25.460 283.380 ;
        RECT 56.290 283.370 57.910 283.380 ;
        RECT 88.740 283.370 90.360 283.380 ;
        RECT 121.190 283.370 122.810 283.380 ;
        RECT 5.840 283.115 6.460 283.300 ;
        RECT 37.440 283.115 38.060 283.300 ;
        RECT 5.840 282.885 38.060 283.115 ;
        RECT 5.840 282.700 6.460 282.885 ;
        RECT 37.440 282.700 38.060 282.885 ;
        RECT 38.290 283.115 38.910 283.300 ;
        RECT 69.890 283.115 70.510 283.300 ;
        RECT 38.290 282.885 70.510 283.115 ;
        RECT 38.290 282.700 38.910 282.885 ;
        RECT 69.890 282.700 70.510 282.885 ;
        RECT 70.740 283.115 71.360 283.300 ;
        RECT 102.340 283.115 102.960 283.300 ;
        RECT 70.740 282.885 102.960 283.115 ;
        RECT 70.740 282.700 71.360 282.885 ;
        RECT 102.340 282.700 102.960 282.885 ;
        RECT 103.190 283.115 103.810 283.300 ;
        RECT 134.790 283.115 135.410 283.300 ;
        RECT 103.190 282.885 135.410 283.115 ;
        RECT 103.190 282.700 103.810 282.885 ;
        RECT 134.790 282.700 135.410 282.885 ;
        RECT 6.690 282.250 37.210 282.630 ;
        RECT 39.140 282.250 69.660 282.630 ;
        RECT 71.590 282.250 102.110 282.630 ;
        RECT 104.040 282.250 134.560 282.630 ;
        RECT 0.960 281.970 3.025 282.200 ;
        RECT 3.255 281.970 4.650 282.200 ;
        RECT 0.130 281.250 1.860 281.480 ;
        RECT 2.160 281.250 3.820 281.480 ;
        RECT 0.130 279.240 0.730 281.250 ;
        RECT 2.160 280.215 2.390 281.250 ;
        RECT 2.795 279.960 3.025 281.005 ;
        RECT 4.050 279.960 4.650 281.970 ;
        RECT 6.690 281.535 37.210 281.905 ;
        RECT 39.140 281.535 69.660 281.905 ;
        RECT 71.590 281.535 102.110 281.905 ;
        RECT 104.040 281.535 134.560 281.905 ;
        RECT 27.680 281.525 29.300 281.535 ;
        RECT 60.130 281.525 61.750 281.535 ;
        RECT 92.580 281.525 94.200 281.535 ;
        RECT 125.030 281.525 126.650 281.535 ;
        RECT 5.840 281.270 6.460 281.455 ;
        RECT 37.440 281.270 38.060 281.455 ;
        RECT 5.840 281.040 38.060 281.270 ;
        RECT 5.840 280.855 6.460 281.040 ;
        RECT 37.440 280.855 38.060 281.040 ;
        RECT 38.290 281.270 38.910 281.455 ;
        RECT 69.890 281.270 70.510 281.455 ;
        RECT 38.290 281.040 70.510 281.270 ;
        RECT 38.290 280.855 38.910 281.040 ;
        RECT 69.890 280.855 70.510 281.040 ;
        RECT 70.740 281.270 71.360 281.455 ;
        RECT 102.340 281.270 102.960 281.455 ;
        RECT 70.740 281.040 102.960 281.270 ;
        RECT 70.740 280.855 71.360 281.040 ;
        RECT 102.340 280.855 102.960 281.040 ;
        RECT 103.190 281.270 103.810 281.455 ;
        RECT 134.790 281.270 135.410 281.455 ;
        RECT 103.190 281.040 135.410 281.270 ;
        RECT 103.190 280.855 103.810 281.040 ;
        RECT 134.790 280.855 135.410 281.040 ;
        RECT 6.690 280.405 37.210 280.785 ;
        RECT 39.140 280.405 69.660 280.785 ;
        RECT 71.590 280.405 102.110 280.785 ;
        RECT 104.040 280.405 134.560 280.785 ;
        RECT 0.960 279.730 3.025 279.960 ;
        RECT 3.255 279.730 4.650 279.960 ;
        RECT 0.130 279.010 1.860 279.240 ;
        RECT 2.160 279.010 3.820 279.240 ;
        RECT 0.130 276.835 0.730 279.010 ;
        RECT 2.160 277.975 2.390 279.010 ;
        RECT 2.795 277.720 3.025 278.765 ;
        RECT 4.050 277.720 4.650 279.730 ;
        RECT 6.700 279.615 37.200 280.055 ;
        RECT 39.150 279.615 69.650 280.055 ;
        RECT 71.600 279.615 102.100 280.055 ;
        RECT 104.050 279.615 134.550 280.055 ;
        RECT 6.690 278.895 37.210 279.265 ;
        RECT 39.140 278.895 69.660 279.265 ;
        RECT 71.590 278.895 102.110 279.265 ;
        RECT 104.040 278.895 134.560 279.265 ;
        RECT 31.520 278.885 33.140 278.895 ;
        RECT 63.970 278.885 65.590 278.895 ;
        RECT 96.420 278.885 98.040 278.895 ;
        RECT 128.870 278.885 130.490 278.895 ;
        RECT 5.840 278.630 6.460 278.815 ;
        RECT 37.440 278.630 38.060 278.815 ;
        RECT 5.840 278.400 38.060 278.630 ;
        RECT 5.840 278.215 6.460 278.400 ;
        RECT 37.440 278.215 38.060 278.400 ;
        RECT 38.290 278.630 38.910 278.815 ;
        RECT 69.890 278.630 70.510 278.815 ;
        RECT 38.290 278.400 70.510 278.630 ;
        RECT 38.290 278.215 38.910 278.400 ;
        RECT 69.890 278.215 70.510 278.400 ;
        RECT 70.740 278.630 71.360 278.815 ;
        RECT 102.340 278.630 102.960 278.815 ;
        RECT 70.740 278.400 102.960 278.630 ;
        RECT 70.740 278.215 71.360 278.400 ;
        RECT 102.340 278.215 102.960 278.400 ;
        RECT 103.190 278.630 103.810 278.815 ;
        RECT 134.790 278.630 135.410 278.815 ;
        RECT 103.190 278.400 135.410 278.630 ;
        RECT 103.190 278.215 103.810 278.400 ;
        RECT 134.790 278.215 135.410 278.400 ;
        RECT 6.690 277.765 37.210 278.145 ;
        RECT 39.140 277.765 69.660 278.145 ;
        RECT 71.590 277.765 102.110 278.145 ;
        RECT 104.040 277.765 134.560 278.145 ;
        RECT 0.960 277.490 3.025 277.720 ;
        RECT 3.255 277.490 4.650 277.720 ;
        RECT 4.050 276.835 4.650 277.490 ;
        RECT 6.690 277.055 37.210 277.425 ;
        RECT 39.140 277.055 69.660 277.425 ;
        RECT 71.590 277.055 102.110 277.425 ;
        RECT 104.040 277.055 134.560 277.425 ;
        RECT 35.360 277.045 36.980 277.055 ;
        RECT 67.810 277.045 69.430 277.055 ;
        RECT 100.260 277.045 101.880 277.055 ;
        RECT 132.710 277.045 134.330 277.055 ;
        RECT 0.130 276.495 2.430 276.835 ;
        RECT 3.160 276.495 4.650 276.835 ;
        RECT 0.130 275.530 0.730 276.495 ;
        RECT 4.050 275.530 4.650 276.495 ;
        RECT 5.840 276.790 6.460 276.975 ;
        RECT 37.440 276.790 38.060 276.975 ;
        RECT 5.840 276.560 38.060 276.790 ;
        RECT 5.840 276.375 6.460 276.560 ;
        RECT 37.440 276.375 38.060 276.560 ;
        RECT 38.290 276.790 38.910 276.975 ;
        RECT 69.890 276.790 70.510 276.975 ;
        RECT 38.290 276.560 70.510 276.790 ;
        RECT 38.290 276.375 38.910 276.560 ;
        RECT 69.890 276.375 70.510 276.560 ;
        RECT 70.740 276.790 71.360 276.975 ;
        RECT 102.340 276.790 102.960 276.975 ;
        RECT 70.740 276.560 102.960 276.790 ;
        RECT 70.740 276.375 71.360 276.560 ;
        RECT 102.340 276.375 102.960 276.560 ;
        RECT 103.190 276.790 103.810 276.975 ;
        RECT 134.790 276.790 135.410 276.975 ;
        RECT 103.190 276.560 135.410 276.790 ;
        RECT 136.340 276.625 136.710 294.555 ;
        RECT 137.360 293.260 137.730 298.880 ;
        RECT 138.380 296.385 138.750 314.895 ;
        RECT 139.400 311.260 139.770 314.895 ;
        RECT 139.395 310.880 139.775 311.260 ;
        RECT 139.400 308.260 139.770 310.880 ;
        RECT 139.395 307.880 139.775 308.260 ;
        RECT 139.400 305.260 139.770 307.880 ;
        RECT 139.395 304.880 139.775 305.260 ;
        RECT 139.400 302.260 139.770 304.880 ;
        RECT 139.395 301.880 139.775 302.260 ;
        RECT 139.400 299.260 139.770 301.880 ;
        RECT 139.395 298.880 139.775 299.260 ;
        RECT 138.380 296.005 138.760 296.385 ;
        RECT 138.380 294.935 138.750 296.005 ;
        RECT 138.380 294.555 138.760 294.935 ;
        RECT 137.355 292.880 137.735 293.260 ;
        RECT 137.360 290.260 137.730 292.880 ;
        RECT 137.355 289.880 137.735 290.260 ;
        RECT 137.360 287.260 137.730 289.880 ;
        RECT 137.355 286.880 137.735 287.260 ;
        RECT 137.360 284.260 137.730 286.880 ;
        RECT 137.355 283.880 137.735 284.260 ;
        RECT 137.360 281.260 137.730 283.880 ;
        RECT 137.355 280.880 137.735 281.260 ;
        RECT 137.360 278.260 137.730 280.880 ;
        RECT 137.355 277.880 137.735 278.260 ;
        RECT 137.360 276.625 137.730 277.880 ;
        RECT 138.380 276.625 138.750 294.555 ;
        RECT 139.400 293.260 139.770 298.880 ;
        RECT 139.395 292.880 139.775 293.260 ;
        RECT 139.400 290.260 139.770 292.880 ;
        RECT 139.395 289.880 139.775 290.260 ;
        RECT 139.400 287.260 139.770 289.880 ;
        RECT 139.395 286.880 139.775 287.260 ;
        RECT 139.400 284.260 139.770 286.880 ;
        RECT 139.395 283.880 139.775 284.260 ;
        RECT 139.400 281.260 139.770 283.880 ;
        RECT 139.395 280.880 139.775 281.260 ;
        RECT 139.400 278.260 139.770 280.880 ;
        RECT 139.395 277.880 139.775 278.260 ;
        RECT 139.400 276.625 139.770 277.880 ;
        RECT 140.420 276.625 140.800 314.895 ;
        RECT 141.150 276.635 141.590 314.885 ;
        RECT 103.190 276.375 103.810 276.560 ;
        RECT 134.790 276.375 135.410 276.560 ;
        RECT 6.690 275.925 37.210 276.305 ;
        RECT 39.140 275.925 69.660 276.305 ;
        RECT 71.590 275.925 102.110 276.305 ;
        RECT 104.040 275.925 134.560 276.305 ;
        RECT 0.130 275.190 2.430 275.530 ;
        RECT 3.160 275.190 4.650 275.530 ;
        RECT 6.690 275.205 37.210 275.585 ;
        RECT 39.140 275.205 69.660 275.585 ;
        RECT 71.590 275.205 102.110 275.585 ;
        RECT 104.040 275.205 134.560 275.585 ;
        RECT 0.130 274.575 0.730 275.190 ;
        RECT 0.130 274.345 1.860 274.575 ;
        RECT 2.160 274.345 3.820 274.575 ;
        RECT 0.130 272.335 0.730 274.345 ;
        RECT 2.160 273.310 2.390 274.345 ;
        RECT 2.795 273.055 3.025 274.100 ;
        RECT 4.050 273.055 4.650 275.190 ;
        RECT 5.840 274.950 6.460 275.135 ;
        RECT 37.440 274.950 38.060 275.135 ;
        RECT 5.840 274.720 38.060 274.950 ;
        RECT 5.840 274.535 6.460 274.720 ;
        RECT 37.440 274.535 38.060 274.720 ;
        RECT 38.290 274.950 38.910 275.135 ;
        RECT 69.890 274.950 70.510 275.135 ;
        RECT 38.290 274.720 70.510 274.950 ;
        RECT 38.290 274.535 38.910 274.720 ;
        RECT 69.890 274.535 70.510 274.720 ;
        RECT 70.740 274.950 71.360 275.135 ;
        RECT 102.340 274.950 102.960 275.135 ;
        RECT 70.740 274.720 102.960 274.950 ;
        RECT 70.740 274.535 71.360 274.720 ;
        RECT 102.340 274.535 102.960 274.720 ;
        RECT 103.190 274.950 103.810 275.135 ;
        RECT 134.790 274.950 135.410 275.135 ;
        RECT 103.190 274.720 135.410 274.950 ;
        RECT 103.190 274.535 103.810 274.720 ;
        RECT 134.790 274.535 135.410 274.720 ;
        RECT 33.440 274.455 35.060 274.465 ;
        RECT 65.890 274.455 67.510 274.465 ;
        RECT 98.340 274.455 99.960 274.465 ;
        RECT 130.790 274.455 132.410 274.465 ;
        RECT 6.690 274.085 37.210 274.455 ;
        RECT 39.140 274.085 69.660 274.455 ;
        RECT 71.590 274.085 102.110 274.455 ;
        RECT 104.040 274.085 134.560 274.455 ;
        RECT 6.690 273.365 37.210 273.745 ;
        RECT 39.140 273.365 69.660 273.745 ;
        RECT 71.590 273.365 102.110 273.745 ;
        RECT 104.040 273.365 134.560 273.745 ;
        RECT 0.960 272.825 3.025 273.055 ;
        RECT 3.255 272.825 4.650 273.055 ;
        RECT 0.130 272.105 1.860 272.335 ;
        RECT 2.160 272.105 3.820 272.335 ;
        RECT 0.130 270.095 0.730 272.105 ;
        RECT 2.160 271.070 2.390 272.105 ;
        RECT 2.795 270.815 3.025 271.860 ;
        RECT 4.050 270.815 4.650 272.825 ;
        RECT 5.840 273.110 6.460 273.295 ;
        RECT 37.440 273.110 38.060 273.295 ;
        RECT 5.840 272.880 38.060 273.110 ;
        RECT 5.840 272.695 6.460 272.880 ;
        RECT 37.440 272.695 38.060 272.880 ;
        RECT 38.290 273.110 38.910 273.295 ;
        RECT 69.890 273.110 70.510 273.295 ;
        RECT 38.290 272.880 70.510 273.110 ;
        RECT 38.290 272.695 38.910 272.880 ;
        RECT 69.890 272.695 70.510 272.880 ;
        RECT 70.740 273.110 71.360 273.295 ;
        RECT 102.340 273.110 102.960 273.295 ;
        RECT 70.740 272.880 102.960 273.110 ;
        RECT 70.740 272.695 71.360 272.880 ;
        RECT 102.340 272.695 102.960 272.880 ;
        RECT 103.190 273.110 103.810 273.295 ;
        RECT 134.790 273.110 135.410 273.295 ;
        RECT 103.190 272.880 135.410 273.110 ;
        RECT 103.190 272.695 103.810 272.880 ;
        RECT 134.790 272.695 135.410 272.880 ;
        RECT 29.600 272.615 31.220 272.625 ;
        RECT 62.050 272.615 63.670 272.625 ;
        RECT 94.500 272.615 96.120 272.625 ;
        RECT 126.950 272.615 128.570 272.625 ;
        RECT 6.690 272.245 37.210 272.615 ;
        RECT 39.140 272.245 69.660 272.615 ;
        RECT 71.590 272.245 102.110 272.615 ;
        RECT 104.040 272.245 134.560 272.615 ;
        RECT 6.700 271.450 37.200 271.890 ;
        RECT 39.150 271.450 69.650 271.890 ;
        RECT 71.600 271.450 102.100 271.890 ;
        RECT 104.050 271.450 134.550 271.890 ;
        RECT 0.960 270.585 3.025 270.815 ;
        RECT 3.255 270.585 4.650 270.815 ;
        RECT 6.690 270.720 37.210 271.100 ;
        RECT 39.140 270.720 69.660 271.100 ;
        RECT 71.590 270.720 102.110 271.100 ;
        RECT 104.040 270.720 134.560 271.100 ;
        RECT 0.130 269.865 1.860 270.095 ;
        RECT 2.160 269.865 3.820 270.095 ;
        RECT 0.130 267.855 0.730 269.865 ;
        RECT 2.160 268.830 2.390 269.865 ;
        RECT 2.795 268.575 3.025 269.620 ;
        RECT 4.050 268.575 4.650 270.585 ;
        RECT 5.840 270.465 6.460 270.650 ;
        RECT 37.440 270.465 38.060 270.650 ;
        RECT 5.840 270.235 38.060 270.465 ;
        RECT 5.840 270.050 6.460 270.235 ;
        RECT 37.440 270.050 38.060 270.235 ;
        RECT 38.290 270.465 38.910 270.650 ;
        RECT 69.890 270.465 70.510 270.650 ;
        RECT 38.290 270.235 70.510 270.465 ;
        RECT 38.290 270.050 38.910 270.235 ;
        RECT 69.890 270.050 70.510 270.235 ;
        RECT 70.740 270.465 71.360 270.650 ;
        RECT 102.340 270.465 102.960 270.650 ;
        RECT 70.740 270.235 102.960 270.465 ;
        RECT 70.740 270.050 71.360 270.235 ;
        RECT 102.340 270.050 102.960 270.235 ;
        RECT 103.190 270.465 103.810 270.650 ;
        RECT 134.790 270.465 135.410 270.650 ;
        RECT 103.190 270.235 135.410 270.465 ;
        RECT 103.190 270.050 103.810 270.235 ;
        RECT 134.790 270.050 135.410 270.235 ;
        RECT 25.760 269.970 27.380 269.980 ;
        RECT 58.210 269.970 59.830 269.980 ;
        RECT 90.660 269.970 92.280 269.980 ;
        RECT 123.110 269.970 124.730 269.980 ;
        RECT 6.690 269.600 37.210 269.970 ;
        RECT 39.140 269.600 69.660 269.970 ;
        RECT 71.590 269.600 102.110 269.970 ;
        RECT 104.040 269.600 134.560 269.970 ;
        RECT 6.690 268.880 37.210 269.260 ;
        RECT 39.140 268.880 69.660 269.260 ;
        RECT 71.590 268.880 102.110 269.260 ;
        RECT 104.040 268.880 134.560 269.260 ;
        RECT 0.960 268.345 3.025 268.575 ;
        RECT 3.255 268.345 4.650 268.575 ;
        RECT 0.130 267.625 1.860 267.855 ;
        RECT 2.160 267.625 3.820 267.855 ;
        RECT 0.130 265.615 0.730 267.625 ;
        RECT 2.160 266.590 2.390 267.625 ;
        RECT 2.795 266.335 3.025 267.380 ;
        RECT 4.050 266.335 4.650 268.345 ;
        RECT 5.840 268.625 6.460 268.810 ;
        RECT 37.440 268.625 38.060 268.810 ;
        RECT 5.840 268.395 38.060 268.625 ;
        RECT 5.840 268.210 6.460 268.395 ;
        RECT 37.440 268.210 38.060 268.395 ;
        RECT 38.290 268.625 38.910 268.810 ;
        RECT 69.890 268.625 70.510 268.810 ;
        RECT 38.290 268.395 70.510 268.625 ;
        RECT 38.290 268.210 38.910 268.395 ;
        RECT 69.890 268.210 70.510 268.395 ;
        RECT 70.740 268.625 71.360 268.810 ;
        RECT 102.340 268.625 102.960 268.810 ;
        RECT 70.740 268.395 102.960 268.625 ;
        RECT 70.740 268.210 71.360 268.395 ;
        RECT 102.340 268.210 102.960 268.395 ;
        RECT 103.190 268.625 103.810 268.810 ;
        RECT 134.790 268.625 135.410 268.810 ;
        RECT 103.190 268.395 135.410 268.625 ;
        RECT 103.190 268.210 103.810 268.395 ;
        RECT 134.790 268.210 135.410 268.395 ;
        RECT 21.920 268.130 23.540 268.140 ;
        RECT 54.370 268.130 55.990 268.140 ;
        RECT 86.820 268.130 88.440 268.140 ;
        RECT 119.270 268.130 120.890 268.140 ;
        RECT 6.690 267.760 37.210 268.130 ;
        RECT 39.140 267.760 69.660 268.130 ;
        RECT 71.590 267.760 102.110 268.130 ;
        RECT 104.040 267.760 134.560 268.130 ;
        RECT 6.690 267.040 37.210 267.420 ;
        RECT 39.140 267.040 69.660 267.420 ;
        RECT 71.590 267.040 102.110 267.420 ;
        RECT 104.040 267.040 134.560 267.420 ;
        RECT 5.840 266.785 6.460 266.970 ;
        RECT 37.440 266.785 38.060 266.970 ;
        RECT 5.840 266.555 38.060 266.785 ;
        RECT 5.840 266.370 6.460 266.555 ;
        RECT 37.440 266.370 38.060 266.555 ;
        RECT 38.290 266.785 38.910 266.970 ;
        RECT 69.890 266.785 70.510 266.970 ;
        RECT 38.290 266.555 70.510 266.785 ;
        RECT 38.290 266.370 38.910 266.555 ;
        RECT 69.890 266.370 70.510 266.555 ;
        RECT 70.740 266.785 71.360 266.970 ;
        RECT 102.340 266.785 102.960 266.970 ;
        RECT 70.740 266.555 102.960 266.785 ;
        RECT 70.740 266.370 71.360 266.555 ;
        RECT 102.340 266.370 102.960 266.555 ;
        RECT 103.190 266.785 103.810 266.970 ;
        RECT 134.790 266.785 135.410 266.970 ;
        RECT 103.190 266.555 135.410 266.785 ;
        RECT 103.190 266.370 103.810 266.555 ;
        RECT 134.790 266.370 135.410 266.555 ;
        RECT 0.960 266.105 3.025 266.335 ;
        RECT 3.255 266.105 4.650 266.335 ;
        RECT 18.080 266.290 19.700 266.300 ;
        RECT 50.530 266.290 52.150 266.300 ;
        RECT 82.980 266.290 84.600 266.300 ;
        RECT 115.430 266.290 117.050 266.300 ;
        RECT 0.130 265.385 1.860 265.615 ;
        RECT 2.160 265.385 3.820 265.615 ;
        RECT 0.130 263.230 0.730 265.385 ;
        RECT 2.160 264.350 2.390 265.385 ;
        RECT 2.795 264.095 3.025 265.140 ;
        RECT 4.050 264.095 4.650 266.105 ;
        RECT 6.690 265.920 37.210 266.290 ;
        RECT 39.140 265.920 69.660 266.290 ;
        RECT 71.590 265.920 102.110 266.290 ;
        RECT 104.040 265.920 134.560 266.290 ;
        RECT 6.700 265.125 37.200 265.565 ;
        RECT 39.150 265.125 69.650 265.565 ;
        RECT 71.600 265.125 102.100 265.565 ;
        RECT 104.050 265.125 134.550 265.565 ;
        RECT 6.690 264.395 37.210 264.775 ;
        RECT 39.140 264.395 69.660 264.775 ;
        RECT 71.590 264.395 102.110 264.775 ;
        RECT 104.040 264.395 134.560 264.775 ;
        RECT 0.960 263.865 3.025 264.095 ;
        RECT 3.255 263.865 4.650 264.095 ;
        RECT 4.050 263.230 4.650 263.865 ;
        RECT 5.840 264.140 6.460 264.325 ;
        RECT 37.440 264.140 38.060 264.325 ;
        RECT 5.840 263.910 38.060 264.140 ;
        RECT 5.840 263.725 6.460 263.910 ;
        RECT 37.440 263.725 38.060 263.910 ;
        RECT 38.290 264.140 38.910 264.325 ;
        RECT 69.890 264.140 70.510 264.325 ;
        RECT 38.290 263.910 70.510 264.140 ;
        RECT 38.290 263.725 38.910 263.910 ;
        RECT 69.890 263.725 70.510 263.910 ;
        RECT 70.740 264.140 71.360 264.325 ;
        RECT 102.340 264.140 102.960 264.325 ;
        RECT 70.740 263.910 102.960 264.140 ;
        RECT 70.740 263.725 71.360 263.910 ;
        RECT 102.340 263.725 102.960 263.910 ;
        RECT 103.190 264.140 103.810 264.325 ;
        RECT 134.790 264.140 135.410 264.325 ;
        RECT 103.190 263.910 135.410 264.140 ;
        RECT 103.190 263.725 103.810 263.910 ;
        RECT 134.790 263.725 135.410 263.910 ;
        RECT 14.240 263.645 15.860 263.655 ;
        RECT 46.690 263.645 48.310 263.655 ;
        RECT 79.140 263.645 80.760 263.655 ;
        RECT 111.590 263.645 113.210 263.655 ;
        RECT 6.690 263.275 37.210 263.645 ;
        RECT 39.140 263.275 69.660 263.645 ;
        RECT 71.590 263.275 102.110 263.645 ;
        RECT 104.040 263.275 134.560 263.645 ;
        RECT 0.130 262.890 2.420 263.230 ;
        RECT 3.165 262.890 4.650 263.230 ;
        RECT 0.130 262.255 0.730 262.890 ;
        RECT 0.130 262.025 1.860 262.255 ;
        RECT 2.160 262.025 3.820 262.255 ;
        RECT 0.130 260.015 0.730 262.025 ;
        RECT 2.160 260.990 2.390 262.025 ;
        RECT 2.795 260.735 3.025 261.780 ;
        RECT 4.050 260.735 4.650 262.890 ;
        RECT 6.690 262.555 37.210 262.935 ;
        RECT 39.140 262.555 69.660 262.935 ;
        RECT 71.590 262.555 102.110 262.935 ;
        RECT 104.040 262.555 134.560 262.935 ;
        RECT 5.840 262.300 6.460 262.485 ;
        RECT 37.440 262.300 38.060 262.485 ;
        RECT 5.840 262.070 38.060 262.300 ;
        RECT 5.840 261.885 6.460 262.070 ;
        RECT 37.440 261.885 38.060 262.070 ;
        RECT 38.290 262.300 38.910 262.485 ;
        RECT 69.890 262.300 70.510 262.485 ;
        RECT 38.290 262.070 70.510 262.300 ;
        RECT 38.290 261.885 38.910 262.070 ;
        RECT 69.890 261.885 70.510 262.070 ;
        RECT 70.740 262.300 71.360 262.485 ;
        RECT 102.340 262.300 102.960 262.485 ;
        RECT 70.740 262.070 102.960 262.300 ;
        RECT 70.740 261.885 71.360 262.070 ;
        RECT 102.340 261.885 102.960 262.070 ;
        RECT 103.190 262.300 103.810 262.485 ;
        RECT 134.790 262.300 135.410 262.485 ;
        RECT 103.190 262.070 135.410 262.300 ;
        RECT 103.190 261.885 103.810 262.070 ;
        RECT 134.790 261.885 135.410 262.070 ;
        RECT 10.400 261.805 12.020 261.815 ;
        RECT 42.850 261.805 44.470 261.815 ;
        RECT 75.300 261.805 76.920 261.815 ;
        RECT 107.750 261.805 109.370 261.815 ;
        RECT 6.690 261.435 37.210 261.805 ;
        RECT 39.140 261.435 69.660 261.805 ;
        RECT 71.590 261.435 102.110 261.805 ;
        RECT 104.040 261.435 134.560 261.805 ;
        RECT 0.960 260.505 3.025 260.735 ;
        RECT 3.255 260.505 4.650 260.735 ;
        RECT 6.690 260.715 37.210 261.095 ;
        RECT 39.140 260.715 69.660 261.095 ;
        RECT 71.590 260.715 102.110 261.095 ;
        RECT 104.040 260.715 134.560 261.095 ;
        RECT 0.130 259.785 1.860 260.015 ;
        RECT 2.160 259.785 3.820 260.015 ;
        RECT 0.130 257.630 0.730 259.785 ;
        RECT 2.160 258.750 2.390 259.785 ;
        RECT 2.795 258.495 3.025 259.540 ;
        RECT 4.050 258.495 4.650 260.505 ;
        RECT 5.840 260.460 6.460 260.645 ;
        RECT 37.440 260.460 38.060 260.645 ;
        RECT 5.840 260.230 38.060 260.460 ;
        RECT 5.840 260.045 6.460 260.230 ;
        RECT 37.440 260.045 38.060 260.230 ;
        RECT 38.290 260.460 38.910 260.645 ;
        RECT 69.890 260.460 70.510 260.645 ;
        RECT 38.290 260.230 70.510 260.460 ;
        RECT 38.290 260.045 38.910 260.230 ;
        RECT 69.890 260.045 70.510 260.230 ;
        RECT 70.740 260.460 71.360 260.645 ;
        RECT 102.340 260.460 102.960 260.645 ;
        RECT 70.740 260.230 102.960 260.460 ;
        RECT 70.740 260.045 71.360 260.230 ;
        RECT 102.340 260.045 102.960 260.230 ;
        RECT 103.190 260.460 103.810 260.645 ;
        RECT 134.790 260.460 135.410 260.645 ;
        RECT 103.190 260.230 135.410 260.460 ;
        RECT 103.190 260.045 103.810 260.230 ;
        RECT 134.790 260.045 135.410 260.230 ;
        RECT 6.690 259.595 37.210 259.965 ;
        RECT 39.140 259.595 69.660 259.965 ;
        RECT 71.590 259.595 102.110 259.965 ;
        RECT 104.040 259.595 134.560 259.965 ;
        RECT 0.960 258.265 3.025 258.495 ;
        RECT 3.255 258.265 4.650 258.495 ;
        RECT 4.050 257.630 4.650 258.265 ;
        RECT 0.130 257.290 2.420 257.630 ;
        RECT 3.165 257.290 4.650 257.630 ;
        RECT 0.130 256.655 0.730 257.290 ;
        RECT 0.130 256.425 1.710 256.655 ;
        RECT 0.130 254.385 0.730 256.425 ;
        RECT 2.140 256.195 2.500 256.280 ;
        RECT 1.010 255.965 2.500 256.195 ;
        RECT 1.010 255.815 1.370 255.965 ;
        RECT 0.960 255.180 1.910 255.585 ;
        RECT 0.130 254.155 1.420 254.385 ;
        RECT 0.130 253.195 0.730 254.155 ;
        RECT 1.650 253.835 1.910 255.180 ;
        RECT 2.140 254.530 2.500 255.965 ;
        RECT 2.730 254.630 3.080 255.830 ;
        RECT 3.440 255.220 3.820 256.865 ;
        RECT 2.520 253.835 2.870 253.895 ;
        RECT 3.440 253.835 3.780 254.440 ;
        RECT 1.650 253.575 3.780 253.835 ;
        RECT 2.520 253.515 2.870 253.575 ;
        RECT 4.050 253.295 4.650 257.290 ;
        RECT 6.495 256.810 8.245 259.595 ;
        RECT 8.885 256.810 9.695 257.810 ;
        RECT 10.335 256.810 12.085 259.105 ;
        RECT 12.725 256.810 13.535 257.810 ;
        RECT 14.175 256.810 15.925 259.105 ;
        RECT 16.565 256.810 17.375 257.810 ;
        RECT 18.015 256.810 19.765 259.105 ;
        RECT 20.405 256.810 21.215 257.810 ;
        RECT 21.855 256.810 23.605 259.105 ;
        RECT 24.245 256.810 25.055 257.810 ;
        RECT 25.695 256.810 27.445 259.105 ;
        RECT 28.085 256.810 28.895 257.810 ;
        RECT 29.535 256.810 31.285 259.105 ;
        RECT 31.925 256.810 32.735 257.810 ;
        RECT 33.375 256.810 35.125 259.105 ;
        RECT 35.765 256.810 36.575 257.810 ;
        RECT 38.945 256.810 40.695 259.595 ;
        RECT 41.335 256.810 42.145 257.810 ;
        RECT 42.785 256.810 44.535 259.105 ;
        RECT 45.175 256.810 45.985 257.810 ;
        RECT 46.625 256.810 48.375 259.105 ;
        RECT 49.015 256.810 49.825 257.810 ;
        RECT 50.465 256.810 52.215 259.105 ;
        RECT 52.855 256.810 53.665 257.810 ;
        RECT 54.305 256.810 56.055 259.105 ;
        RECT 56.695 256.810 57.505 257.810 ;
        RECT 58.145 256.810 59.895 259.105 ;
        RECT 60.535 256.810 61.345 257.810 ;
        RECT 61.985 256.810 63.735 259.105 ;
        RECT 64.375 256.810 65.185 257.810 ;
        RECT 65.825 256.810 67.575 259.105 ;
        RECT 68.215 256.810 69.025 257.810 ;
        RECT 71.395 256.810 73.145 259.595 ;
        RECT 73.785 256.810 74.595 257.810 ;
        RECT 75.235 256.810 76.985 259.105 ;
        RECT 77.625 256.810 78.435 257.810 ;
        RECT 79.075 256.810 80.825 259.105 ;
        RECT 81.465 256.810 82.275 257.810 ;
        RECT 82.915 256.810 84.665 259.105 ;
        RECT 85.305 256.810 86.115 257.810 ;
        RECT 86.755 256.810 88.505 259.105 ;
        RECT 89.145 256.810 89.955 257.810 ;
        RECT 90.595 256.810 92.345 259.105 ;
        RECT 92.985 256.810 93.795 257.810 ;
        RECT 94.435 256.810 96.185 259.105 ;
        RECT 96.825 256.810 97.635 257.810 ;
        RECT 98.275 256.810 100.025 259.105 ;
        RECT 100.665 256.810 101.475 257.810 ;
        RECT 103.845 256.810 105.595 259.595 ;
        RECT 106.235 256.810 107.045 257.810 ;
        RECT 107.685 256.810 109.435 259.105 ;
        RECT 110.075 256.810 110.885 257.810 ;
        RECT 111.525 256.810 113.275 259.105 ;
        RECT 113.915 256.810 114.725 257.810 ;
        RECT 115.365 256.810 117.115 259.105 ;
        RECT 117.755 256.810 118.565 257.810 ;
        RECT 119.205 256.810 120.955 259.105 ;
        RECT 121.595 256.810 122.405 257.810 ;
        RECT 123.045 256.810 124.795 259.105 ;
        RECT 125.435 256.810 126.245 257.810 ;
        RECT 126.885 256.810 128.635 259.105 ;
        RECT 129.275 256.810 130.085 257.810 ;
        RECT 130.725 256.810 132.475 259.105 ;
        RECT 133.115 256.810 133.925 257.810 ;
        RECT 136.340 257.000 136.710 275.510 ;
        RECT 137.360 271.875 137.730 275.510 ;
        RECT 137.355 271.495 137.735 271.875 ;
        RECT 137.360 268.875 137.730 271.495 ;
        RECT 137.355 268.495 137.735 268.875 ;
        RECT 137.360 265.875 137.730 268.495 ;
        RECT 137.355 265.495 137.735 265.875 ;
        RECT 137.360 262.875 137.730 265.495 ;
        RECT 137.355 262.495 137.735 262.875 ;
        RECT 137.360 259.875 137.730 262.495 ;
        RECT 137.355 259.495 137.735 259.875 ;
        RECT 136.340 256.620 136.720 257.000 ;
        RECT 136.340 255.550 136.710 256.620 ;
        RECT 6.965 254.360 7.775 255.360 ;
        RECT 0.130 252.965 1.820 253.195 ;
        RECT 3.190 253.065 4.650 253.295 ;
        RECT 0.130 250.955 0.730 252.965 ;
        RECT 2.150 252.505 3.150 252.830 ;
        RECT 0.960 251.945 3.820 252.275 ;
        RECT 0.130 250.725 1.820 250.955 ;
        RECT 0.130 248.715 0.730 250.725 ;
        RECT 2.535 250.590 2.800 251.945 ;
        RECT 4.050 251.055 4.650 253.065 ;
        RECT 8.415 252.530 10.165 255.360 ;
        RECT 10.805 254.360 11.615 255.360 ;
        RECT 12.255 253.065 14.005 255.360 ;
        RECT 14.645 254.360 15.455 255.360 ;
        RECT 16.095 253.065 17.845 255.360 ;
        RECT 18.485 254.360 19.295 255.360 ;
        RECT 19.935 253.065 21.685 255.360 ;
        RECT 22.325 254.360 23.135 255.360 ;
        RECT 23.775 253.065 25.525 255.360 ;
        RECT 26.165 254.360 26.975 255.360 ;
        RECT 27.615 253.065 29.365 255.360 ;
        RECT 30.005 254.360 30.815 255.360 ;
        RECT 31.455 253.065 33.205 255.360 ;
        RECT 33.845 254.360 34.655 255.360 ;
        RECT 35.295 253.065 37.045 255.360 ;
        RECT 39.415 254.360 40.225 255.360 ;
        RECT 40.865 252.530 42.615 255.360 ;
        RECT 43.255 254.360 44.065 255.360 ;
        RECT 44.705 253.065 46.455 255.360 ;
        RECT 47.095 254.360 47.905 255.360 ;
        RECT 48.545 253.065 50.295 255.360 ;
        RECT 50.935 254.360 51.745 255.360 ;
        RECT 52.385 253.065 54.135 255.360 ;
        RECT 54.775 254.360 55.585 255.360 ;
        RECT 56.225 253.065 57.975 255.360 ;
        RECT 58.615 254.360 59.425 255.360 ;
        RECT 60.065 253.065 61.815 255.360 ;
        RECT 62.455 254.360 63.265 255.360 ;
        RECT 63.905 253.065 65.655 255.360 ;
        RECT 66.295 254.360 67.105 255.360 ;
        RECT 67.745 253.065 69.495 255.360 ;
        RECT 71.865 254.360 72.675 255.360 ;
        RECT 73.315 252.530 75.065 255.360 ;
        RECT 75.705 254.360 76.515 255.360 ;
        RECT 77.155 253.065 78.905 255.360 ;
        RECT 79.545 254.360 80.355 255.360 ;
        RECT 80.995 253.065 82.745 255.360 ;
        RECT 83.385 254.360 84.195 255.360 ;
        RECT 84.835 253.065 86.585 255.360 ;
        RECT 87.225 254.360 88.035 255.360 ;
        RECT 88.675 253.065 90.425 255.360 ;
        RECT 91.065 254.360 91.875 255.360 ;
        RECT 92.515 253.065 94.265 255.360 ;
        RECT 94.905 254.360 95.715 255.360 ;
        RECT 96.355 253.065 98.105 255.360 ;
        RECT 98.745 254.360 99.555 255.360 ;
        RECT 100.195 253.065 101.945 255.360 ;
        RECT 104.315 254.360 105.125 255.360 ;
        RECT 105.765 252.530 107.515 255.360 ;
        RECT 108.155 254.360 108.965 255.360 ;
        RECT 109.605 253.065 111.355 255.360 ;
        RECT 111.995 254.360 112.805 255.360 ;
        RECT 113.445 253.065 115.195 255.360 ;
        RECT 115.835 254.360 116.645 255.360 ;
        RECT 117.285 253.065 119.035 255.360 ;
        RECT 119.675 254.360 120.485 255.360 ;
        RECT 121.125 253.065 122.875 255.360 ;
        RECT 123.515 254.360 124.325 255.360 ;
        RECT 124.965 253.065 126.715 255.360 ;
        RECT 127.355 254.360 128.165 255.360 ;
        RECT 128.805 253.065 130.555 255.360 ;
        RECT 131.195 254.360 132.005 255.360 ;
        RECT 132.645 253.065 134.395 255.360 ;
        RECT 136.340 255.170 136.720 255.550 ;
        RECT 6.690 252.160 37.210 252.530 ;
        RECT 39.140 252.160 69.660 252.530 ;
        RECT 71.590 252.160 102.110 252.530 ;
        RECT 104.040 252.160 134.560 252.530 ;
        RECT 5.840 251.895 6.460 252.080 ;
        RECT 37.440 251.895 38.060 252.080 ;
        RECT 5.840 251.665 38.060 251.895 ;
        RECT 5.840 251.480 6.460 251.665 ;
        RECT 37.440 251.480 38.060 251.665 ;
        RECT 38.290 251.895 38.910 252.080 ;
        RECT 69.890 251.895 70.510 252.080 ;
        RECT 38.290 251.665 70.510 251.895 ;
        RECT 38.290 251.480 38.910 251.665 ;
        RECT 69.890 251.480 70.510 251.665 ;
        RECT 70.740 251.895 71.360 252.080 ;
        RECT 102.340 251.895 102.960 252.080 ;
        RECT 70.740 251.665 102.960 251.895 ;
        RECT 70.740 251.480 71.360 251.665 ;
        RECT 102.340 251.480 102.960 251.665 ;
        RECT 103.190 251.895 103.810 252.080 ;
        RECT 134.790 251.895 135.410 252.080 ;
        RECT 103.190 251.665 135.410 251.895 ;
        RECT 103.190 251.480 103.810 251.665 ;
        RECT 134.790 251.480 135.410 251.665 ;
        RECT 3.190 250.825 4.650 251.055 ;
        RECT 6.690 251.030 37.210 251.410 ;
        RECT 39.140 251.030 69.660 251.410 ;
        RECT 71.590 251.030 102.110 251.410 ;
        RECT 104.040 251.030 134.560 251.410 ;
        RECT 2.150 250.265 3.150 250.590 ;
        RECT 0.960 249.705 3.820 250.035 ;
        RECT 4.050 248.815 4.650 250.825 ;
        RECT 6.690 250.320 37.210 250.690 ;
        RECT 39.140 250.320 69.660 250.690 ;
        RECT 71.590 250.320 102.110 250.690 ;
        RECT 104.040 250.320 134.560 250.690 ;
        RECT 12.320 250.310 13.940 250.320 ;
        RECT 44.770 250.310 46.390 250.320 ;
        RECT 77.220 250.310 78.840 250.320 ;
        RECT 109.670 250.310 111.290 250.320 ;
        RECT 5.840 250.055 6.460 250.240 ;
        RECT 37.440 250.055 38.060 250.240 ;
        RECT 5.840 249.825 38.060 250.055 ;
        RECT 5.840 249.640 6.460 249.825 ;
        RECT 37.440 249.640 38.060 249.825 ;
        RECT 38.290 250.055 38.910 250.240 ;
        RECT 69.890 250.055 70.510 250.240 ;
        RECT 38.290 249.825 70.510 250.055 ;
        RECT 38.290 249.640 38.910 249.825 ;
        RECT 69.890 249.640 70.510 249.825 ;
        RECT 70.740 250.055 71.360 250.240 ;
        RECT 102.340 250.055 102.960 250.240 ;
        RECT 70.740 249.825 102.960 250.055 ;
        RECT 70.740 249.640 71.360 249.825 ;
        RECT 102.340 249.640 102.960 249.825 ;
        RECT 103.190 250.055 103.810 250.240 ;
        RECT 134.790 250.055 135.410 250.240 ;
        RECT 103.190 249.825 135.410 250.055 ;
        RECT 103.190 249.640 103.810 249.825 ;
        RECT 134.790 249.640 135.410 249.825 ;
        RECT 6.690 249.190 37.210 249.570 ;
        RECT 39.140 249.190 69.660 249.570 ;
        RECT 71.590 249.190 102.110 249.570 ;
        RECT 104.040 249.190 134.560 249.570 ;
        RECT 0.130 248.485 1.820 248.715 ;
        RECT 3.190 248.585 4.650 248.815 ;
        RECT 0.130 246.430 0.730 248.485 ;
        RECT 2.150 248.025 3.150 248.350 ;
        RECT 0.960 247.465 3.820 247.795 ;
        RECT 2.300 247.340 2.680 247.465 ;
        RECT 4.050 246.430 4.650 248.585 ;
        RECT 6.690 248.475 37.210 248.845 ;
        RECT 39.140 248.475 69.660 248.845 ;
        RECT 71.590 248.475 102.110 248.845 ;
        RECT 104.040 248.475 134.560 248.845 ;
        RECT 16.160 248.465 17.780 248.475 ;
        RECT 48.610 248.465 50.230 248.475 ;
        RECT 81.060 248.465 82.680 248.475 ;
        RECT 113.510 248.465 115.130 248.475 ;
        RECT 5.840 248.210 6.460 248.395 ;
        RECT 37.440 248.210 38.060 248.395 ;
        RECT 5.840 247.980 38.060 248.210 ;
        RECT 5.840 247.795 6.460 247.980 ;
        RECT 37.440 247.795 38.060 247.980 ;
        RECT 38.290 248.210 38.910 248.395 ;
        RECT 69.890 248.210 70.510 248.395 ;
        RECT 38.290 247.980 70.510 248.210 ;
        RECT 38.290 247.795 38.910 247.980 ;
        RECT 69.890 247.795 70.510 247.980 ;
        RECT 70.740 248.210 71.360 248.395 ;
        RECT 102.340 248.210 102.960 248.395 ;
        RECT 70.740 247.980 102.960 248.210 ;
        RECT 70.740 247.795 71.360 247.980 ;
        RECT 102.340 247.795 102.960 247.980 ;
        RECT 103.190 248.210 103.810 248.395 ;
        RECT 134.790 248.210 135.410 248.395 ;
        RECT 103.190 247.980 135.410 248.210 ;
        RECT 103.190 247.795 103.810 247.980 ;
        RECT 134.790 247.795 135.410 247.980 ;
        RECT 6.690 247.345 37.210 247.725 ;
        RECT 39.140 247.345 69.660 247.725 ;
        RECT 71.590 247.345 102.110 247.725 ;
        RECT 104.040 247.345 134.560 247.725 ;
        RECT 6.700 246.555 37.200 246.995 ;
        RECT 39.150 246.555 69.650 246.995 ;
        RECT 71.600 246.555 102.100 246.995 ;
        RECT 104.050 246.555 134.550 246.995 ;
        RECT 0.130 246.090 2.420 246.430 ;
        RECT 3.165 246.090 4.650 246.430 ;
        RECT 0.130 245.310 0.730 246.090 ;
        RECT 4.050 245.310 4.650 246.090 ;
        RECT 6.690 245.835 37.210 246.205 ;
        RECT 39.140 245.835 69.660 246.205 ;
        RECT 71.590 245.835 102.110 246.205 ;
        RECT 104.040 245.835 134.560 246.205 ;
        RECT 20.000 245.825 21.620 245.835 ;
        RECT 52.450 245.825 54.070 245.835 ;
        RECT 84.900 245.825 86.520 245.835 ;
        RECT 117.350 245.825 118.970 245.835 ;
        RECT 0.130 244.970 2.420 245.310 ;
        RECT 3.165 244.970 4.650 245.310 ;
        RECT 5.840 245.570 6.460 245.755 ;
        RECT 37.440 245.570 38.060 245.755 ;
        RECT 5.840 245.340 38.060 245.570 ;
        RECT 5.840 245.155 6.460 245.340 ;
        RECT 37.440 245.155 38.060 245.340 ;
        RECT 38.290 245.570 38.910 245.755 ;
        RECT 69.890 245.570 70.510 245.755 ;
        RECT 38.290 245.340 70.510 245.570 ;
        RECT 38.290 245.155 38.910 245.340 ;
        RECT 69.890 245.155 70.510 245.340 ;
        RECT 70.740 245.570 71.360 245.755 ;
        RECT 102.340 245.570 102.960 245.755 ;
        RECT 70.740 245.340 102.960 245.570 ;
        RECT 70.740 245.155 71.360 245.340 ;
        RECT 102.340 245.155 102.960 245.340 ;
        RECT 103.190 245.570 103.810 245.755 ;
        RECT 134.790 245.570 135.410 245.755 ;
        RECT 103.190 245.340 135.410 245.570 ;
        RECT 103.190 245.155 103.810 245.340 ;
        RECT 134.790 245.155 135.410 245.340 ;
        RECT 0.130 244.335 0.730 244.970 ;
        RECT 0.130 244.105 1.860 244.335 ;
        RECT 2.160 244.105 3.820 244.335 ;
        RECT 0.130 242.095 0.730 244.105 ;
        RECT 2.160 243.070 2.390 244.105 ;
        RECT 2.795 242.815 3.025 243.860 ;
        RECT 4.050 242.815 4.650 244.970 ;
        RECT 6.690 244.705 37.210 245.085 ;
        RECT 39.140 244.705 69.660 245.085 ;
        RECT 71.590 244.705 102.110 245.085 ;
        RECT 104.040 244.705 134.560 245.085 ;
        RECT 6.690 243.995 37.210 244.365 ;
        RECT 39.140 243.995 69.660 244.365 ;
        RECT 71.590 243.995 102.110 244.365 ;
        RECT 104.040 243.995 134.560 244.365 ;
        RECT 23.840 243.985 25.460 243.995 ;
        RECT 56.290 243.985 57.910 243.995 ;
        RECT 88.740 243.985 90.360 243.995 ;
        RECT 121.190 243.985 122.810 243.995 ;
        RECT 5.840 243.730 6.460 243.915 ;
        RECT 37.440 243.730 38.060 243.915 ;
        RECT 5.840 243.500 38.060 243.730 ;
        RECT 5.840 243.315 6.460 243.500 ;
        RECT 37.440 243.315 38.060 243.500 ;
        RECT 38.290 243.730 38.910 243.915 ;
        RECT 69.890 243.730 70.510 243.915 ;
        RECT 38.290 243.500 70.510 243.730 ;
        RECT 38.290 243.315 38.910 243.500 ;
        RECT 69.890 243.315 70.510 243.500 ;
        RECT 70.740 243.730 71.360 243.915 ;
        RECT 102.340 243.730 102.960 243.915 ;
        RECT 70.740 243.500 102.960 243.730 ;
        RECT 70.740 243.315 71.360 243.500 ;
        RECT 102.340 243.315 102.960 243.500 ;
        RECT 103.190 243.730 103.810 243.915 ;
        RECT 134.790 243.730 135.410 243.915 ;
        RECT 103.190 243.500 135.410 243.730 ;
        RECT 103.190 243.315 103.810 243.500 ;
        RECT 134.790 243.315 135.410 243.500 ;
        RECT 6.690 242.865 37.210 243.245 ;
        RECT 39.140 242.865 69.660 243.245 ;
        RECT 71.590 242.865 102.110 243.245 ;
        RECT 104.040 242.865 134.560 243.245 ;
        RECT 0.960 242.585 3.025 242.815 ;
        RECT 3.255 242.585 4.650 242.815 ;
        RECT 0.130 241.865 1.860 242.095 ;
        RECT 2.160 241.865 3.820 242.095 ;
        RECT 0.130 239.855 0.730 241.865 ;
        RECT 2.160 240.830 2.390 241.865 ;
        RECT 2.795 240.575 3.025 241.620 ;
        RECT 4.050 240.575 4.650 242.585 ;
        RECT 6.690 242.150 37.210 242.520 ;
        RECT 39.140 242.150 69.660 242.520 ;
        RECT 71.590 242.150 102.110 242.520 ;
        RECT 104.040 242.150 134.560 242.520 ;
        RECT 27.680 242.140 29.300 242.150 ;
        RECT 60.130 242.140 61.750 242.150 ;
        RECT 92.580 242.140 94.200 242.150 ;
        RECT 125.030 242.140 126.650 242.150 ;
        RECT 5.840 241.885 6.460 242.070 ;
        RECT 37.440 241.885 38.060 242.070 ;
        RECT 5.840 241.655 38.060 241.885 ;
        RECT 5.840 241.470 6.460 241.655 ;
        RECT 37.440 241.470 38.060 241.655 ;
        RECT 38.290 241.885 38.910 242.070 ;
        RECT 69.890 241.885 70.510 242.070 ;
        RECT 38.290 241.655 70.510 241.885 ;
        RECT 38.290 241.470 38.910 241.655 ;
        RECT 69.890 241.470 70.510 241.655 ;
        RECT 70.740 241.885 71.360 242.070 ;
        RECT 102.340 241.885 102.960 242.070 ;
        RECT 70.740 241.655 102.960 241.885 ;
        RECT 70.740 241.470 71.360 241.655 ;
        RECT 102.340 241.470 102.960 241.655 ;
        RECT 103.190 241.885 103.810 242.070 ;
        RECT 134.790 241.885 135.410 242.070 ;
        RECT 103.190 241.655 135.410 241.885 ;
        RECT 103.190 241.470 103.810 241.655 ;
        RECT 134.790 241.470 135.410 241.655 ;
        RECT 6.690 241.020 37.210 241.400 ;
        RECT 39.140 241.020 69.660 241.400 ;
        RECT 71.590 241.020 102.110 241.400 ;
        RECT 104.040 241.020 134.560 241.400 ;
        RECT 0.960 240.345 3.025 240.575 ;
        RECT 3.255 240.345 4.650 240.575 ;
        RECT 0.130 239.625 1.860 239.855 ;
        RECT 2.160 239.625 3.820 239.855 ;
        RECT 0.130 237.450 0.730 239.625 ;
        RECT 2.160 238.590 2.390 239.625 ;
        RECT 2.795 238.335 3.025 239.380 ;
        RECT 4.050 238.335 4.650 240.345 ;
        RECT 6.700 240.230 37.200 240.670 ;
        RECT 39.150 240.230 69.650 240.670 ;
        RECT 71.600 240.230 102.100 240.670 ;
        RECT 104.050 240.230 134.550 240.670 ;
        RECT 6.690 239.510 37.210 239.880 ;
        RECT 39.140 239.510 69.660 239.880 ;
        RECT 71.590 239.510 102.110 239.880 ;
        RECT 104.040 239.510 134.560 239.880 ;
        RECT 31.520 239.500 33.140 239.510 ;
        RECT 63.970 239.500 65.590 239.510 ;
        RECT 96.420 239.500 98.040 239.510 ;
        RECT 128.870 239.500 130.490 239.510 ;
        RECT 5.840 239.245 6.460 239.430 ;
        RECT 37.440 239.245 38.060 239.430 ;
        RECT 5.840 239.015 38.060 239.245 ;
        RECT 5.840 238.830 6.460 239.015 ;
        RECT 37.440 238.830 38.060 239.015 ;
        RECT 38.290 239.245 38.910 239.430 ;
        RECT 69.890 239.245 70.510 239.430 ;
        RECT 38.290 239.015 70.510 239.245 ;
        RECT 38.290 238.830 38.910 239.015 ;
        RECT 69.890 238.830 70.510 239.015 ;
        RECT 70.740 239.245 71.360 239.430 ;
        RECT 102.340 239.245 102.960 239.430 ;
        RECT 70.740 239.015 102.960 239.245 ;
        RECT 70.740 238.830 71.360 239.015 ;
        RECT 102.340 238.830 102.960 239.015 ;
        RECT 103.190 239.245 103.810 239.430 ;
        RECT 134.790 239.245 135.410 239.430 ;
        RECT 103.190 239.015 135.410 239.245 ;
        RECT 103.190 238.830 103.810 239.015 ;
        RECT 134.790 238.830 135.410 239.015 ;
        RECT 6.690 238.380 37.210 238.760 ;
        RECT 39.140 238.380 69.660 238.760 ;
        RECT 71.590 238.380 102.110 238.760 ;
        RECT 104.040 238.380 134.560 238.760 ;
        RECT 0.960 238.105 3.025 238.335 ;
        RECT 3.255 238.105 4.650 238.335 ;
        RECT 4.050 237.450 4.650 238.105 ;
        RECT 6.690 237.670 37.210 238.040 ;
        RECT 39.140 237.670 69.660 238.040 ;
        RECT 71.590 237.670 102.110 238.040 ;
        RECT 104.040 237.670 134.560 238.040 ;
        RECT 35.360 237.660 36.980 237.670 ;
        RECT 67.810 237.660 69.430 237.670 ;
        RECT 100.260 237.660 101.880 237.670 ;
        RECT 132.710 237.660 134.330 237.670 ;
        RECT 0.130 237.110 2.430 237.450 ;
        RECT 3.160 237.110 4.650 237.450 ;
        RECT 0.130 236.145 0.730 237.110 ;
        RECT 4.050 236.145 4.650 237.110 ;
        RECT 5.840 237.405 6.460 237.590 ;
        RECT 37.440 237.405 38.060 237.590 ;
        RECT 5.840 237.175 38.060 237.405 ;
        RECT 5.840 236.990 6.460 237.175 ;
        RECT 37.440 236.990 38.060 237.175 ;
        RECT 38.290 237.405 38.910 237.590 ;
        RECT 69.890 237.405 70.510 237.590 ;
        RECT 38.290 237.175 70.510 237.405 ;
        RECT 38.290 236.990 38.910 237.175 ;
        RECT 69.890 236.990 70.510 237.175 ;
        RECT 70.740 237.405 71.360 237.590 ;
        RECT 102.340 237.405 102.960 237.590 ;
        RECT 70.740 237.175 102.960 237.405 ;
        RECT 70.740 236.990 71.360 237.175 ;
        RECT 102.340 236.990 102.960 237.175 ;
        RECT 103.190 237.405 103.810 237.590 ;
        RECT 134.790 237.405 135.410 237.590 ;
        RECT 103.190 237.175 135.410 237.405 ;
        RECT 136.340 237.240 136.710 255.170 ;
        RECT 137.360 253.875 137.730 259.495 ;
        RECT 138.380 257.000 138.750 275.510 ;
        RECT 139.400 271.875 139.770 275.510 ;
        RECT 139.395 271.495 139.775 271.875 ;
        RECT 139.400 268.875 139.770 271.495 ;
        RECT 139.395 268.495 139.775 268.875 ;
        RECT 139.400 265.875 139.770 268.495 ;
        RECT 139.395 265.495 139.775 265.875 ;
        RECT 139.400 262.875 139.770 265.495 ;
        RECT 139.395 262.495 139.775 262.875 ;
        RECT 139.400 259.875 139.770 262.495 ;
        RECT 139.395 259.495 139.775 259.875 ;
        RECT 138.380 256.620 138.760 257.000 ;
        RECT 138.380 255.550 138.750 256.620 ;
        RECT 138.380 255.170 138.760 255.550 ;
        RECT 137.355 253.495 137.735 253.875 ;
        RECT 137.360 250.875 137.730 253.495 ;
        RECT 137.355 250.495 137.735 250.875 ;
        RECT 137.360 247.875 137.730 250.495 ;
        RECT 137.355 247.495 137.735 247.875 ;
        RECT 137.360 244.875 137.730 247.495 ;
        RECT 137.355 244.495 137.735 244.875 ;
        RECT 137.360 241.875 137.730 244.495 ;
        RECT 137.355 241.495 137.735 241.875 ;
        RECT 137.360 238.875 137.730 241.495 ;
        RECT 137.355 238.495 137.735 238.875 ;
        RECT 137.360 237.240 137.730 238.495 ;
        RECT 138.380 237.240 138.750 255.170 ;
        RECT 139.400 253.875 139.770 259.495 ;
        RECT 139.395 253.495 139.775 253.875 ;
        RECT 139.400 250.875 139.770 253.495 ;
        RECT 139.395 250.495 139.775 250.875 ;
        RECT 139.400 247.875 139.770 250.495 ;
        RECT 139.395 247.495 139.775 247.875 ;
        RECT 139.400 244.875 139.770 247.495 ;
        RECT 139.395 244.495 139.775 244.875 ;
        RECT 139.400 241.875 139.770 244.495 ;
        RECT 139.395 241.495 139.775 241.875 ;
        RECT 139.400 238.875 139.770 241.495 ;
        RECT 139.395 238.495 139.775 238.875 ;
        RECT 139.400 237.240 139.770 238.495 ;
        RECT 140.420 237.240 140.800 275.510 ;
        RECT 141.150 237.250 141.590 275.500 ;
        RECT 103.190 236.990 103.810 237.175 ;
        RECT 134.790 236.990 135.410 237.175 ;
        RECT 6.690 236.540 37.210 236.920 ;
        RECT 39.140 236.540 69.660 236.920 ;
        RECT 71.590 236.540 102.110 236.920 ;
        RECT 104.040 236.540 134.560 236.920 ;
        RECT 0.130 235.805 2.430 236.145 ;
        RECT 3.160 235.805 4.650 236.145 ;
        RECT 6.690 235.820 37.210 236.200 ;
        RECT 39.140 235.820 69.660 236.200 ;
        RECT 71.590 235.820 102.110 236.200 ;
        RECT 104.040 235.820 134.560 236.200 ;
        RECT 0.130 235.190 0.730 235.805 ;
        RECT 0.130 234.960 1.860 235.190 ;
        RECT 2.160 234.960 3.820 235.190 ;
        RECT 0.130 232.950 0.730 234.960 ;
        RECT 2.160 233.925 2.390 234.960 ;
        RECT 2.795 233.670 3.025 234.715 ;
        RECT 4.050 233.670 4.650 235.805 ;
        RECT 5.840 235.565 6.460 235.750 ;
        RECT 37.440 235.565 38.060 235.750 ;
        RECT 5.840 235.335 38.060 235.565 ;
        RECT 5.840 235.150 6.460 235.335 ;
        RECT 37.440 235.150 38.060 235.335 ;
        RECT 38.290 235.565 38.910 235.750 ;
        RECT 69.890 235.565 70.510 235.750 ;
        RECT 38.290 235.335 70.510 235.565 ;
        RECT 38.290 235.150 38.910 235.335 ;
        RECT 69.890 235.150 70.510 235.335 ;
        RECT 70.740 235.565 71.360 235.750 ;
        RECT 102.340 235.565 102.960 235.750 ;
        RECT 70.740 235.335 102.960 235.565 ;
        RECT 70.740 235.150 71.360 235.335 ;
        RECT 102.340 235.150 102.960 235.335 ;
        RECT 103.190 235.565 103.810 235.750 ;
        RECT 134.790 235.565 135.410 235.750 ;
        RECT 103.190 235.335 135.410 235.565 ;
        RECT 103.190 235.150 103.810 235.335 ;
        RECT 134.790 235.150 135.410 235.335 ;
        RECT 33.440 235.070 35.060 235.080 ;
        RECT 65.890 235.070 67.510 235.080 ;
        RECT 98.340 235.070 99.960 235.080 ;
        RECT 130.790 235.070 132.410 235.080 ;
        RECT 6.690 234.700 37.210 235.070 ;
        RECT 39.140 234.700 69.660 235.070 ;
        RECT 71.590 234.700 102.110 235.070 ;
        RECT 104.040 234.700 134.560 235.070 ;
        RECT 6.690 233.980 37.210 234.360 ;
        RECT 39.140 233.980 69.660 234.360 ;
        RECT 71.590 233.980 102.110 234.360 ;
        RECT 104.040 233.980 134.560 234.360 ;
        RECT 0.960 233.440 3.025 233.670 ;
        RECT 3.255 233.440 4.650 233.670 ;
        RECT 0.130 232.720 1.860 232.950 ;
        RECT 2.160 232.720 3.820 232.950 ;
        RECT 0.130 230.710 0.730 232.720 ;
        RECT 2.160 231.685 2.390 232.720 ;
        RECT 2.795 231.430 3.025 232.475 ;
        RECT 4.050 231.430 4.650 233.440 ;
        RECT 5.840 233.725 6.460 233.910 ;
        RECT 37.440 233.725 38.060 233.910 ;
        RECT 5.840 233.495 38.060 233.725 ;
        RECT 5.840 233.310 6.460 233.495 ;
        RECT 37.440 233.310 38.060 233.495 ;
        RECT 38.290 233.725 38.910 233.910 ;
        RECT 69.890 233.725 70.510 233.910 ;
        RECT 38.290 233.495 70.510 233.725 ;
        RECT 38.290 233.310 38.910 233.495 ;
        RECT 69.890 233.310 70.510 233.495 ;
        RECT 70.740 233.725 71.360 233.910 ;
        RECT 102.340 233.725 102.960 233.910 ;
        RECT 70.740 233.495 102.960 233.725 ;
        RECT 70.740 233.310 71.360 233.495 ;
        RECT 102.340 233.310 102.960 233.495 ;
        RECT 103.190 233.725 103.810 233.910 ;
        RECT 134.790 233.725 135.410 233.910 ;
        RECT 103.190 233.495 135.410 233.725 ;
        RECT 103.190 233.310 103.810 233.495 ;
        RECT 134.790 233.310 135.410 233.495 ;
        RECT 29.600 233.230 31.220 233.240 ;
        RECT 62.050 233.230 63.670 233.240 ;
        RECT 94.500 233.230 96.120 233.240 ;
        RECT 126.950 233.230 128.570 233.240 ;
        RECT 6.690 232.860 37.210 233.230 ;
        RECT 39.140 232.860 69.660 233.230 ;
        RECT 71.590 232.860 102.110 233.230 ;
        RECT 104.040 232.860 134.560 233.230 ;
        RECT 6.700 232.065 37.200 232.505 ;
        RECT 39.150 232.065 69.650 232.505 ;
        RECT 71.600 232.065 102.100 232.505 ;
        RECT 104.050 232.065 134.550 232.505 ;
        RECT 0.960 231.200 3.025 231.430 ;
        RECT 3.255 231.200 4.650 231.430 ;
        RECT 6.690 231.335 37.210 231.715 ;
        RECT 39.140 231.335 69.660 231.715 ;
        RECT 71.590 231.335 102.110 231.715 ;
        RECT 104.040 231.335 134.560 231.715 ;
        RECT 0.130 230.480 1.860 230.710 ;
        RECT 2.160 230.480 3.820 230.710 ;
        RECT 0.130 228.470 0.730 230.480 ;
        RECT 2.160 229.445 2.390 230.480 ;
        RECT 2.795 229.190 3.025 230.235 ;
        RECT 4.050 229.190 4.650 231.200 ;
        RECT 5.840 231.080 6.460 231.265 ;
        RECT 37.440 231.080 38.060 231.265 ;
        RECT 5.840 230.850 38.060 231.080 ;
        RECT 5.840 230.665 6.460 230.850 ;
        RECT 37.440 230.665 38.060 230.850 ;
        RECT 38.290 231.080 38.910 231.265 ;
        RECT 69.890 231.080 70.510 231.265 ;
        RECT 38.290 230.850 70.510 231.080 ;
        RECT 38.290 230.665 38.910 230.850 ;
        RECT 69.890 230.665 70.510 230.850 ;
        RECT 70.740 231.080 71.360 231.265 ;
        RECT 102.340 231.080 102.960 231.265 ;
        RECT 70.740 230.850 102.960 231.080 ;
        RECT 70.740 230.665 71.360 230.850 ;
        RECT 102.340 230.665 102.960 230.850 ;
        RECT 103.190 231.080 103.810 231.265 ;
        RECT 134.790 231.080 135.410 231.265 ;
        RECT 103.190 230.850 135.410 231.080 ;
        RECT 103.190 230.665 103.810 230.850 ;
        RECT 134.790 230.665 135.410 230.850 ;
        RECT 25.760 230.585 27.380 230.595 ;
        RECT 58.210 230.585 59.830 230.595 ;
        RECT 90.660 230.585 92.280 230.595 ;
        RECT 123.110 230.585 124.730 230.595 ;
        RECT 6.690 230.215 37.210 230.585 ;
        RECT 39.140 230.215 69.660 230.585 ;
        RECT 71.590 230.215 102.110 230.585 ;
        RECT 104.040 230.215 134.560 230.585 ;
        RECT 6.690 229.495 37.210 229.875 ;
        RECT 39.140 229.495 69.660 229.875 ;
        RECT 71.590 229.495 102.110 229.875 ;
        RECT 104.040 229.495 134.560 229.875 ;
        RECT 0.960 228.960 3.025 229.190 ;
        RECT 3.255 228.960 4.650 229.190 ;
        RECT 0.130 228.240 1.860 228.470 ;
        RECT 2.160 228.240 3.820 228.470 ;
        RECT 0.130 226.230 0.730 228.240 ;
        RECT 2.160 227.205 2.390 228.240 ;
        RECT 2.795 226.950 3.025 227.995 ;
        RECT 4.050 226.950 4.650 228.960 ;
        RECT 5.840 229.240 6.460 229.425 ;
        RECT 37.440 229.240 38.060 229.425 ;
        RECT 5.840 229.010 38.060 229.240 ;
        RECT 5.840 228.825 6.460 229.010 ;
        RECT 37.440 228.825 38.060 229.010 ;
        RECT 38.290 229.240 38.910 229.425 ;
        RECT 69.890 229.240 70.510 229.425 ;
        RECT 38.290 229.010 70.510 229.240 ;
        RECT 38.290 228.825 38.910 229.010 ;
        RECT 69.890 228.825 70.510 229.010 ;
        RECT 70.740 229.240 71.360 229.425 ;
        RECT 102.340 229.240 102.960 229.425 ;
        RECT 70.740 229.010 102.960 229.240 ;
        RECT 70.740 228.825 71.360 229.010 ;
        RECT 102.340 228.825 102.960 229.010 ;
        RECT 103.190 229.240 103.810 229.425 ;
        RECT 134.790 229.240 135.410 229.425 ;
        RECT 103.190 229.010 135.410 229.240 ;
        RECT 103.190 228.825 103.810 229.010 ;
        RECT 134.790 228.825 135.410 229.010 ;
        RECT 21.920 228.745 23.540 228.755 ;
        RECT 54.370 228.745 55.990 228.755 ;
        RECT 86.820 228.745 88.440 228.755 ;
        RECT 119.270 228.745 120.890 228.755 ;
        RECT 6.690 228.375 37.210 228.745 ;
        RECT 39.140 228.375 69.660 228.745 ;
        RECT 71.590 228.375 102.110 228.745 ;
        RECT 104.040 228.375 134.560 228.745 ;
        RECT 6.690 227.655 37.210 228.035 ;
        RECT 39.140 227.655 69.660 228.035 ;
        RECT 71.590 227.655 102.110 228.035 ;
        RECT 104.040 227.655 134.560 228.035 ;
        RECT 5.840 227.400 6.460 227.585 ;
        RECT 37.440 227.400 38.060 227.585 ;
        RECT 5.840 227.170 38.060 227.400 ;
        RECT 5.840 226.985 6.460 227.170 ;
        RECT 37.440 226.985 38.060 227.170 ;
        RECT 38.290 227.400 38.910 227.585 ;
        RECT 69.890 227.400 70.510 227.585 ;
        RECT 38.290 227.170 70.510 227.400 ;
        RECT 38.290 226.985 38.910 227.170 ;
        RECT 69.890 226.985 70.510 227.170 ;
        RECT 70.740 227.400 71.360 227.585 ;
        RECT 102.340 227.400 102.960 227.585 ;
        RECT 70.740 227.170 102.960 227.400 ;
        RECT 70.740 226.985 71.360 227.170 ;
        RECT 102.340 226.985 102.960 227.170 ;
        RECT 103.190 227.400 103.810 227.585 ;
        RECT 134.790 227.400 135.410 227.585 ;
        RECT 103.190 227.170 135.410 227.400 ;
        RECT 103.190 226.985 103.810 227.170 ;
        RECT 134.790 226.985 135.410 227.170 ;
        RECT 0.960 226.720 3.025 226.950 ;
        RECT 3.255 226.720 4.650 226.950 ;
        RECT 18.080 226.905 19.700 226.915 ;
        RECT 50.530 226.905 52.150 226.915 ;
        RECT 82.980 226.905 84.600 226.915 ;
        RECT 115.430 226.905 117.050 226.915 ;
        RECT 0.130 226.000 1.860 226.230 ;
        RECT 2.160 226.000 3.820 226.230 ;
        RECT 0.130 223.845 0.730 226.000 ;
        RECT 2.160 224.965 2.390 226.000 ;
        RECT 2.795 224.710 3.025 225.755 ;
        RECT 4.050 224.710 4.650 226.720 ;
        RECT 6.690 226.535 37.210 226.905 ;
        RECT 39.140 226.535 69.660 226.905 ;
        RECT 71.590 226.535 102.110 226.905 ;
        RECT 104.040 226.535 134.560 226.905 ;
        RECT 6.700 225.740 37.200 226.180 ;
        RECT 39.150 225.740 69.650 226.180 ;
        RECT 71.600 225.740 102.100 226.180 ;
        RECT 104.050 225.740 134.550 226.180 ;
        RECT 6.690 225.010 37.210 225.390 ;
        RECT 39.140 225.010 69.660 225.390 ;
        RECT 71.590 225.010 102.110 225.390 ;
        RECT 104.040 225.010 134.560 225.390 ;
        RECT 0.960 224.480 3.025 224.710 ;
        RECT 3.255 224.480 4.650 224.710 ;
        RECT 4.050 223.845 4.650 224.480 ;
        RECT 5.840 224.755 6.460 224.940 ;
        RECT 37.440 224.755 38.060 224.940 ;
        RECT 5.840 224.525 38.060 224.755 ;
        RECT 5.840 224.340 6.460 224.525 ;
        RECT 37.440 224.340 38.060 224.525 ;
        RECT 38.290 224.755 38.910 224.940 ;
        RECT 69.890 224.755 70.510 224.940 ;
        RECT 38.290 224.525 70.510 224.755 ;
        RECT 38.290 224.340 38.910 224.525 ;
        RECT 69.890 224.340 70.510 224.525 ;
        RECT 70.740 224.755 71.360 224.940 ;
        RECT 102.340 224.755 102.960 224.940 ;
        RECT 70.740 224.525 102.960 224.755 ;
        RECT 70.740 224.340 71.360 224.525 ;
        RECT 102.340 224.340 102.960 224.525 ;
        RECT 103.190 224.755 103.810 224.940 ;
        RECT 134.790 224.755 135.410 224.940 ;
        RECT 103.190 224.525 135.410 224.755 ;
        RECT 103.190 224.340 103.810 224.525 ;
        RECT 134.790 224.340 135.410 224.525 ;
        RECT 14.240 224.260 15.860 224.270 ;
        RECT 46.690 224.260 48.310 224.270 ;
        RECT 79.140 224.260 80.760 224.270 ;
        RECT 111.590 224.260 113.210 224.270 ;
        RECT 6.690 223.890 37.210 224.260 ;
        RECT 39.140 223.890 69.660 224.260 ;
        RECT 71.590 223.890 102.110 224.260 ;
        RECT 104.040 223.890 134.560 224.260 ;
        RECT 0.130 223.505 2.420 223.845 ;
        RECT 3.165 223.505 4.650 223.845 ;
        RECT 0.130 222.870 0.730 223.505 ;
        RECT 0.130 222.640 1.860 222.870 ;
        RECT 2.160 222.640 3.820 222.870 ;
        RECT 0.130 220.630 0.730 222.640 ;
        RECT 2.160 221.605 2.390 222.640 ;
        RECT 2.795 221.350 3.025 222.395 ;
        RECT 4.050 221.350 4.650 223.505 ;
        RECT 6.690 223.170 37.210 223.550 ;
        RECT 39.140 223.170 69.660 223.550 ;
        RECT 71.590 223.170 102.110 223.550 ;
        RECT 104.040 223.170 134.560 223.550 ;
        RECT 5.840 222.915 6.460 223.100 ;
        RECT 37.440 222.915 38.060 223.100 ;
        RECT 5.840 222.685 38.060 222.915 ;
        RECT 5.840 222.500 6.460 222.685 ;
        RECT 37.440 222.500 38.060 222.685 ;
        RECT 38.290 222.915 38.910 223.100 ;
        RECT 69.890 222.915 70.510 223.100 ;
        RECT 38.290 222.685 70.510 222.915 ;
        RECT 38.290 222.500 38.910 222.685 ;
        RECT 69.890 222.500 70.510 222.685 ;
        RECT 70.740 222.915 71.360 223.100 ;
        RECT 102.340 222.915 102.960 223.100 ;
        RECT 70.740 222.685 102.960 222.915 ;
        RECT 70.740 222.500 71.360 222.685 ;
        RECT 102.340 222.500 102.960 222.685 ;
        RECT 103.190 222.915 103.810 223.100 ;
        RECT 134.790 222.915 135.410 223.100 ;
        RECT 103.190 222.685 135.410 222.915 ;
        RECT 103.190 222.500 103.810 222.685 ;
        RECT 134.790 222.500 135.410 222.685 ;
        RECT 10.400 222.420 12.020 222.430 ;
        RECT 42.850 222.420 44.470 222.430 ;
        RECT 75.300 222.420 76.920 222.430 ;
        RECT 107.750 222.420 109.370 222.430 ;
        RECT 6.690 222.050 37.210 222.420 ;
        RECT 39.140 222.050 69.660 222.420 ;
        RECT 71.590 222.050 102.110 222.420 ;
        RECT 104.040 222.050 134.560 222.420 ;
        RECT 0.960 221.120 3.025 221.350 ;
        RECT 3.255 221.120 4.650 221.350 ;
        RECT 6.690 221.330 37.210 221.710 ;
        RECT 39.140 221.330 69.660 221.710 ;
        RECT 71.590 221.330 102.110 221.710 ;
        RECT 104.040 221.330 134.560 221.710 ;
        RECT 0.130 220.400 1.860 220.630 ;
        RECT 2.160 220.400 3.820 220.630 ;
        RECT 0.130 218.245 0.730 220.400 ;
        RECT 2.160 219.365 2.390 220.400 ;
        RECT 2.795 219.110 3.025 220.155 ;
        RECT 4.050 219.110 4.650 221.120 ;
        RECT 5.840 221.075 6.460 221.260 ;
        RECT 37.440 221.075 38.060 221.260 ;
        RECT 5.840 220.845 38.060 221.075 ;
        RECT 5.840 220.660 6.460 220.845 ;
        RECT 37.440 220.660 38.060 220.845 ;
        RECT 38.290 221.075 38.910 221.260 ;
        RECT 69.890 221.075 70.510 221.260 ;
        RECT 38.290 220.845 70.510 221.075 ;
        RECT 38.290 220.660 38.910 220.845 ;
        RECT 69.890 220.660 70.510 220.845 ;
        RECT 70.740 221.075 71.360 221.260 ;
        RECT 102.340 221.075 102.960 221.260 ;
        RECT 70.740 220.845 102.960 221.075 ;
        RECT 70.740 220.660 71.360 220.845 ;
        RECT 102.340 220.660 102.960 220.845 ;
        RECT 103.190 221.075 103.810 221.260 ;
        RECT 134.790 221.075 135.410 221.260 ;
        RECT 103.190 220.845 135.410 221.075 ;
        RECT 103.190 220.660 103.810 220.845 ;
        RECT 134.790 220.660 135.410 220.845 ;
        RECT 6.690 220.210 37.210 220.580 ;
        RECT 39.140 220.210 69.660 220.580 ;
        RECT 71.590 220.210 102.110 220.580 ;
        RECT 104.040 220.210 134.560 220.580 ;
        RECT 0.960 218.880 3.025 219.110 ;
        RECT 3.255 218.880 4.650 219.110 ;
        RECT 4.050 218.245 4.650 218.880 ;
        RECT 0.130 217.905 2.420 218.245 ;
        RECT 3.165 217.905 4.650 218.245 ;
        RECT 0.130 217.270 0.730 217.905 ;
        RECT 0.130 217.040 1.710 217.270 ;
        RECT 0.130 215.000 0.730 217.040 ;
        RECT 2.140 216.810 2.500 216.895 ;
        RECT 1.010 216.580 2.500 216.810 ;
        RECT 1.010 216.430 1.370 216.580 ;
        RECT 0.960 215.795 1.910 216.200 ;
        RECT 0.130 214.770 1.420 215.000 ;
        RECT 0.130 213.810 0.730 214.770 ;
        RECT 1.650 214.450 1.910 215.795 ;
        RECT 2.140 215.145 2.500 216.580 ;
        RECT 2.730 215.245 3.080 216.445 ;
        RECT 3.440 215.835 3.820 217.480 ;
        RECT 2.520 214.450 2.870 214.510 ;
        RECT 3.440 214.450 3.780 215.055 ;
        RECT 1.650 214.190 3.780 214.450 ;
        RECT 2.520 214.130 2.870 214.190 ;
        RECT 4.050 213.910 4.650 217.905 ;
        RECT 6.495 217.425 8.245 220.210 ;
        RECT 8.885 217.425 9.695 218.425 ;
        RECT 10.335 217.425 12.085 219.720 ;
        RECT 12.725 217.425 13.535 218.425 ;
        RECT 14.175 217.425 15.925 219.720 ;
        RECT 16.565 217.425 17.375 218.425 ;
        RECT 18.015 217.425 19.765 219.720 ;
        RECT 20.405 217.425 21.215 218.425 ;
        RECT 21.855 217.425 23.605 219.720 ;
        RECT 24.245 217.425 25.055 218.425 ;
        RECT 25.695 217.425 27.445 219.720 ;
        RECT 28.085 217.425 28.895 218.425 ;
        RECT 29.535 217.425 31.285 219.720 ;
        RECT 31.925 217.425 32.735 218.425 ;
        RECT 33.375 217.425 35.125 219.720 ;
        RECT 35.765 217.425 36.575 218.425 ;
        RECT 38.945 217.425 40.695 220.210 ;
        RECT 41.335 217.425 42.145 218.425 ;
        RECT 42.785 217.425 44.535 219.720 ;
        RECT 45.175 217.425 45.985 218.425 ;
        RECT 46.625 217.425 48.375 219.720 ;
        RECT 49.015 217.425 49.825 218.425 ;
        RECT 50.465 217.425 52.215 219.720 ;
        RECT 52.855 217.425 53.665 218.425 ;
        RECT 54.305 217.425 56.055 219.720 ;
        RECT 56.695 217.425 57.505 218.425 ;
        RECT 58.145 217.425 59.895 219.720 ;
        RECT 60.535 217.425 61.345 218.425 ;
        RECT 61.985 217.425 63.735 219.720 ;
        RECT 64.375 217.425 65.185 218.425 ;
        RECT 65.825 217.425 67.575 219.720 ;
        RECT 68.215 217.425 69.025 218.425 ;
        RECT 71.395 217.425 73.145 220.210 ;
        RECT 73.785 217.425 74.595 218.425 ;
        RECT 75.235 217.425 76.985 219.720 ;
        RECT 77.625 217.425 78.435 218.425 ;
        RECT 79.075 217.425 80.825 219.720 ;
        RECT 81.465 217.425 82.275 218.425 ;
        RECT 82.915 217.425 84.665 219.720 ;
        RECT 85.305 217.425 86.115 218.425 ;
        RECT 86.755 217.425 88.505 219.720 ;
        RECT 89.145 217.425 89.955 218.425 ;
        RECT 90.595 217.425 92.345 219.720 ;
        RECT 92.985 217.425 93.795 218.425 ;
        RECT 94.435 217.425 96.185 219.720 ;
        RECT 96.825 217.425 97.635 218.425 ;
        RECT 98.275 217.425 100.025 219.720 ;
        RECT 100.665 217.425 101.475 218.425 ;
        RECT 103.845 217.425 105.595 220.210 ;
        RECT 106.235 217.425 107.045 218.425 ;
        RECT 107.685 217.425 109.435 219.720 ;
        RECT 110.075 217.425 110.885 218.425 ;
        RECT 111.525 217.425 113.275 219.720 ;
        RECT 113.915 217.425 114.725 218.425 ;
        RECT 115.365 217.425 117.115 219.720 ;
        RECT 117.755 217.425 118.565 218.425 ;
        RECT 119.205 217.425 120.955 219.720 ;
        RECT 121.595 217.425 122.405 218.425 ;
        RECT 123.045 217.425 124.795 219.720 ;
        RECT 125.435 217.425 126.245 218.425 ;
        RECT 126.885 217.425 128.635 219.720 ;
        RECT 129.275 217.425 130.085 218.425 ;
        RECT 130.725 217.425 132.475 219.720 ;
        RECT 133.115 217.425 133.925 218.425 ;
        RECT 136.340 217.615 136.710 236.125 ;
        RECT 137.360 232.490 137.730 236.125 ;
        RECT 137.355 232.110 137.735 232.490 ;
        RECT 137.360 229.490 137.730 232.110 ;
        RECT 137.355 229.110 137.735 229.490 ;
        RECT 137.360 226.490 137.730 229.110 ;
        RECT 137.355 226.110 137.735 226.490 ;
        RECT 137.360 223.490 137.730 226.110 ;
        RECT 137.355 223.110 137.735 223.490 ;
        RECT 137.360 220.490 137.730 223.110 ;
        RECT 137.355 220.110 137.735 220.490 ;
        RECT 136.340 217.235 136.720 217.615 ;
        RECT 136.340 216.165 136.710 217.235 ;
        RECT 6.965 214.975 7.775 215.975 ;
        RECT 0.130 213.580 1.820 213.810 ;
        RECT 3.190 213.680 4.650 213.910 ;
        RECT 0.130 211.570 0.730 213.580 ;
        RECT 2.150 213.120 3.150 213.445 ;
        RECT 0.960 212.560 3.820 212.890 ;
        RECT 0.130 211.340 1.820 211.570 ;
        RECT 0.130 209.330 0.730 211.340 ;
        RECT 2.535 211.205 2.800 212.560 ;
        RECT 4.050 211.670 4.650 213.680 ;
        RECT 8.415 213.145 10.165 215.975 ;
        RECT 10.805 214.975 11.615 215.975 ;
        RECT 12.255 213.680 14.005 215.975 ;
        RECT 14.645 214.975 15.455 215.975 ;
        RECT 16.095 213.680 17.845 215.975 ;
        RECT 18.485 214.975 19.295 215.975 ;
        RECT 19.935 213.680 21.685 215.975 ;
        RECT 22.325 214.975 23.135 215.975 ;
        RECT 23.775 213.680 25.525 215.975 ;
        RECT 26.165 214.975 26.975 215.975 ;
        RECT 27.615 213.680 29.365 215.975 ;
        RECT 30.005 214.975 30.815 215.975 ;
        RECT 31.455 213.680 33.205 215.975 ;
        RECT 33.845 214.975 34.655 215.975 ;
        RECT 35.295 213.680 37.045 215.975 ;
        RECT 39.415 214.975 40.225 215.975 ;
        RECT 40.865 213.145 42.615 215.975 ;
        RECT 43.255 214.975 44.065 215.975 ;
        RECT 44.705 213.680 46.455 215.975 ;
        RECT 47.095 214.975 47.905 215.975 ;
        RECT 48.545 213.680 50.295 215.975 ;
        RECT 50.935 214.975 51.745 215.975 ;
        RECT 52.385 213.680 54.135 215.975 ;
        RECT 54.775 214.975 55.585 215.975 ;
        RECT 56.225 213.680 57.975 215.975 ;
        RECT 58.615 214.975 59.425 215.975 ;
        RECT 60.065 213.680 61.815 215.975 ;
        RECT 62.455 214.975 63.265 215.975 ;
        RECT 63.905 213.680 65.655 215.975 ;
        RECT 66.295 214.975 67.105 215.975 ;
        RECT 67.745 213.680 69.495 215.975 ;
        RECT 71.865 214.975 72.675 215.975 ;
        RECT 73.315 213.145 75.065 215.975 ;
        RECT 75.705 214.975 76.515 215.975 ;
        RECT 77.155 213.680 78.905 215.975 ;
        RECT 79.545 214.975 80.355 215.975 ;
        RECT 80.995 213.680 82.745 215.975 ;
        RECT 83.385 214.975 84.195 215.975 ;
        RECT 84.835 213.680 86.585 215.975 ;
        RECT 87.225 214.975 88.035 215.975 ;
        RECT 88.675 213.680 90.425 215.975 ;
        RECT 91.065 214.975 91.875 215.975 ;
        RECT 92.515 213.680 94.265 215.975 ;
        RECT 94.905 214.975 95.715 215.975 ;
        RECT 96.355 213.680 98.105 215.975 ;
        RECT 98.745 214.975 99.555 215.975 ;
        RECT 100.195 213.680 101.945 215.975 ;
        RECT 104.315 214.975 105.125 215.975 ;
        RECT 105.765 213.145 107.515 215.975 ;
        RECT 108.155 214.975 108.965 215.975 ;
        RECT 109.605 213.680 111.355 215.975 ;
        RECT 111.995 214.975 112.805 215.975 ;
        RECT 113.445 213.680 115.195 215.975 ;
        RECT 115.835 214.975 116.645 215.975 ;
        RECT 117.285 213.680 119.035 215.975 ;
        RECT 119.675 214.975 120.485 215.975 ;
        RECT 121.125 213.680 122.875 215.975 ;
        RECT 123.515 214.975 124.325 215.975 ;
        RECT 124.965 213.680 126.715 215.975 ;
        RECT 127.355 214.975 128.165 215.975 ;
        RECT 128.805 213.680 130.555 215.975 ;
        RECT 131.195 214.975 132.005 215.975 ;
        RECT 132.645 213.680 134.395 215.975 ;
        RECT 136.340 215.785 136.720 216.165 ;
        RECT 6.690 212.775 37.210 213.145 ;
        RECT 39.140 212.775 69.660 213.145 ;
        RECT 71.590 212.775 102.110 213.145 ;
        RECT 104.040 212.775 134.560 213.145 ;
        RECT 5.840 212.510 6.460 212.695 ;
        RECT 37.440 212.510 38.060 212.695 ;
        RECT 5.840 212.280 38.060 212.510 ;
        RECT 5.840 212.095 6.460 212.280 ;
        RECT 37.440 212.095 38.060 212.280 ;
        RECT 38.290 212.510 38.910 212.695 ;
        RECT 69.890 212.510 70.510 212.695 ;
        RECT 38.290 212.280 70.510 212.510 ;
        RECT 38.290 212.095 38.910 212.280 ;
        RECT 69.890 212.095 70.510 212.280 ;
        RECT 70.740 212.510 71.360 212.695 ;
        RECT 102.340 212.510 102.960 212.695 ;
        RECT 70.740 212.280 102.960 212.510 ;
        RECT 70.740 212.095 71.360 212.280 ;
        RECT 102.340 212.095 102.960 212.280 ;
        RECT 103.190 212.510 103.810 212.695 ;
        RECT 134.790 212.510 135.410 212.695 ;
        RECT 103.190 212.280 135.410 212.510 ;
        RECT 103.190 212.095 103.810 212.280 ;
        RECT 134.790 212.095 135.410 212.280 ;
        RECT 3.190 211.440 4.650 211.670 ;
        RECT 6.690 211.645 37.210 212.025 ;
        RECT 39.140 211.645 69.660 212.025 ;
        RECT 71.590 211.645 102.110 212.025 ;
        RECT 104.040 211.645 134.560 212.025 ;
        RECT 2.150 210.880 3.150 211.205 ;
        RECT 0.960 210.320 3.820 210.650 ;
        RECT 4.050 209.430 4.650 211.440 ;
        RECT 6.690 210.935 37.210 211.305 ;
        RECT 39.140 210.935 69.660 211.305 ;
        RECT 71.590 210.935 102.110 211.305 ;
        RECT 104.040 210.935 134.560 211.305 ;
        RECT 12.320 210.925 13.940 210.935 ;
        RECT 44.770 210.925 46.390 210.935 ;
        RECT 77.220 210.925 78.840 210.935 ;
        RECT 109.670 210.925 111.290 210.935 ;
        RECT 5.840 210.670 6.460 210.855 ;
        RECT 37.440 210.670 38.060 210.855 ;
        RECT 5.840 210.440 38.060 210.670 ;
        RECT 5.840 210.255 6.460 210.440 ;
        RECT 37.440 210.255 38.060 210.440 ;
        RECT 38.290 210.670 38.910 210.855 ;
        RECT 69.890 210.670 70.510 210.855 ;
        RECT 38.290 210.440 70.510 210.670 ;
        RECT 38.290 210.255 38.910 210.440 ;
        RECT 69.890 210.255 70.510 210.440 ;
        RECT 70.740 210.670 71.360 210.855 ;
        RECT 102.340 210.670 102.960 210.855 ;
        RECT 70.740 210.440 102.960 210.670 ;
        RECT 70.740 210.255 71.360 210.440 ;
        RECT 102.340 210.255 102.960 210.440 ;
        RECT 103.190 210.670 103.810 210.855 ;
        RECT 134.790 210.670 135.410 210.855 ;
        RECT 103.190 210.440 135.410 210.670 ;
        RECT 103.190 210.255 103.810 210.440 ;
        RECT 134.790 210.255 135.410 210.440 ;
        RECT 6.690 209.805 37.210 210.185 ;
        RECT 39.140 209.805 69.660 210.185 ;
        RECT 71.590 209.805 102.110 210.185 ;
        RECT 104.040 209.805 134.560 210.185 ;
        RECT 0.130 209.100 1.820 209.330 ;
        RECT 3.190 209.200 4.650 209.430 ;
        RECT 0.130 207.045 0.730 209.100 ;
        RECT 2.150 208.640 3.150 208.965 ;
        RECT 0.960 208.080 3.820 208.410 ;
        RECT 2.300 207.955 2.680 208.080 ;
        RECT 4.050 207.045 4.650 209.200 ;
        RECT 6.690 209.090 37.210 209.460 ;
        RECT 39.140 209.090 69.660 209.460 ;
        RECT 71.590 209.090 102.110 209.460 ;
        RECT 104.040 209.090 134.560 209.460 ;
        RECT 16.160 209.080 17.780 209.090 ;
        RECT 48.610 209.080 50.230 209.090 ;
        RECT 81.060 209.080 82.680 209.090 ;
        RECT 113.510 209.080 115.130 209.090 ;
        RECT 5.840 208.825 6.460 209.010 ;
        RECT 37.440 208.825 38.060 209.010 ;
        RECT 5.840 208.595 38.060 208.825 ;
        RECT 5.840 208.410 6.460 208.595 ;
        RECT 37.440 208.410 38.060 208.595 ;
        RECT 38.290 208.825 38.910 209.010 ;
        RECT 69.890 208.825 70.510 209.010 ;
        RECT 38.290 208.595 70.510 208.825 ;
        RECT 38.290 208.410 38.910 208.595 ;
        RECT 69.890 208.410 70.510 208.595 ;
        RECT 70.740 208.825 71.360 209.010 ;
        RECT 102.340 208.825 102.960 209.010 ;
        RECT 70.740 208.595 102.960 208.825 ;
        RECT 70.740 208.410 71.360 208.595 ;
        RECT 102.340 208.410 102.960 208.595 ;
        RECT 103.190 208.825 103.810 209.010 ;
        RECT 134.790 208.825 135.410 209.010 ;
        RECT 103.190 208.595 135.410 208.825 ;
        RECT 103.190 208.410 103.810 208.595 ;
        RECT 134.790 208.410 135.410 208.595 ;
        RECT 6.690 207.960 37.210 208.340 ;
        RECT 39.140 207.960 69.660 208.340 ;
        RECT 71.590 207.960 102.110 208.340 ;
        RECT 104.040 207.960 134.560 208.340 ;
        RECT 6.700 207.170 37.200 207.610 ;
        RECT 39.150 207.170 69.650 207.610 ;
        RECT 71.600 207.170 102.100 207.610 ;
        RECT 104.050 207.170 134.550 207.610 ;
        RECT 0.130 206.705 2.420 207.045 ;
        RECT 3.165 206.705 4.650 207.045 ;
        RECT 0.130 205.925 0.730 206.705 ;
        RECT 4.050 205.925 4.650 206.705 ;
        RECT 6.690 206.450 37.210 206.820 ;
        RECT 39.140 206.450 69.660 206.820 ;
        RECT 71.590 206.450 102.110 206.820 ;
        RECT 104.040 206.450 134.560 206.820 ;
        RECT 20.000 206.440 21.620 206.450 ;
        RECT 52.450 206.440 54.070 206.450 ;
        RECT 84.900 206.440 86.520 206.450 ;
        RECT 117.350 206.440 118.970 206.450 ;
        RECT 0.130 205.585 2.420 205.925 ;
        RECT 3.165 205.585 4.650 205.925 ;
        RECT 5.840 206.185 6.460 206.370 ;
        RECT 37.440 206.185 38.060 206.370 ;
        RECT 5.840 205.955 38.060 206.185 ;
        RECT 5.840 205.770 6.460 205.955 ;
        RECT 37.440 205.770 38.060 205.955 ;
        RECT 38.290 206.185 38.910 206.370 ;
        RECT 69.890 206.185 70.510 206.370 ;
        RECT 38.290 205.955 70.510 206.185 ;
        RECT 38.290 205.770 38.910 205.955 ;
        RECT 69.890 205.770 70.510 205.955 ;
        RECT 70.740 206.185 71.360 206.370 ;
        RECT 102.340 206.185 102.960 206.370 ;
        RECT 70.740 205.955 102.960 206.185 ;
        RECT 70.740 205.770 71.360 205.955 ;
        RECT 102.340 205.770 102.960 205.955 ;
        RECT 103.190 206.185 103.810 206.370 ;
        RECT 134.790 206.185 135.410 206.370 ;
        RECT 103.190 205.955 135.410 206.185 ;
        RECT 103.190 205.770 103.810 205.955 ;
        RECT 134.790 205.770 135.410 205.955 ;
        RECT 0.130 204.950 0.730 205.585 ;
        RECT 0.130 204.720 1.860 204.950 ;
        RECT 2.160 204.720 3.820 204.950 ;
        RECT 0.130 202.710 0.730 204.720 ;
        RECT 2.160 203.685 2.390 204.720 ;
        RECT 2.795 203.430 3.025 204.475 ;
        RECT 4.050 203.430 4.650 205.585 ;
        RECT 6.690 205.320 37.210 205.700 ;
        RECT 39.140 205.320 69.660 205.700 ;
        RECT 71.590 205.320 102.110 205.700 ;
        RECT 104.040 205.320 134.560 205.700 ;
        RECT 6.690 204.610 37.210 204.980 ;
        RECT 39.140 204.610 69.660 204.980 ;
        RECT 71.590 204.610 102.110 204.980 ;
        RECT 104.040 204.610 134.560 204.980 ;
        RECT 23.840 204.600 25.460 204.610 ;
        RECT 56.290 204.600 57.910 204.610 ;
        RECT 88.740 204.600 90.360 204.610 ;
        RECT 121.190 204.600 122.810 204.610 ;
        RECT 5.840 204.345 6.460 204.530 ;
        RECT 37.440 204.345 38.060 204.530 ;
        RECT 5.840 204.115 38.060 204.345 ;
        RECT 5.840 203.930 6.460 204.115 ;
        RECT 37.440 203.930 38.060 204.115 ;
        RECT 38.290 204.345 38.910 204.530 ;
        RECT 69.890 204.345 70.510 204.530 ;
        RECT 38.290 204.115 70.510 204.345 ;
        RECT 38.290 203.930 38.910 204.115 ;
        RECT 69.890 203.930 70.510 204.115 ;
        RECT 70.740 204.345 71.360 204.530 ;
        RECT 102.340 204.345 102.960 204.530 ;
        RECT 70.740 204.115 102.960 204.345 ;
        RECT 70.740 203.930 71.360 204.115 ;
        RECT 102.340 203.930 102.960 204.115 ;
        RECT 103.190 204.345 103.810 204.530 ;
        RECT 134.790 204.345 135.410 204.530 ;
        RECT 103.190 204.115 135.410 204.345 ;
        RECT 103.190 203.930 103.810 204.115 ;
        RECT 134.790 203.930 135.410 204.115 ;
        RECT 6.690 203.480 37.210 203.860 ;
        RECT 39.140 203.480 69.660 203.860 ;
        RECT 71.590 203.480 102.110 203.860 ;
        RECT 104.040 203.480 134.560 203.860 ;
        RECT 0.960 203.200 3.025 203.430 ;
        RECT 3.255 203.200 4.650 203.430 ;
        RECT 0.130 202.480 1.860 202.710 ;
        RECT 2.160 202.480 3.820 202.710 ;
        RECT 0.130 200.470 0.730 202.480 ;
        RECT 2.160 201.445 2.390 202.480 ;
        RECT 2.795 201.190 3.025 202.235 ;
        RECT 4.050 201.190 4.650 203.200 ;
        RECT 6.690 202.765 37.210 203.135 ;
        RECT 39.140 202.765 69.660 203.135 ;
        RECT 71.590 202.765 102.110 203.135 ;
        RECT 104.040 202.765 134.560 203.135 ;
        RECT 27.680 202.755 29.300 202.765 ;
        RECT 60.130 202.755 61.750 202.765 ;
        RECT 92.580 202.755 94.200 202.765 ;
        RECT 125.030 202.755 126.650 202.765 ;
        RECT 5.840 202.500 6.460 202.685 ;
        RECT 37.440 202.500 38.060 202.685 ;
        RECT 5.840 202.270 38.060 202.500 ;
        RECT 5.840 202.085 6.460 202.270 ;
        RECT 37.440 202.085 38.060 202.270 ;
        RECT 38.290 202.500 38.910 202.685 ;
        RECT 69.890 202.500 70.510 202.685 ;
        RECT 38.290 202.270 70.510 202.500 ;
        RECT 38.290 202.085 38.910 202.270 ;
        RECT 69.890 202.085 70.510 202.270 ;
        RECT 70.740 202.500 71.360 202.685 ;
        RECT 102.340 202.500 102.960 202.685 ;
        RECT 70.740 202.270 102.960 202.500 ;
        RECT 70.740 202.085 71.360 202.270 ;
        RECT 102.340 202.085 102.960 202.270 ;
        RECT 103.190 202.500 103.810 202.685 ;
        RECT 134.790 202.500 135.410 202.685 ;
        RECT 103.190 202.270 135.410 202.500 ;
        RECT 103.190 202.085 103.810 202.270 ;
        RECT 134.790 202.085 135.410 202.270 ;
        RECT 6.690 201.635 37.210 202.015 ;
        RECT 39.140 201.635 69.660 202.015 ;
        RECT 71.590 201.635 102.110 202.015 ;
        RECT 104.040 201.635 134.560 202.015 ;
        RECT 0.960 200.960 3.025 201.190 ;
        RECT 3.255 200.960 4.650 201.190 ;
        RECT 0.130 200.240 1.860 200.470 ;
        RECT 2.160 200.240 3.820 200.470 ;
        RECT 0.130 198.065 0.730 200.240 ;
        RECT 2.160 199.205 2.390 200.240 ;
        RECT 2.795 198.950 3.025 199.995 ;
        RECT 4.050 198.950 4.650 200.960 ;
        RECT 6.700 200.845 37.200 201.285 ;
        RECT 39.150 200.845 69.650 201.285 ;
        RECT 71.600 200.845 102.100 201.285 ;
        RECT 104.050 200.845 134.550 201.285 ;
        RECT 6.690 200.125 37.210 200.495 ;
        RECT 39.140 200.125 69.660 200.495 ;
        RECT 71.590 200.125 102.110 200.495 ;
        RECT 104.040 200.125 134.560 200.495 ;
        RECT 31.520 200.115 33.140 200.125 ;
        RECT 63.970 200.115 65.590 200.125 ;
        RECT 96.420 200.115 98.040 200.125 ;
        RECT 128.870 200.115 130.490 200.125 ;
        RECT 5.840 199.860 6.460 200.045 ;
        RECT 37.440 199.860 38.060 200.045 ;
        RECT 5.840 199.630 38.060 199.860 ;
        RECT 5.840 199.445 6.460 199.630 ;
        RECT 37.440 199.445 38.060 199.630 ;
        RECT 38.290 199.860 38.910 200.045 ;
        RECT 69.890 199.860 70.510 200.045 ;
        RECT 38.290 199.630 70.510 199.860 ;
        RECT 38.290 199.445 38.910 199.630 ;
        RECT 69.890 199.445 70.510 199.630 ;
        RECT 70.740 199.860 71.360 200.045 ;
        RECT 102.340 199.860 102.960 200.045 ;
        RECT 70.740 199.630 102.960 199.860 ;
        RECT 70.740 199.445 71.360 199.630 ;
        RECT 102.340 199.445 102.960 199.630 ;
        RECT 103.190 199.860 103.810 200.045 ;
        RECT 134.790 199.860 135.410 200.045 ;
        RECT 103.190 199.630 135.410 199.860 ;
        RECT 103.190 199.445 103.810 199.630 ;
        RECT 134.790 199.445 135.410 199.630 ;
        RECT 6.690 198.995 37.210 199.375 ;
        RECT 39.140 198.995 69.660 199.375 ;
        RECT 71.590 198.995 102.110 199.375 ;
        RECT 104.040 198.995 134.560 199.375 ;
        RECT 0.960 198.720 3.025 198.950 ;
        RECT 3.255 198.720 4.650 198.950 ;
        RECT 4.050 198.065 4.650 198.720 ;
        RECT 6.690 198.285 37.210 198.655 ;
        RECT 39.140 198.285 69.660 198.655 ;
        RECT 71.590 198.285 102.110 198.655 ;
        RECT 104.040 198.285 134.560 198.655 ;
        RECT 35.360 198.275 36.980 198.285 ;
        RECT 67.810 198.275 69.430 198.285 ;
        RECT 100.260 198.275 101.880 198.285 ;
        RECT 132.710 198.275 134.330 198.285 ;
        RECT 0.130 197.725 2.430 198.065 ;
        RECT 3.160 197.725 4.650 198.065 ;
        RECT 0.130 196.760 0.730 197.725 ;
        RECT 4.050 196.760 4.650 197.725 ;
        RECT 5.840 198.020 6.460 198.205 ;
        RECT 37.440 198.020 38.060 198.205 ;
        RECT 5.840 197.790 38.060 198.020 ;
        RECT 5.840 197.605 6.460 197.790 ;
        RECT 37.440 197.605 38.060 197.790 ;
        RECT 38.290 198.020 38.910 198.205 ;
        RECT 69.890 198.020 70.510 198.205 ;
        RECT 38.290 197.790 70.510 198.020 ;
        RECT 38.290 197.605 38.910 197.790 ;
        RECT 69.890 197.605 70.510 197.790 ;
        RECT 70.740 198.020 71.360 198.205 ;
        RECT 102.340 198.020 102.960 198.205 ;
        RECT 70.740 197.790 102.960 198.020 ;
        RECT 70.740 197.605 71.360 197.790 ;
        RECT 102.340 197.605 102.960 197.790 ;
        RECT 103.190 198.020 103.810 198.205 ;
        RECT 134.790 198.020 135.410 198.205 ;
        RECT 103.190 197.790 135.410 198.020 ;
        RECT 136.340 197.855 136.710 215.785 ;
        RECT 137.360 214.490 137.730 220.110 ;
        RECT 138.380 217.615 138.750 236.125 ;
        RECT 139.400 232.490 139.770 236.125 ;
        RECT 139.395 232.110 139.775 232.490 ;
        RECT 139.400 229.490 139.770 232.110 ;
        RECT 139.395 229.110 139.775 229.490 ;
        RECT 139.400 226.490 139.770 229.110 ;
        RECT 139.395 226.110 139.775 226.490 ;
        RECT 139.400 223.490 139.770 226.110 ;
        RECT 139.395 223.110 139.775 223.490 ;
        RECT 139.400 220.490 139.770 223.110 ;
        RECT 139.395 220.110 139.775 220.490 ;
        RECT 138.380 217.235 138.760 217.615 ;
        RECT 138.380 216.165 138.750 217.235 ;
        RECT 138.380 215.785 138.760 216.165 ;
        RECT 137.355 214.110 137.735 214.490 ;
        RECT 137.360 211.490 137.730 214.110 ;
        RECT 137.355 211.110 137.735 211.490 ;
        RECT 137.360 208.490 137.730 211.110 ;
        RECT 137.355 208.110 137.735 208.490 ;
        RECT 137.360 205.490 137.730 208.110 ;
        RECT 137.355 205.110 137.735 205.490 ;
        RECT 137.360 202.490 137.730 205.110 ;
        RECT 137.355 202.110 137.735 202.490 ;
        RECT 137.360 199.490 137.730 202.110 ;
        RECT 137.355 199.110 137.735 199.490 ;
        RECT 137.360 197.855 137.730 199.110 ;
        RECT 138.380 197.855 138.750 215.785 ;
        RECT 139.400 214.490 139.770 220.110 ;
        RECT 139.395 214.110 139.775 214.490 ;
        RECT 139.400 211.490 139.770 214.110 ;
        RECT 139.395 211.110 139.775 211.490 ;
        RECT 139.400 208.490 139.770 211.110 ;
        RECT 139.395 208.110 139.775 208.490 ;
        RECT 139.400 205.490 139.770 208.110 ;
        RECT 139.395 205.110 139.775 205.490 ;
        RECT 139.400 202.490 139.770 205.110 ;
        RECT 139.395 202.110 139.775 202.490 ;
        RECT 139.400 199.490 139.770 202.110 ;
        RECT 139.395 199.110 139.775 199.490 ;
        RECT 139.400 197.855 139.770 199.110 ;
        RECT 140.420 197.855 140.800 236.125 ;
        RECT 141.150 197.865 141.590 236.115 ;
        RECT 103.190 197.605 103.810 197.790 ;
        RECT 134.790 197.605 135.410 197.790 ;
        RECT 6.690 197.155 37.210 197.535 ;
        RECT 39.140 197.155 69.660 197.535 ;
        RECT 71.590 197.155 102.110 197.535 ;
        RECT 104.040 197.155 134.560 197.535 ;
        RECT 0.130 196.420 2.430 196.760 ;
        RECT 3.160 196.420 4.650 196.760 ;
        RECT 6.690 196.435 37.210 196.815 ;
        RECT 39.140 196.435 69.660 196.815 ;
        RECT 71.590 196.435 102.110 196.815 ;
        RECT 104.040 196.435 134.560 196.815 ;
        RECT 0.130 195.805 0.730 196.420 ;
        RECT 0.130 195.575 1.860 195.805 ;
        RECT 2.160 195.575 3.820 195.805 ;
        RECT 0.130 193.565 0.730 195.575 ;
        RECT 2.160 194.540 2.390 195.575 ;
        RECT 2.795 194.285 3.025 195.330 ;
        RECT 4.050 194.285 4.650 196.420 ;
        RECT 5.840 196.180 6.460 196.365 ;
        RECT 37.440 196.180 38.060 196.365 ;
        RECT 5.840 195.950 38.060 196.180 ;
        RECT 5.840 195.765 6.460 195.950 ;
        RECT 37.440 195.765 38.060 195.950 ;
        RECT 38.290 196.180 38.910 196.365 ;
        RECT 69.890 196.180 70.510 196.365 ;
        RECT 38.290 195.950 70.510 196.180 ;
        RECT 38.290 195.765 38.910 195.950 ;
        RECT 69.890 195.765 70.510 195.950 ;
        RECT 70.740 196.180 71.360 196.365 ;
        RECT 102.340 196.180 102.960 196.365 ;
        RECT 70.740 195.950 102.960 196.180 ;
        RECT 70.740 195.765 71.360 195.950 ;
        RECT 102.340 195.765 102.960 195.950 ;
        RECT 103.190 196.180 103.810 196.365 ;
        RECT 134.790 196.180 135.410 196.365 ;
        RECT 103.190 195.950 135.410 196.180 ;
        RECT 103.190 195.765 103.810 195.950 ;
        RECT 134.790 195.765 135.410 195.950 ;
        RECT 33.440 195.685 35.060 195.695 ;
        RECT 65.890 195.685 67.510 195.695 ;
        RECT 98.340 195.685 99.960 195.695 ;
        RECT 130.790 195.685 132.410 195.695 ;
        RECT 6.690 195.315 37.210 195.685 ;
        RECT 39.140 195.315 69.660 195.685 ;
        RECT 71.590 195.315 102.110 195.685 ;
        RECT 104.040 195.315 134.560 195.685 ;
        RECT 6.690 194.595 37.210 194.975 ;
        RECT 39.140 194.595 69.660 194.975 ;
        RECT 71.590 194.595 102.110 194.975 ;
        RECT 104.040 194.595 134.560 194.975 ;
        RECT 0.960 194.055 3.025 194.285 ;
        RECT 3.255 194.055 4.650 194.285 ;
        RECT 0.130 193.335 1.860 193.565 ;
        RECT 2.160 193.335 3.820 193.565 ;
        RECT 0.130 191.325 0.730 193.335 ;
        RECT 2.160 192.300 2.390 193.335 ;
        RECT 2.795 192.045 3.025 193.090 ;
        RECT 4.050 192.045 4.650 194.055 ;
        RECT 5.840 194.340 6.460 194.525 ;
        RECT 37.440 194.340 38.060 194.525 ;
        RECT 5.840 194.110 38.060 194.340 ;
        RECT 5.840 193.925 6.460 194.110 ;
        RECT 37.440 193.925 38.060 194.110 ;
        RECT 38.290 194.340 38.910 194.525 ;
        RECT 69.890 194.340 70.510 194.525 ;
        RECT 38.290 194.110 70.510 194.340 ;
        RECT 38.290 193.925 38.910 194.110 ;
        RECT 69.890 193.925 70.510 194.110 ;
        RECT 70.740 194.340 71.360 194.525 ;
        RECT 102.340 194.340 102.960 194.525 ;
        RECT 70.740 194.110 102.960 194.340 ;
        RECT 70.740 193.925 71.360 194.110 ;
        RECT 102.340 193.925 102.960 194.110 ;
        RECT 103.190 194.340 103.810 194.525 ;
        RECT 134.790 194.340 135.410 194.525 ;
        RECT 103.190 194.110 135.410 194.340 ;
        RECT 103.190 193.925 103.810 194.110 ;
        RECT 134.790 193.925 135.410 194.110 ;
        RECT 29.600 193.845 31.220 193.855 ;
        RECT 62.050 193.845 63.670 193.855 ;
        RECT 94.500 193.845 96.120 193.855 ;
        RECT 126.950 193.845 128.570 193.855 ;
        RECT 6.690 193.475 37.210 193.845 ;
        RECT 39.140 193.475 69.660 193.845 ;
        RECT 71.590 193.475 102.110 193.845 ;
        RECT 104.040 193.475 134.560 193.845 ;
        RECT 6.700 192.680 37.200 193.120 ;
        RECT 39.150 192.680 69.650 193.120 ;
        RECT 71.600 192.680 102.100 193.120 ;
        RECT 104.050 192.680 134.550 193.120 ;
        RECT 0.960 191.815 3.025 192.045 ;
        RECT 3.255 191.815 4.650 192.045 ;
        RECT 6.690 191.950 37.210 192.330 ;
        RECT 39.140 191.950 69.660 192.330 ;
        RECT 71.590 191.950 102.110 192.330 ;
        RECT 104.040 191.950 134.560 192.330 ;
        RECT 0.130 191.095 1.860 191.325 ;
        RECT 2.160 191.095 3.820 191.325 ;
        RECT 0.130 189.085 0.730 191.095 ;
        RECT 2.160 190.060 2.390 191.095 ;
        RECT 2.795 189.805 3.025 190.850 ;
        RECT 4.050 189.805 4.650 191.815 ;
        RECT 5.840 191.695 6.460 191.880 ;
        RECT 37.440 191.695 38.060 191.880 ;
        RECT 5.840 191.465 38.060 191.695 ;
        RECT 5.840 191.280 6.460 191.465 ;
        RECT 37.440 191.280 38.060 191.465 ;
        RECT 38.290 191.695 38.910 191.880 ;
        RECT 69.890 191.695 70.510 191.880 ;
        RECT 38.290 191.465 70.510 191.695 ;
        RECT 38.290 191.280 38.910 191.465 ;
        RECT 69.890 191.280 70.510 191.465 ;
        RECT 70.740 191.695 71.360 191.880 ;
        RECT 102.340 191.695 102.960 191.880 ;
        RECT 70.740 191.465 102.960 191.695 ;
        RECT 70.740 191.280 71.360 191.465 ;
        RECT 102.340 191.280 102.960 191.465 ;
        RECT 103.190 191.695 103.810 191.880 ;
        RECT 134.790 191.695 135.410 191.880 ;
        RECT 103.190 191.465 135.410 191.695 ;
        RECT 103.190 191.280 103.810 191.465 ;
        RECT 134.790 191.280 135.410 191.465 ;
        RECT 25.760 191.200 27.380 191.210 ;
        RECT 58.210 191.200 59.830 191.210 ;
        RECT 90.660 191.200 92.280 191.210 ;
        RECT 123.110 191.200 124.730 191.210 ;
        RECT 6.690 190.830 37.210 191.200 ;
        RECT 39.140 190.830 69.660 191.200 ;
        RECT 71.590 190.830 102.110 191.200 ;
        RECT 104.040 190.830 134.560 191.200 ;
        RECT 6.690 190.110 37.210 190.490 ;
        RECT 39.140 190.110 69.660 190.490 ;
        RECT 71.590 190.110 102.110 190.490 ;
        RECT 104.040 190.110 134.560 190.490 ;
        RECT 0.960 189.575 3.025 189.805 ;
        RECT 3.255 189.575 4.650 189.805 ;
        RECT 0.130 188.855 1.860 189.085 ;
        RECT 2.160 188.855 3.820 189.085 ;
        RECT 0.130 186.845 0.730 188.855 ;
        RECT 2.160 187.820 2.390 188.855 ;
        RECT 2.795 187.565 3.025 188.610 ;
        RECT 4.050 187.565 4.650 189.575 ;
        RECT 5.840 189.855 6.460 190.040 ;
        RECT 37.440 189.855 38.060 190.040 ;
        RECT 5.840 189.625 38.060 189.855 ;
        RECT 5.840 189.440 6.460 189.625 ;
        RECT 37.440 189.440 38.060 189.625 ;
        RECT 38.290 189.855 38.910 190.040 ;
        RECT 69.890 189.855 70.510 190.040 ;
        RECT 38.290 189.625 70.510 189.855 ;
        RECT 38.290 189.440 38.910 189.625 ;
        RECT 69.890 189.440 70.510 189.625 ;
        RECT 70.740 189.855 71.360 190.040 ;
        RECT 102.340 189.855 102.960 190.040 ;
        RECT 70.740 189.625 102.960 189.855 ;
        RECT 70.740 189.440 71.360 189.625 ;
        RECT 102.340 189.440 102.960 189.625 ;
        RECT 103.190 189.855 103.810 190.040 ;
        RECT 134.790 189.855 135.410 190.040 ;
        RECT 103.190 189.625 135.410 189.855 ;
        RECT 103.190 189.440 103.810 189.625 ;
        RECT 134.790 189.440 135.410 189.625 ;
        RECT 21.920 189.360 23.540 189.370 ;
        RECT 54.370 189.360 55.990 189.370 ;
        RECT 86.820 189.360 88.440 189.370 ;
        RECT 119.270 189.360 120.890 189.370 ;
        RECT 6.690 188.990 37.210 189.360 ;
        RECT 39.140 188.990 69.660 189.360 ;
        RECT 71.590 188.990 102.110 189.360 ;
        RECT 104.040 188.990 134.560 189.360 ;
        RECT 6.690 188.270 37.210 188.650 ;
        RECT 39.140 188.270 69.660 188.650 ;
        RECT 71.590 188.270 102.110 188.650 ;
        RECT 104.040 188.270 134.560 188.650 ;
        RECT 5.840 188.015 6.460 188.200 ;
        RECT 37.440 188.015 38.060 188.200 ;
        RECT 5.840 187.785 38.060 188.015 ;
        RECT 5.840 187.600 6.460 187.785 ;
        RECT 37.440 187.600 38.060 187.785 ;
        RECT 38.290 188.015 38.910 188.200 ;
        RECT 69.890 188.015 70.510 188.200 ;
        RECT 38.290 187.785 70.510 188.015 ;
        RECT 38.290 187.600 38.910 187.785 ;
        RECT 69.890 187.600 70.510 187.785 ;
        RECT 70.740 188.015 71.360 188.200 ;
        RECT 102.340 188.015 102.960 188.200 ;
        RECT 70.740 187.785 102.960 188.015 ;
        RECT 70.740 187.600 71.360 187.785 ;
        RECT 102.340 187.600 102.960 187.785 ;
        RECT 103.190 188.015 103.810 188.200 ;
        RECT 134.790 188.015 135.410 188.200 ;
        RECT 103.190 187.785 135.410 188.015 ;
        RECT 103.190 187.600 103.810 187.785 ;
        RECT 134.790 187.600 135.410 187.785 ;
        RECT 0.960 187.335 3.025 187.565 ;
        RECT 3.255 187.335 4.650 187.565 ;
        RECT 18.080 187.520 19.700 187.530 ;
        RECT 50.530 187.520 52.150 187.530 ;
        RECT 82.980 187.520 84.600 187.530 ;
        RECT 115.430 187.520 117.050 187.530 ;
        RECT 0.130 186.615 1.860 186.845 ;
        RECT 2.160 186.615 3.820 186.845 ;
        RECT 0.130 184.460 0.730 186.615 ;
        RECT 2.160 185.580 2.390 186.615 ;
        RECT 2.795 185.325 3.025 186.370 ;
        RECT 4.050 185.325 4.650 187.335 ;
        RECT 6.690 187.150 37.210 187.520 ;
        RECT 39.140 187.150 69.660 187.520 ;
        RECT 71.590 187.150 102.110 187.520 ;
        RECT 104.040 187.150 134.560 187.520 ;
        RECT 6.700 186.355 37.200 186.795 ;
        RECT 39.150 186.355 69.650 186.795 ;
        RECT 71.600 186.355 102.100 186.795 ;
        RECT 104.050 186.355 134.550 186.795 ;
        RECT 6.690 185.625 37.210 186.005 ;
        RECT 39.140 185.625 69.660 186.005 ;
        RECT 71.590 185.625 102.110 186.005 ;
        RECT 104.040 185.625 134.560 186.005 ;
        RECT 0.960 185.095 3.025 185.325 ;
        RECT 3.255 185.095 4.650 185.325 ;
        RECT 4.050 184.460 4.650 185.095 ;
        RECT 5.840 185.370 6.460 185.555 ;
        RECT 37.440 185.370 38.060 185.555 ;
        RECT 5.840 185.140 38.060 185.370 ;
        RECT 5.840 184.955 6.460 185.140 ;
        RECT 37.440 184.955 38.060 185.140 ;
        RECT 38.290 185.370 38.910 185.555 ;
        RECT 69.890 185.370 70.510 185.555 ;
        RECT 38.290 185.140 70.510 185.370 ;
        RECT 38.290 184.955 38.910 185.140 ;
        RECT 69.890 184.955 70.510 185.140 ;
        RECT 70.740 185.370 71.360 185.555 ;
        RECT 102.340 185.370 102.960 185.555 ;
        RECT 70.740 185.140 102.960 185.370 ;
        RECT 70.740 184.955 71.360 185.140 ;
        RECT 102.340 184.955 102.960 185.140 ;
        RECT 103.190 185.370 103.810 185.555 ;
        RECT 134.790 185.370 135.410 185.555 ;
        RECT 103.190 185.140 135.410 185.370 ;
        RECT 103.190 184.955 103.810 185.140 ;
        RECT 134.790 184.955 135.410 185.140 ;
        RECT 14.240 184.875 15.860 184.885 ;
        RECT 46.690 184.875 48.310 184.885 ;
        RECT 79.140 184.875 80.760 184.885 ;
        RECT 111.590 184.875 113.210 184.885 ;
        RECT 6.690 184.505 37.210 184.875 ;
        RECT 39.140 184.505 69.660 184.875 ;
        RECT 71.590 184.505 102.110 184.875 ;
        RECT 104.040 184.505 134.560 184.875 ;
        RECT 0.130 184.120 2.420 184.460 ;
        RECT 3.165 184.120 4.650 184.460 ;
        RECT 0.130 183.485 0.730 184.120 ;
        RECT 0.130 183.255 1.860 183.485 ;
        RECT 2.160 183.255 3.820 183.485 ;
        RECT 0.130 181.245 0.730 183.255 ;
        RECT 2.160 182.220 2.390 183.255 ;
        RECT 2.795 181.965 3.025 183.010 ;
        RECT 4.050 181.965 4.650 184.120 ;
        RECT 6.690 183.785 37.210 184.165 ;
        RECT 39.140 183.785 69.660 184.165 ;
        RECT 71.590 183.785 102.110 184.165 ;
        RECT 104.040 183.785 134.560 184.165 ;
        RECT 5.840 183.530 6.460 183.715 ;
        RECT 37.440 183.530 38.060 183.715 ;
        RECT 5.840 183.300 38.060 183.530 ;
        RECT 5.840 183.115 6.460 183.300 ;
        RECT 37.440 183.115 38.060 183.300 ;
        RECT 38.290 183.530 38.910 183.715 ;
        RECT 69.890 183.530 70.510 183.715 ;
        RECT 38.290 183.300 70.510 183.530 ;
        RECT 38.290 183.115 38.910 183.300 ;
        RECT 69.890 183.115 70.510 183.300 ;
        RECT 70.740 183.530 71.360 183.715 ;
        RECT 102.340 183.530 102.960 183.715 ;
        RECT 70.740 183.300 102.960 183.530 ;
        RECT 70.740 183.115 71.360 183.300 ;
        RECT 102.340 183.115 102.960 183.300 ;
        RECT 103.190 183.530 103.810 183.715 ;
        RECT 134.790 183.530 135.410 183.715 ;
        RECT 103.190 183.300 135.410 183.530 ;
        RECT 103.190 183.115 103.810 183.300 ;
        RECT 134.790 183.115 135.410 183.300 ;
        RECT 10.400 183.035 12.020 183.045 ;
        RECT 42.850 183.035 44.470 183.045 ;
        RECT 75.300 183.035 76.920 183.045 ;
        RECT 107.750 183.035 109.370 183.045 ;
        RECT 6.690 182.665 37.210 183.035 ;
        RECT 39.140 182.665 69.660 183.035 ;
        RECT 71.590 182.665 102.110 183.035 ;
        RECT 104.040 182.665 134.560 183.035 ;
        RECT 0.960 181.735 3.025 181.965 ;
        RECT 3.255 181.735 4.650 181.965 ;
        RECT 6.690 181.945 37.210 182.325 ;
        RECT 39.140 181.945 69.660 182.325 ;
        RECT 71.590 181.945 102.110 182.325 ;
        RECT 104.040 181.945 134.560 182.325 ;
        RECT 0.130 181.015 1.860 181.245 ;
        RECT 2.160 181.015 3.820 181.245 ;
        RECT 0.130 178.860 0.730 181.015 ;
        RECT 2.160 179.980 2.390 181.015 ;
        RECT 2.795 179.725 3.025 180.770 ;
        RECT 4.050 179.725 4.650 181.735 ;
        RECT 5.840 181.690 6.460 181.875 ;
        RECT 37.440 181.690 38.060 181.875 ;
        RECT 5.840 181.460 38.060 181.690 ;
        RECT 5.840 181.275 6.460 181.460 ;
        RECT 37.440 181.275 38.060 181.460 ;
        RECT 38.290 181.690 38.910 181.875 ;
        RECT 69.890 181.690 70.510 181.875 ;
        RECT 38.290 181.460 70.510 181.690 ;
        RECT 38.290 181.275 38.910 181.460 ;
        RECT 69.890 181.275 70.510 181.460 ;
        RECT 70.740 181.690 71.360 181.875 ;
        RECT 102.340 181.690 102.960 181.875 ;
        RECT 70.740 181.460 102.960 181.690 ;
        RECT 70.740 181.275 71.360 181.460 ;
        RECT 102.340 181.275 102.960 181.460 ;
        RECT 103.190 181.690 103.810 181.875 ;
        RECT 134.790 181.690 135.410 181.875 ;
        RECT 103.190 181.460 135.410 181.690 ;
        RECT 103.190 181.275 103.810 181.460 ;
        RECT 134.790 181.275 135.410 181.460 ;
        RECT 6.690 180.825 37.210 181.195 ;
        RECT 39.140 180.825 69.660 181.195 ;
        RECT 71.590 180.825 102.110 181.195 ;
        RECT 104.040 180.825 134.560 181.195 ;
        RECT 0.960 179.495 3.025 179.725 ;
        RECT 3.255 179.495 4.650 179.725 ;
        RECT 4.050 178.860 4.650 179.495 ;
        RECT 0.130 178.520 2.420 178.860 ;
        RECT 3.165 178.520 4.650 178.860 ;
        RECT 0.130 177.885 0.730 178.520 ;
        RECT 0.130 177.655 1.710 177.885 ;
        RECT 0.130 175.615 0.730 177.655 ;
        RECT 2.140 177.425 2.500 177.510 ;
        RECT 1.010 177.195 2.500 177.425 ;
        RECT 1.010 177.045 1.370 177.195 ;
        RECT 0.960 176.410 1.910 176.815 ;
        RECT 0.130 175.385 1.420 175.615 ;
        RECT 0.130 174.425 0.730 175.385 ;
        RECT 1.650 175.065 1.910 176.410 ;
        RECT 2.140 175.760 2.500 177.195 ;
        RECT 2.730 175.860 3.080 177.060 ;
        RECT 3.440 176.450 3.820 178.095 ;
        RECT 2.520 175.065 2.870 175.125 ;
        RECT 3.440 175.065 3.780 175.670 ;
        RECT 1.650 174.805 3.780 175.065 ;
        RECT 2.520 174.745 2.870 174.805 ;
        RECT 4.050 174.525 4.650 178.520 ;
        RECT 6.495 178.040 8.245 180.825 ;
        RECT 8.885 178.040 9.695 179.040 ;
        RECT 10.335 178.040 12.085 180.335 ;
        RECT 12.725 178.040 13.535 179.040 ;
        RECT 14.175 178.040 15.925 180.335 ;
        RECT 16.565 178.040 17.375 179.040 ;
        RECT 18.015 178.040 19.765 180.335 ;
        RECT 20.405 178.040 21.215 179.040 ;
        RECT 21.855 178.040 23.605 180.335 ;
        RECT 24.245 178.040 25.055 179.040 ;
        RECT 25.695 178.040 27.445 180.335 ;
        RECT 28.085 178.040 28.895 179.040 ;
        RECT 29.535 178.040 31.285 180.335 ;
        RECT 31.925 178.040 32.735 179.040 ;
        RECT 33.375 178.040 35.125 180.335 ;
        RECT 35.765 178.040 36.575 179.040 ;
        RECT 38.945 178.040 40.695 180.825 ;
        RECT 41.335 178.040 42.145 179.040 ;
        RECT 42.785 178.040 44.535 180.335 ;
        RECT 45.175 178.040 45.985 179.040 ;
        RECT 46.625 178.040 48.375 180.335 ;
        RECT 49.015 178.040 49.825 179.040 ;
        RECT 50.465 178.040 52.215 180.335 ;
        RECT 52.855 178.040 53.665 179.040 ;
        RECT 54.305 178.040 56.055 180.335 ;
        RECT 56.695 178.040 57.505 179.040 ;
        RECT 58.145 178.040 59.895 180.335 ;
        RECT 60.535 178.040 61.345 179.040 ;
        RECT 61.985 178.040 63.735 180.335 ;
        RECT 64.375 178.040 65.185 179.040 ;
        RECT 65.825 178.040 67.575 180.335 ;
        RECT 68.215 178.040 69.025 179.040 ;
        RECT 71.395 178.040 73.145 180.825 ;
        RECT 73.785 178.040 74.595 179.040 ;
        RECT 75.235 178.040 76.985 180.335 ;
        RECT 77.625 178.040 78.435 179.040 ;
        RECT 79.075 178.040 80.825 180.335 ;
        RECT 81.465 178.040 82.275 179.040 ;
        RECT 82.915 178.040 84.665 180.335 ;
        RECT 85.305 178.040 86.115 179.040 ;
        RECT 86.755 178.040 88.505 180.335 ;
        RECT 89.145 178.040 89.955 179.040 ;
        RECT 90.595 178.040 92.345 180.335 ;
        RECT 92.985 178.040 93.795 179.040 ;
        RECT 94.435 178.040 96.185 180.335 ;
        RECT 96.825 178.040 97.635 179.040 ;
        RECT 98.275 178.040 100.025 180.335 ;
        RECT 100.665 178.040 101.475 179.040 ;
        RECT 103.845 178.040 105.595 180.825 ;
        RECT 106.235 178.040 107.045 179.040 ;
        RECT 107.685 178.040 109.435 180.335 ;
        RECT 110.075 178.040 110.885 179.040 ;
        RECT 111.525 178.040 113.275 180.335 ;
        RECT 113.915 178.040 114.725 179.040 ;
        RECT 115.365 178.040 117.115 180.335 ;
        RECT 117.755 178.040 118.565 179.040 ;
        RECT 119.205 178.040 120.955 180.335 ;
        RECT 121.595 178.040 122.405 179.040 ;
        RECT 123.045 178.040 124.795 180.335 ;
        RECT 125.435 178.040 126.245 179.040 ;
        RECT 126.885 178.040 128.635 180.335 ;
        RECT 129.275 178.040 130.085 179.040 ;
        RECT 130.725 178.040 132.475 180.335 ;
        RECT 133.115 178.040 133.925 179.040 ;
        RECT 136.340 178.230 136.710 196.740 ;
        RECT 137.360 193.105 137.730 196.740 ;
        RECT 137.355 192.725 137.735 193.105 ;
        RECT 137.360 190.105 137.730 192.725 ;
        RECT 137.355 189.725 137.735 190.105 ;
        RECT 137.360 187.105 137.730 189.725 ;
        RECT 137.355 186.725 137.735 187.105 ;
        RECT 137.360 184.105 137.730 186.725 ;
        RECT 137.355 183.725 137.735 184.105 ;
        RECT 137.360 181.105 137.730 183.725 ;
        RECT 137.355 180.725 137.735 181.105 ;
        RECT 136.340 177.850 136.720 178.230 ;
        RECT 136.340 176.780 136.710 177.850 ;
        RECT 6.965 175.590 7.775 176.590 ;
        RECT 0.130 174.195 1.820 174.425 ;
        RECT 3.190 174.295 4.650 174.525 ;
        RECT 0.130 172.185 0.730 174.195 ;
        RECT 2.150 173.735 3.150 174.060 ;
        RECT 0.960 173.175 3.820 173.505 ;
        RECT 0.130 171.955 1.820 172.185 ;
        RECT 0.130 169.945 0.730 171.955 ;
        RECT 2.535 171.820 2.800 173.175 ;
        RECT 4.050 172.285 4.650 174.295 ;
        RECT 8.415 173.760 10.165 176.590 ;
        RECT 10.805 175.590 11.615 176.590 ;
        RECT 12.255 174.295 14.005 176.590 ;
        RECT 14.645 175.590 15.455 176.590 ;
        RECT 16.095 174.295 17.845 176.590 ;
        RECT 18.485 175.590 19.295 176.590 ;
        RECT 19.935 174.295 21.685 176.590 ;
        RECT 22.325 175.590 23.135 176.590 ;
        RECT 23.775 174.295 25.525 176.590 ;
        RECT 26.165 175.590 26.975 176.590 ;
        RECT 27.615 174.295 29.365 176.590 ;
        RECT 30.005 175.590 30.815 176.590 ;
        RECT 31.455 174.295 33.205 176.590 ;
        RECT 33.845 175.590 34.655 176.590 ;
        RECT 35.295 174.295 37.045 176.590 ;
        RECT 39.415 175.590 40.225 176.590 ;
        RECT 40.865 173.760 42.615 176.590 ;
        RECT 43.255 175.590 44.065 176.590 ;
        RECT 44.705 174.295 46.455 176.590 ;
        RECT 47.095 175.590 47.905 176.590 ;
        RECT 48.545 174.295 50.295 176.590 ;
        RECT 50.935 175.590 51.745 176.590 ;
        RECT 52.385 174.295 54.135 176.590 ;
        RECT 54.775 175.590 55.585 176.590 ;
        RECT 56.225 174.295 57.975 176.590 ;
        RECT 58.615 175.590 59.425 176.590 ;
        RECT 60.065 174.295 61.815 176.590 ;
        RECT 62.455 175.590 63.265 176.590 ;
        RECT 63.905 174.295 65.655 176.590 ;
        RECT 66.295 175.590 67.105 176.590 ;
        RECT 67.745 174.295 69.495 176.590 ;
        RECT 71.865 175.590 72.675 176.590 ;
        RECT 73.315 173.760 75.065 176.590 ;
        RECT 75.705 175.590 76.515 176.590 ;
        RECT 77.155 174.295 78.905 176.590 ;
        RECT 79.545 175.590 80.355 176.590 ;
        RECT 80.995 174.295 82.745 176.590 ;
        RECT 83.385 175.590 84.195 176.590 ;
        RECT 84.835 174.295 86.585 176.590 ;
        RECT 87.225 175.590 88.035 176.590 ;
        RECT 88.675 174.295 90.425 176.590 ;
        RECT 91.065 175.590 91.875 176.590 ;
        RECT 92.515 174.295 94.265 176.590 ;
        RECT 94.905 175.590 95.715 176.590 ;
        RECT 96.355 174.295 98.105 176.590 ;
        RECT 98.745 175.590 99.555 176.590 ;
        RECT 100.195 174.295 101.945 176.590 ;
        RECT 104.315 175.590 105.125 176.590 ;
        RECT 105.765 173.760 107.515 176.590 ;
        RECT 108.155 175.590 108.965 176.590 ;
        RECT 109.605 174.295 111.355 176.590 ;
        RECT 111.995 175.590 112.805 176.590 ;
        RECT 113.445 174.295 115.195 176.590 ;
        RECT 115.835 175.590 116.645 176.590 ;
        RECT 117.285 174.295 119.035 176.590 ;
        RECT 119.675 175.590 120.485 176.590 ;
        RECT 121.125 174.295 122.875 176.590 ;
        RECT 123.515 175.590 124.325 176.590 ;
        RECT 124.965 174.295 126.715 176.590 ;
        RECT 127.355 175.590 128.165 176.590 ;
        RECT 128.805 174.295 130.555 176.590 ;
        RECT 131.195 175.590 132.005 176.590 ;
        RECT 132.645 174.295 134.395 176.590 ;
        RECT 136.340 176.400 136.720 176.780 ;
        RECT 6.690 173.390 37.210 173.760 ;
        RECT 39.140 173.390 69.660 173.760 ;
        RECT 71.590 173.390 102.110 173.760 ;
        RECT 104.040 173.390 134.560 173.760 ;
        RECT 5.840 173.125 6.460 173.310 ;
        RECT 37.440 173.125 38.060 173.310 ;
        RECT 5.840 172.895 38.060 173.125 ;
        RECT 5.840 172.710 6.460 172.895 ;
        RECT 37.440 172.710 38.060 172.895 ;
        RECT 38.290 173.125 38.910 173.310 ;
        RECT 69.890 173.125 70.510 173.310 ;
        RECT 38.290 172.895 70.510 173.125 ;
        RECT 38.290 172.710 38.910 172.895 ;
        RECT 69.890 172.710 70.510 172.895 ;
        RECT 70.740 173.125 71.360 173.310 ;
        RECT 102.340 173.125 102.960 173.310 ;
        RECT 70.740 172.895 102.960 173.125 ;
        RECT 70.740 172.710 71.360 172.895 ;
        RECT 102.340 172.710 102.960 172.895 ;
        RECT 103.190 173.125 103.810 173.310 ;
        RECT 134.790 173.125 135.410 173.310 ;
        RECT 103.190 172.895 135.410 173.125 ;
        RECT 103.190 172.710 103.810 172.895 ;
        RECT 134.790 172.710 135.410 172.895 ;
        RECT 3.190 172.055 4.650 172.285 ;
        RECT 6.690 172.260 37.210 172.640 ;
        RECT 39.140 172.260 69.660 172.640 ;
        RECT 71.590 172.260 102.110 172.640 ;
        RECT 104.040 172.260 134.560 172.640 ;
        RECT 2.150 171.495 3.150 171.820 ;
        RECT 0.960 170.935 3.820 171.265 ;
        RECT 4.050 170.045 4.650 172.055 ;
        RECT 6.690 171.550 37.210 171.920 ;
        RECT 39.140 171.550 69.660 171.920 ;
        RECT 71.590 171.550 102.110 171.920 ;
        RECT 104.040 171.550 134.560 171.920 ;
        RECT 12.320 171.540 13.940 171.550 ;
        RECT 44.770 171.540 46.390 171.550 ;
        RECT 77.220 171.540 78.840 171.550 ;
        RECT 109.670 171.540 111.290 171.550 ;
        RECT 5.840 171.285 6.460 171.470 ;
        RECT 37.440 171.285 38.060 171.470 ;
        RECT 5.840 171.055 38.060 171.285 ;
        RECT 5.840 170.870 6.460 171.055 ;
        RECT 37.440 170.870 38.060 171.055 ;
        RECT 38.290 171.285 38.910 171.470 ;
        RECT 69.890 171.285 70.510 171.470 ;
        RECT 38.290 171.055 70.510 171.285 ;
        RECT 38.290 170.870 38.910 171.055 ;
        RECT 69.890 170.870 70.510 171.055 ;
        RECT 70.740 171.285 71.360 171.470 ;
        RECT 102.340 171.285 102.960 171.470 ;
        RECT 70.740 171.055 102.960 171.285 ;
        RECT 70.740 170.870 71.360 171.055 ;
        RECT 102.340 170.870 102.960 171.055 ;
        RECT 103.190 171.285 103.810 171.470 ;
        RECT 134.790 171.285 135.410 171.470 ;
        RECT 103.190 171.055 135.410 171.285 ;
        RECT 103.190 170.870 103.810 171.055 ;
        RECT 134.790 170.870 135.410 171.055 ;
        RECT 6.690 170.420 37.210 170.800 ;
        RECT 39.140 170.420 69.660 170.800 ;
        RECT 71.590 170.420 102.110 170.800 ;
        RECT 104.040 170.420 134.560 170.800 ;
        RECT 0.130 169.715 1.820 169.945 ;
        RECT 3.190 169.815 4.650 170.045 ;
        RECT 0.130 167.660 0.730 169.715 ;
        RECT 2.150 169.255 3.150 169.580 ;
        RECT 0.960 168.695 3.820 169.025 ;
        RECT 2.300 168.570 2.680 168.695 ;
        RECT 4.050 167.660 4.650 169.815 ;
        RECT 6.690 169.705 37.210 170.075 ;
        RECT 39.140 169.705 69.660 170.075 ;
        RECT 71.590 169.705 102.110 170.075 ;
        RECT 104.040 169.705 134.560 170.075 ;
        RECT 16.160 169.695 17.780 169.705 ;
        RECT 48.610 169.695 50.230 169.705 ;
        RECT 81.060 169.695 82.680 169.705 ;
        RECT 113.510 169.695 115.130 169.705 ;
        RECT 5.840 169.440 6.460 169.625 ;
        RECT 37.440 169.440 38.060 169.625 ;
        RECT 5.840 169.210 38.060 169.440 ;
        RECT 5.840 169.025 6.460 169.210 ;
        RECT 37.440 169.025 38.060 169.210 ;
        RECT 38.290 169.440 38.910 169.625 ;
        RECT 69.890 169.440 70.510 169.625 ;
        RECT 38.290 169.210 70.510 169.440 ;
        RECT 38.290 169.025 38.910 169.210 ;
        RECT 69.890 169.025 70.510 169.210 ;
        RECT 70.740 169.440 71.360 169.625 ;
        RECT 102.340 169.440 102.960 169.625 ;
        RECT 70.740 169.210 102.960 169.440 ;
        RECT 70.740 169.025 71.360 169.210 ;
        RECT 102.340 169.025 102.960 169.210 ;
        RECT 103.190 169.440 103.810 169.625 ;
        RECT 134.790 169.440 135.410 169.625 ;
        RECT 103.190 169.210 135.410 169.440 ;
        RECT 103.190 169.025 103.810 169.210 ;
        RECT 134.790 169.025 135.410 169.210 ;
        RECT 6.690 168.575 37.210 168.955 ;
        RECT 39.140 168.575 69.660 168.955 ;
        RECT 71.590 168.575 102.110 168.955 ;
        RECT 104.040 168.575 134.560 168.955 ;
        RECT 6.700 167.785 37.200 168.225 ;
        RECT 39.150 167.785 69.650 168.225 ;
        RECT 71.600 167.785 102.100 168.225 ;
        RECT 104.050 167.785 134.550 168.225 ;
        RECT 0.130 167.320 2.420 167.660 ;
        RECT 3.165 167.320 4.650 167.660 ;
        RECT 0.130 166.540 0.730 167.320 ;
        RECT 4.050 166.540 4.650 167.320 ;
        RECT 6.690 167.065 37.210 167.435 ;
        RECT 39.140 167.065 69.660 167.435 ;
        RECT 71.590 167.065 102.110 167.435 ;
        RECT 104.040 167.065 134.560 167.435 ;
        RECT 20.000 167.055 21.620 167.065 ;
        RECT 52.450 167.055 54.070 167.065 ;
        RECT 84.900 167.055 86.520 167.065 ;
        RECT 117.350 167.055 118.970 167.065 ;
        RECT 0.130 166.200 2.420 166.540 ;
        RECT 3.165 166.200 4.650 166.540 ;
        RECT 5.840 166.800 6.460 166.985 ;
        RECT 37.440 166.800 38.060 166.985 ;
        RECT 5.840 166.570 38.060 166.800 ;
        RECT 5.840 166.385 6.460 166.570 ;
        RECT 37.440 166.385 38.060 166.570 ;
        RECT 38.290 166.800 38.910 166.985 ;
        RECT 69.890 166.800 70.510 166.985 ;
        RECT 38.290 166.570 70.510 166.800 ;
        RECT 38.290 166.385 38.910 166.570 ;
        RECT 69.890 166.385 70.510 166.570 ;
        RECT 70.740 166.800 71.360 166.985 ;
        RECT 102.340 166.800 102.960 166.985 ;
        RECT 70.740 166.570 102.960 166.800 ;
        RECT 70.740 166.385 71.360 166.570 ;
        RECT 102.340 166.385 102.960 166.570 ;
        RECT 103.190 166.800 103.810 166.985 ;
        RECT 134.790 166.800 135.410 166.985 ;
        RECT 103.190 166.570 135.410 166.800 ;
        RECT 103.190 166.385 103.810 166.570 ;
        RECT 134.790 166.385 135.410 166.570 ;
        RECT 0.130 165.565 0.730 166.200 ;
        RECT 0.130 165.335 1.860 165.565 ;
        RECT 2.160 165.335 3.820 165.565 ;
        RECT 0.130 163.325 0.730 165.335 ;
        RECT 2.160 164.300 2.390 165.335 ;
        RECT 2.795 164.045 3.025 165.090 ;
        RECT 4.050 164.045 4.650 166.200 ;
        RECT 6.690 165.935 37.210 166.315 ;
        RECT 39.140 165.935 69.660 166.315 ;
        RECT 71.590 165.935 102.110 166.315 ;
        RECT 104.040 165.935 134.560 166.315 ;
        RECT 6.690 165.225 37.210 165.595 ;
        RECT 39.140 165.225 69.660 165.595 ;
        RECT 71.590 165.225 102.110 165.595 ;
        RECT 104.040 165.225 134.560 165.595 ;
        RECT 23.840 165.215 25.460 165.225 ;
        RECT 56.290 165.215 57.910 165.225 ;
        RECT 88.740 165.215 90.360 165.225 ;
        RECT 121.190 165.215 122.810 165.225 ;
        RECT 5.840 164.960 6.460 165.145 ;
        RECT 37.440 164.960 38.060 165.145 ;
        RECT 5.840 164.730 38.060 164.960 ;
        RECT 5.840 164.545 6.460 164.730 ;
        RECT 37.440 164.545 38.060 164.730 ;
        RECT 38.290 164.960 38.910 165.145 ;
        RECT 69.890 164.960 70.510 165.145 ;
        RECT 38.290 164.730 70.510 164.960 ;
        RECT 38.290 164.545 38.910 164.730 ;
        RECT 69.890 164.545 70.510 164.730 ;
        RECT 70.740 164.960 71.360 165.145 ;
        RECT 102.340 164.960 102.960 165.145 ;
        RECT 70.740 164.730 102.960 164.960 ;
        RECT 70.740 164.545 71.360 164.730 ;
        RECT 102.340 164.545 102.960 164.730 ;
        RECT 103.190 164.960 103.810 165.145 ;
        RECT 134.790 164.960 135.410 165.145 ;
        RECT 103.190 164.730 135.410 164.960 ;
        RECT 103.190 164.545 103.810 164.730 ;
        RECT 134.790 164.545 135.410 164.730 ;
        RECT 6.690 164.095 37.210 164.475 ;
        RECT 39.140 164.095 69.660 164.475 ;
        RECT 71.590 164.095 102.110 164.475 ;
        RECT 104.040 164.095 134.560 164.475 ;
        RECT 0.960 163.815 3.025 164.045 ;
        RECT 3.255 163.815 4.650 164.045 ;
        RECT 0.130 163.095 1.860 163.325 ;
        RECT 2.160 163.095 3.820 163.325 ;
        RECT 0.130 161.085 0.730 163.095 ;
        RECT 2.160 162.060 2.390 163.095 ;
        RECT 2.795 161.805 3.025 162.850 ;
        RECT 4.050 161.805 4.650 163.815 ;
        RECT 6.690 163.380 37.210 163.750 ;
        RECT 39.140 163.380 69.660 163.750 ;
        RECT 71.590 163.380 102.110 163.750 ;
        RECT 104.040 163.380 134.560 163.750 ;
        RECT 27.680 163.370 29.300 163.380 ;
        RECT 60.130 163.370 61.750 163.380 ;
        RECT 92.580 163.370 94.200 163.380 ;
        RECT 125.030 163.370 126.650 163.380 ;
        RECT 5.840 163.115 6.460 163.300 ;
        RECT 37.440 163.115 38.060 163.300 ;
        RECT 5.840 162.885 38.060 163.115 ;
        RECT 5.840 162.700 6.460 162.885 ;
        RECT 37.440 162.700 38.060 162.885 ;
        RECT 38.290 163.115 38.910 163.300 ;
        RECT 69.890 163.115 70.510 163.300 ;
        RECT 38.290 162.885 70.510 163.115 ;
        RECT 38.290 162.700 38.910 162.885 ;
        RECT 69.890 162.700 70.510 162.885 ;
        RECT 70.740 163.115 71.360 163.300 ;
        RECT 102.340 163.115 102.960 163.300 ;
        RECT 70.740 162.885 102.960 163.115 ;
        RECT 70.740 162.700 71.360 162.885 ;
        RECT 102.340 162.700 102.960 162.885 ;
        RECT 103.190 163.115 103.810 163.300 ;
        RECT 134.790 163.115 135.410 163.300 ;
        RECT 103.190 162.885 135.410 163.115 ;
        RECT 103.190 162.700 103.810 162.885 ;
        RECT 134.790 162.700 135.410 162.885 ;
        RECT 6.690 162.250 37.210 162.630 ;
        RECT 39.140 162.250 69.660 162.630 ;
        RECT 71.590 162.250 102.110 162.630 ;
        RECT 104.040 162.250 134.560 162.630 ;
        RECT 0.960 161.575 3.025 161.805 ;
        RECT 3.255 161.575 4.650 161.805 ;
        RECT 0.130 160.855 1.860 161.085 ;
        RECT 2.160 160.855 3.820 161.085 ;
        RECT 0.130 158.680 0.730 160.855 ;
        RECT 2.160 159.820 2.390 160.855 ;
        RECT 2.795 159.565 3.025 160.610 ;
        RECT 4.050 159.565 4.650 161.575 ;
        RECT 6.700 161.460 37.200 161.900 ;
        RECT 39.150 161.460 69.650 161.900 ;
        RECT 71.600 161.460 102.100 161.900 ;
        RECT 104.050 161.460 134.550 161.900 ;
        RECT 6.690 160.740 37.210 161.110 ;
        RECT 39.140 160.740 69.660 161.110 ;
        RECT 71.590 160.740 102.110 161.110 ;
        RECT 104.040 160.740 134.560 161.110 ;
        RECT 31.520 160.730 33.140 160.740 ;
        RECT 63.970 160.730 65.590 160.740 ;
        RECT 96.420 160.730 98.040 160.740 ;
        RECT 128.870 160.730 130.490 160.740 ;
        RECT 5.840 160.475 6.460 160.660 ;
        RECT 37.440 160.475 38.060 160.660 ;
        RECT 5.840 160.245 38.060 160.475 ;
        RECT 5.840 160.060 6.460 160.245 ;
        RECT 37.440 160.060 38.060 160.245 ;
        RECT 38.290 160.475 38.910 160.660 ;
        RECT 69.890 160.475 70.510 160.660 ;
        RECT 38.290 160.245 70.510 160.475 ;
        RECT 38.290 160.060 38.910 160.245 ;
        RECT 69.890 160.060 70.510 160.245 ;
        RECT 70.740 160.475 71.360 160.660 ;
        RECT 102.340 160.475 102.960 160.660 ;
        RECT 70.740 160.245 102.960 160.475 ;
        RECT 70.740 160.060 71.360 160.245 ;
        RECT 102.340 160.060 102.960 160.245 ;
        RECT 103.190 160.475 103.810 160.660 ;
        RECT 134.790 160.475 135.410 160.660 ;
        RECT 103.190 160.245 135.410 160.475 ;
        RECT 103.190 160.060 103.810 160.245 ;
        RECT 134.790 160.060 135.410 160.245 ;
        RECT 6.690 159.610 37.210 159.990 ;
        RECT 39.140 159.610 69.660 159.990 ;
        RECT 71.590 159.610 102.110 159.990 ;
        RECT 104.040 159.610 134.560 159.990 ;
        RECT 0.960 159.335 3.025 159.565 ;
        RECT 3.255 159.335 4.650 159.565 ;
        RECT 4.050 158.680 4.650 159.335 ;
        RECT 6.690 158.900 37.210 159.270 ;
        RECT 39.140 158.900 69.660 159.270 ;
        RECT 71.590 158.900 102.110 159.270 ;
        RECT 104.040 158.900 134.560 159.270 ;
        RECT 35.360 158.890 36.980 158.900 ;
        RECT 67.810 158.890 69.430 158.900 ;
        RECT 100.260 158.890 101.880 158.900 ;
        RECT 132.710 158.890 134.330 158.900 ;
        RECT 0.130 158.340 2.430 158.680 ;
        RECT 3.160 158.340 4.650 158.680 ;
        RECT 0.130 157.375 0.730 158.340 ;
        RECT 4.050 157.375 4.650 158.340 ;
        RECT 5.840 158.635 6.460 158.820 ;
        RECT 37.440 158.635 38.060 158.820 ;
        RECT 5.840 158.405 38.060 158.635 ;
        RECT 5.840 158.220 6.460 158.405 ;
        RECT 37.440 158.220 38.060 158.405 ;
        RECT 38.290 158.635 38.910 158.820 ;
        RECT 69.890 158.635 70.510 158.820 ;
        RECT 38.290 158.405 70.510 158.635 ;
        RECT 38.290 158.220 38.910 158.405 ;
        RECT 69.890 158.220 70.510 158.405 ;
        RECT 70.740 158.635 71.360 158.820 ;
        RECT 102.340 158.635 102.960 158.820 ;
        RECT 70.740 158.405 102.960 158.635 ;
        RECT 70.740 158.220 71.360 158.405 ;
        RECT 102.340 158.220 102.960 158.405 ;
        RECT 103.190 158.635 103.810 158.820 ;
        RECT 134.790 158.635 135.410 158.820 ;
        RECT 103.190 158.405 135.410 158.635 ;
        RECT 136.340 158.470 136.710 176.400 ;
        RECT 137.360 175.105 137.730 180.725 ;
        RECT 138.380 178.230 138.750 196.740 ;
        RECT 139.400 193.105 139.770 196.740 ;
        RECT 139.395 192.725 139.775 193.105 ;
        RECT 139.400 190.105 139.770 192.725 ;
        RECT 139.395 189.725 139.775 190.105 ;
        RECT 139.400 187.105 139.770 189.725 ;
        RECT 139.395 186.725 139.775 187.105 ;
        RECT 139.400 184.105 139.770 186.725 ;
        RECT 139.395 183.725 139.775 184.105 ;
        RECT 139.400 181.105 139.770 183.725 ;
        RECT 139.395 180.725 139.775 181.105 ;
        RECT 138.380 177.850 138.760 178.230 ;
        RECT 138.380 176.780 138.750 177.850 ;
        RECT 138.380 176.400 138.760 176.780 ;
        RECT 137.355 174.725 137.735 175.105 ;
        RECT 137.360 172.105 137.730 174.725 ;
        RECT 137.355 171.725 137.735 172.105 ;
        RECT 137.360 169.105 137.730 171.725 ;
        RECT 137.355 168.725 137.735 169.105 ;
        RECT 137.360 166.105 137.730 168.725 ;
        RECT 137.355 165.725 137.735 166.105 ;
        RECT 137.360 163.105 137.730 165.725 ;
        RECT 137.355 162.725 137.735 163.105 ;
        RECT 137.360 160.105 137.730 162.725 ;
        RECT 137.355 159.725 137.735 160.105 ;
        RECT 137.360 158.470 137.730 159.725 ;
        RECT 138.380 158.470 138.750 176.400 ;
        RECT 139.400 175.105 139.770 180.725 ;
        RECT 139.395 174.725 139.775 175.105 ;
        RECT 139.400 172.105 139.770 174.725 ;
        RECT 139.395 171.725 139.775 172.105 ;
        RECT 139.400 169.105 139.770 171.725 ;
        RECT 139.395 168.725 139.775 169.105 ;
        RECT 139.400 166.105 139.770 168.725 ;
        RECT 139.395 165.725 139.775 166.105 ;
        RECT 139.400 163.105 139.770 165.725 ;
        RECT 139.395 162.725 139.775 163.105 ;
        RECT 139.400 160.105 139.770 162.725 ;
        RECT 139.395 159.725 139.775 160.105 ;
        RECT 139.400 158.470 139.770 159.725 ;
        RECT 140.420 158.470 140.800 196.740 ;
        RECT 141.150 158.480 141.590 196.730 ;
        RECT 103.190 158.220 103.810 158.405 ;
        RECT 134.790 158.220 135.410 158.405 ;
        RECT 6.690 157.770 37.210 158.150 ;
        RECT 39.140 157.770 69.660 158.150 ;
        RECT 71.590 157.770 102.110 158.150 ;
        RECT 104.040 157.770 134.560 158.150 ;
        RECT 0.130 157.035 2.430 157.375 ;
        RECT 3.160 157.035 4.650 157.375 ;
        RECT 6.690 157.050 37.210 157.430 ;
        RECT 39.140 157.050 69.660 157.430 ;
        RECT 71.590 157.050 102.110 157.430 ;
        RECT 104.040 157.050 134.560 157.430 ;
        RECT 0.130 156.420 0.730 157.035 ;
        RECT 0.130 156.190 1.860 156.420 ;
        RECT 2.160 156.190 3.820 156.420 ;
        RECT 0.130 154.180 0.730 156.190 ;
        RECT 2.160 155.155 2.390 156.190 ;
        RECT 2.795 154.900 3.025 155.945 ;
        RECT 4.050 154.900 4.650 157.035 ;
        RECT 5.840 156.795 6.460 156.980 ;
        RECT 37.440 156.795 38.060 156.980 ;
        RECT 5.840 156.565 38.060 156.795 ;
        RECT 5.840 156.380 6.460 156.565 ;
        RECT 37.440 156.380 38.060 156.565 ;
        RECT 38.290 156.795 38.910 156.980 ;
        RECT 69.890 156.795 70.510 156.980 ;
        RECT 38.290 156.565 70.510 156.795 ;
        RECT 38.290 156.380 38.910 156.565 ;
        RECT 69.890 156.380 70.510 156.565 ;
        RECT 70.740 156.795 71.360 156.980 ;
        RECT 102.340 156.795 102.960 156.980 ;
        RECT 70.740 156.565 102.960 156.795 ;
        RECT 70.740 156.380 71.360 156.565 ;
        RECT 102.340 156.380 102.960 156.565 ;
        RECT 103.190 156.795 103.810 156.980 ;
        RECT 134.790 156.795 135.410 156.980 ;
        RECT 103.190 156.565 135.410 156.795 ;
        RECT 103.190 156.380 103.810 156.565 ;
        RECT 134.790 156.380 135.410 156.565 ;
        RECT 33.440 156.300 35.060 156.310 ;
        RECT 65.890 156.300 67.510 156.310 ;
        RECT 98.340 156.300 99.960 156.310 ;
        RECT 130.790 156.300 132.410 156.310 ;
        RECT 6.690 155.930 37.210 156.300 ;
        RECT 39.140 155.930 69.660 156.300 ;
        RECT 71.590 155.930 102.110 156.300 ;
        RECT 104.040 155.930 134.560 156.300 ;
        RECT 6.690 155.210 37.210 155.590 ;
        RECT 39.140 155.210 69.660 155.590 ;
        RECT 71.590 155.210 102.110 155.590 ;
        RECT 104.040 155.210 134.560 155.590 ;
        RECT 0.960 154.670 3.025 154.900 ;
        RECT 3.255 154.670 4.650 154.900 ;
        RECT 0.130 153.950 1.860 154.180 ;
        RECT 2.160 153.950 3.820 154.180 ;
        RECT 0.130 151.940 0.730 153.950 ;
        RECT 2.160 152.915 2.390 153.950 ;
        RECT 2.795 152.660 3.025 153.705 ;
        RECT 4.050 152.660 4.650 154.670 ;
        RECT 5.840 154.955 6.460 155.140 ;
        RECT 37.440 154.955 38.060 155.140 ;
        RECT 5.840 154.725 38.060 154.955 ;
        RECT 5.840 154.540 6.460 154.725 ;
        RECT 37.440 154.540 38.060 154.725 ;
        RECT 38.290 154.955 38.910 155.140 ;
        RECT 69.890 154.955 70.510 155.140 ;
        RECT 38.290 154.725 70.510 154.955 ;
        RECT 38.290 154.540 38.910 154.725 ;
        RECT 69.890 154.540 70.510 154.725 ;
        RECT 70.740 154.955 71.360 155.140 ;
        RECT 102.340 154.955 102.960 155.140 ;
        RECT 70.740 154.725 102.960 154.955 ;
        RECT 70.740 154.540 71.360 154.725 ;
        RECT 102.340 154.540 102.960 154.725 ;
        RECT 103.190 154.955 103.810 155.140 ;
        RECT 134.790 154.955 135.410 155.140 ;
        RECT 103.190 154.725 135.410 154.955 ;
        RECT 103.190 154.540 103.810 154.725 ;
        RECT 134.790 154.540 135.410 154.725 ;
        RECT 29.600 154.460 31.220 154.470 ;
        RECT 62.050 154.460 63.670 154.470 ;
        RECT 94.500 154.460 96.120 154.470 ;
        RECT 126.950 154.460 128.570 154.470 ;
        RECT 6.690 154.090 37.210 154.460 ;
        RECT 39.140 154.090 69.660 154.460 ;
        RECT 71.590 154.090 102.110 154.460 ;
        RECT 104.040 154.090 134.560 154.460 ;
        RECT 6.700 153.295 37.200 153.735 ;
        RECT 39.150 153.295 69.650 153.735 ;
        RECT 71.600 153.295 102.100 153.735 ;
        RECT 104.050 153.295 134.550 153.735 ;
        RECT 0.960 152.430 3.025 152.660 ;
        RECT 3.255 152.430 4.650 152.660 ;
        RECT 6.690 152.565 37.210 152.945 ;
        RECT 39.140 152.565 69.660 152.945 ;
        RECT 71.590 152.565 102.110 152.945 ;
        RECT 104.040 152.565 134.560 152.945 ;
        RECT 0.130 151.710 1.860 151.940 ;
        RECT 2.160 151.710 3.820 151.940 ;
        RECT 0.130 149.700 0.730 151.710 ;
        RECT 2.160 150.675 2.390 151.710 ;
        RECT 2.795 150.420 3.025 151.465 ;
        RECT 4.050 150.420 4.650 152.430 ;
        RECT 5.840 152.310 6.460 152.495 ;
        RECT 37.440 152.310 38.060 152.495 ;
        RECT 5.840 152.080 38.060 152.310 ;
        RECT 5.840 151.895 6.460 152.080 ;
        RECT 37.440 151.895 38.060 152.080 ;
        RECT 38.290 152.310 38.910 152.495 ;
        RECT 69.890 152.310 70.510 152.495 ;
        RECT 38.290 152.080 70.510 152.310 ;
        RECT 38.290 151.895 38.910 152.080 ;
        RECT 69.890 151.895 70.510 152.080 ;
        RECT 70.740 152.310 71.360 152.495 ;
        RECT 102.340 152.310 102.960 152.495 ;
        RECT 70.740 152.080 102.960 152.310 ;
        RECT 70.740 151.895 71.360 152.080 ;
        RECT 102.340 151.895 102.960 152.080 ;
        RECT 103.190 152.310 103.810 152.495 ;
        RECT 134.790 152.310 135.410 152.495 ;
        RECT 103.190 152.080 135.410 152.310 ;
        RECT 103.190 151.895 103.810 152.080 ;
        RECT 134.790 151.895 135.410 152.080 ;
        RECT 25.760 151.815 27.380 151.825 ;
        RECT 58.210 151.815 59.830 151.825 ;
        RECT 90.660 151.815 92.280 151.825 ;
        RECT 123.110 151.815 124.730 151.825 ;
        RECT 6.690 151.445 37.210 151.815 ;
        RECT 39.140 151.445 69.660 151.815 ;
        RECT 71.590 151.445 102.110 151.815 ;
        RECT 104.040 151.445 134.560 151.815 ;
        RECT 6.690 150.725 37.210 151.105 ;
        RECT 39.140 150.725 69.660 151.105 ;
        RECT 71.590 150.725 102.110 151.105 ;
        RECT 104.040 150.725 134.560 151.105 ;
        RECT 0.960 150.190 3.025 150.420 ;
        RECT 3.255 150.190 4.650 150.420 ;
        RECT 0.130 149.470 1.860 149.700 ;
        RECT 2.160 149.470 3.820 149.700 ;
        RECT 0.130 147.460 0.730 149.470 ;
        RECT 2.160 148.435 2.390 149.470 ;
        RECT 2.795 148.180 3.025 149.225 ;
        RECT 4.050 148.180 4.650 150.190 ;
        RECT 5.840 150.470 6.460 150.655 ;
        RECT 37.440 150.470 38.060 150.655 ;
        RECT 5.840 150.240 38.060 150.470 ;
        RECT 5.840 150.055 6.460 150.240 ;
        RECT 37.440 150.055 38.060 150.240 ;
        RECT 38.290 150.470 38.910 150.655 ;
        RECT 69.890 150.470 70.510 150.655 ;
        RECT 38.290 150.240 70.510 150.470 ;
        RECT 38.290 150.055 38.910 150.240 ;
        RECT 69.890 150.055 70.510 150.240 ;
        RECT 70.740 150.470 71.360 150.655 ;
        RECT 102.340 150.470 102.960 150.655 ;
        RECT 70.740 150.240 102.960 150.470 ;
        RECT 70.740 150.055 71.360 150.240 ;
        RECT 102.340 150.055 102.960 150.240 ;
        RECT 103.190 150.470 103.810 150.655 ;
        RECT 134.790 150.470 135.410 150.655 ;
        RECT 103.190 150.240 135.410 150.470 ;
        RECT 103.190 150.055 103.810 150.240 ;
        RECT 134.790 150.055 135.410 150.240 ;
        RECT 21.920 149.975 23.540 149.985 ;
        RECT 54.370 149.975 55.990 149.985 ;
        RECT 86.820 149.975 88.440 149.985 ;
        RECT 119.270 149.975 120.890 149.985 ;
        RECT 6.690 149.605 37.210 149.975 ;
        RECT 39.140 149.605 69.660 149.975 ;
        RECT 71.590 149.605 102.110 149.975 ;
        RECT 104.040 149.605 134.560 149.975 ;
        RECT 6.690 148.885 37.210 149.265 ;
        RECT 39.140 148.885 69.660 149.265 ;
        RECT 71.590 148.885 102.110 149.265 ;
        RECT 104.040 148.885 134.560 149.265 ;
        RECT 5.840 148.630 6.460 148.815 ;
        RECT 37.440 148.630 38.060 148.815 ;
        RECT 5.840 148.400 38.060 148.630 ;
        RECT 5.840 148.215 6.460 148.400 ;
        RECT 37.440 148.215 38.060 148.400 ;
        RECT 38.290 148.630 38.910 148.815 ;
        RECT 69.890 148.630 70.510 148.815 ;
        RECT 38.290 148.400 70.510 148.630 ;
        RECT 38.290 148.215 38.910 148.400 ;
        RECT 69.890 148.215 70.510 148.400 ;
        RECT 70.740 148.630 71.360 148.815 ;
        RECT 102.340 148.630 102.960 148.815 ;
        RECT 70.740 148.400 102.960 148.630 ;
        RECT 70.740 148.215 71.360 148.400 ;
        RECT 102.340 148.215 102.960 148.400 ;
        RECT 103.190 148.630 103.810 148.815 ;
        RECT 134.790 148.630 135.410 148.815 ;
        RECT 103.190 148.400 135.410 148.630 ;
        RECT 103.190 148.215 103.810 148.400 ;
        RECT 134.790 148.215 135.410 148.400 ;
        RECT 0.960 147.950 3.025 148.180 ;
        RECT 3.255 147.950 4.650 148.180 ;
        RECT 18.080 148.135 19.700 148.145 ;
        RECT 50.530 148.135 52.150 148.145 ;
        RECT 82.980 148.135 84.600 148.145 ;
        RECT 115.430 148.135 117.050 148.145 ;
        RECT 0.130 147.230 1.860 147.460 ;
        RECT 2.160 147.230 3.820 147.460 ;
        RECT 0.130 145.075 0.730 147.230 ;
        RECT 2.160 146.195 2.390 147.230 ;
        RECT 2.795 145.940 3.025 146.985 ;
        RECT 4.050 145.940 4.650 147.950 ;
        RECT 6.690 147.765 37.210 148.135 ;
        RECT 39.140 147.765 69.660 148.135 ;
        RECT 71.590 147.765 102.110 148.135 ;
        RECT 104.040 147.765 134.560 148.135 ;
        RECT 6.700 146.970 37.200 147.410 ;
        RECT 39.150 146.970 69.650 147.410 ;
        RECT 71.600 146.970 102.100 147.410 ;
        RECT 104.050 146.970 134.550 147.410 ;
        RECT 6.690 146.240 37.210 146.620 ;
        RECT 39.140 146.240 69.660 146.620 ;
        RECT 71.590 146.240 102.110 146.620 ;
        RECT 104.040 146.240 134.560 146.620 ;
        RECT 0.960 145.710 3.025 145.940 ;
        RECT 3.255 145.710 4.650 145.940 ;
        RECT 4.050 145.075 4.650 145.710 ;
        RECT 5.840 145.985 6.460 146.170 ;
        RECT 37.440 145.985 38.060 146.170 ;
        RECT 5.840 145.755 38.060 145.985 ;
        RECT 5.840 145.570 6.460 145.755 ;
        RECT 37.440 145.570 38.060 145.755 ;
        RECT 38.290 145.985 38.910 146.170 ;
        RECT 69.890 145.985 70.510 146.170 ;
        RECT 38.290 145.755 70.510 145.985 ;
        RECT 38.290 145.570 38.910 145.755 ;
        RECT 69.890 145.570 70.510 145.755 ;
        RECT 70.740 145.985 71.360 146.170 ;
        RECT 102.340 145.985 102.960 146.170 ;
        RECT 70.740 145.755 102.960 145.985 ;
        RECT 70.740 145.570 71.360 145.755 ;
        RECT 102.340 145.570 102.960 145.755 ;
        RECT 103.190 145.985 103.810 146.170 ;
        RECT 134.790 145.985 135.410 146.170 ;
        RECT 103.190 145.755 135.410 145.985 ;
        RECT 103.190 145.570 103.810 145.755 ;
        RECT 134.790 145.570 135.410 145.755 ;
        RECT 14.240 145.490 15.860 145.500 ;
        RECT 46.690 145.490 48.310 145.500 ;
        RECT 79.140 145.490 80.760 145.500 ;
        RECT 111.590 145.490 113.210 145.500 ;
        RECT 6.690 145.120 37.210 145.490 ;
        RECT 39.140 145.120 69.660 145.490 ;
        RECT 71.590 145.120 102.110 145.490 ;
        RECT 104.040 145.120 134.560 145.490 ;
        RECT 0.130 144.735 2.420 145.075 ;
        RECT 3.165 144.735 4.650 145.075 ;
        RECT 0.130 144.100 0.730 144.735 ;
        RECT 0.130 143.870 1.860 144.100 ;
        RECT 2.160 143.870 3.820 144.100 ;
        RECT 0.130 141.860 0.730 143.870 ;
        RECT 2.160 142.835 2.390 143.870 ;
        RECT 2.795 142.580 3.025 143.625 ;
        RECT 4.050 142.580 4.650 144.735 ;
        RECT 6.690 144.400 37.210 144.780 ;
        RECT 39.140 144.400 69.660 144.780 ;
        RECT 71.590 144.400 102.110 144.780 ;
        RECT 104.040 144.400 134.560 144.780 ;
        RECT 5.840 144.145 6.460 144.330 ;
        RECT 37.440 144.145 38.060 144.330 ;
        RECT 5.840 143.915 38.060 144.145 ;
        RECT 5.840 143.730 6.460 143.915 ;
        RECT 37.440 143.730 38.060 143.915 ;
        RECT 38.290 144.145 38.910 144.330 ;
        RECT 69.890 144.145 70.510 144.330 ;
        RECT 38.290 143.915 70.510 144.145 ;
        RECT 38.290 143.730 38.910 143.915 ;
        RECT 69.890 143.730 70.510 143.915 ;
        RECT 70.740 144.145 71.360 144.330 ;
        RECT 102.340 144.145 102.960 144.330 ;
        RECT 70.740 143.915 102.960 144.145 ;
        RECT 70.740 143.730 71.360 143.915 ;
        RECT 102.340 143.730 102.960 143.915 ;
        RECT 103.190 144.145 103.810 144.330 ;
        RECT 134.790 144.145 135.410 144.330 ;
        RECT 103.190 143.915 135.410 144.145 ;
        RECT 103.190 143.730 103.810 143.915 ;
        RECT 134.790 143.730 135.410 143.915 ;
        RECT 10.400 143.650 12.020 143.660 ;
        RECT 42.850 143.650 44.470 143.660 ;
        RECT 75.300 143.650 76.920 143.660 ;
        RECT 107.750 143.650 109.370 143.660 ;
        RECT 6.690 143.280 37.210 143.650 ;
        RECT 39.140 143.280 69.660 143.650 ;
        RECT 71.590 143.280 102.110 143.650 ;
        RECT 104.040 143.280 134.560 143.650 ;
        RECT 0.960 142.350 3.025 142.580 ;
        RECT 3.255 142.350 4.650 142.580 ;
        RECT 6.690 142.560 37.210 142.940 ;
        RECT 39.140 142.560 69.660 142.940 ;
        RECT 71.590 142.560 102.110 142.940 ;
        RECT 104.040 142.560 134.560 142.940 ;
        RECT 0.130 141.630 1.860 141.860 ;
        RECT 2.160 141.630 3.820 141.860 ;
        RECT 0.130 139.475 0.730 141.630 ;
        RECT 2.160 140.595 2.390 141.630 ;
        RECT 2.795 140.340 3.025 141.385 ;
        RECT 4.050 140.340 4.650 142.350 ;
        RECT 5.840 142.305 6.460 142.490 ;
        RECT 37.440 142.305 38.060 142.490 ;
        RECT 5.840 142.075 38.060 142.305 ;
        RECT 5.840 141.890 6.460 142.075 ;
        RECT 37.440 141.890 38.060 142.075 ;
        RECT 38.290 142.305 38.910 142.490 ;
        RECT 69.890 142.305 70.510 142.490 ;
        RECT 38.290 142.075 70.510 142.305 ;
        RECT 38.290 141.890 38.910 142.075 ;
        RECT 69.890 141.890 70.510 142.075 ;
        RECT 70.740 142.305 71.360 142.490 ;
        RECT 102.340 142.305 102.960 142.490 ;
        RECT 70.740 142.075 102.960 142.305 ;
        RECT 70.740 141.890 71.360 142.075 ;
        RECT 102.340 141.890 102.960 142.075 ;
        RECT 103.190 142.305 103.810 142.490 ;
        RECT 134.790 142.305 135.410 142.490 ;
        RECT 103.190 142.075 135.410 142.305 ;
        RECT 103.190 141.890 103.810 142.075 ;
        RECT 134.790 141.890 135.410 142.075 ;
        RECT 6.690 141.440 37.210 141.810 ;
        RECT 39.140 141.440 69.660 141.810 ;
        RECT 71.590 141.440 102.110 141.810 ;
        RECT 104.040 141.440 134.560 141.810 ;
        RECT 0.960 140.110 3.025 140.340 ;
        RECT 3.255 140.110 4.650 140.340 ;
        RECT 4.050 139.475 4.650 140.110 ;
        RECT 0.130 139.135 2.420 139.475 ;
        RECT 3.165 139.135 4.650 139.475 ;
        RECT 0.130 138.500 0.730 139.135 ;
        RECT 0.130 138.270 1.710 138.500 ;
        RECT 0.130 136.230 0.730 138.270 ;
        RECT 2.140 138.040 2.500 138.125 ;
        RECT 1.010 137.810 2.500 138.040 ;
        RECT 1.010 137.660 1.370 137.810 ;
        RECT 0.960 137.025 1.910 137.430 ;
        RECT 0.130 136.000 1.420 136.230 ;
        RECT 0.130 135.040 0.730 136.000 ;
        RECT 1.650 135.680 1.910 137.025 ;
        RECT 2.140 136.375 2.500 137.810 ;
        RECT 2.730 136.475 3.080 137.675 ;
        RECT 3.440 137.065 3.820 138.710 ;
        RECT 2.520 135.680 2.870 135.740 ;
        RECT 3.440 135.680 3.780 136.285 ;
        RECT 1.650 135.420 3.780 135.680 ;
        RECT 2.520 135.360 2.870 135.420 ;
        RECT 4.050 135.140 4.650 139.135 ;
        RECT 6.495 138.655 8.245 141.440 ;
        RECT 8.885 138.655 9.695 139.655 ;
        RECT 10.335 138.655 12.085 140.950 ;
        RECT 12.725 138.655 13.535 139.655 ;
        RECT 14.175 138.655 15.925 140.950 ;
        RECT 16.565 138.655 17.375 139.655 ;
        RECT 18.015 138.655 19.765 140.950 ;
        RECT 20.405 138.655 21.215 139.655 ;
        RECT 21.855 138.655 23.605 140.950 ;
        RECT 24.245 138.655 25.055 139.655 ;
        RECT 25.695 138.655 27.445 140.950 ;
        RECT 28.085 138.655 28.895 139.655 ;
        RECT 29.535 138.655 31.285 140.950 ;
        RECT 31.925 138.655 32.735 139.655 ;
        RECT 33.375 138.655 35.125 140.950 ;
        RECT 35.765 138.655 36.575 139.655 ;
        RECT 38.945 138.655 40.695 141.440 ;
        RECT 41.335 138.655 42.145 139.655 ;
        RECT 42.785 138.655 44.535 140.950 ;
        RECT 45.175 138.655 45.985 139.655 ;
        RECT 46.625 138.655 48.375 140.950 ;
        RECT 49.015 138.655 49.825 139.655 ;
        RECT 50.465 138.655 52.215 140.950 ;
        RECT 52.855 138.655 53.665 139.655 ;
        RECT 54.305 138.655 56.055 140.950 ;
        RECT 56.695 138.655 57.505 139.655 ;
        RECT 58.145 138.655 59.895 140.950 ;
        RECT 60.535 138.655 61.345 139.655 ;
        RECT 61.985 138.655 63.735 140.950 ;
        RECT 64.375 138.655 65.185 139.655 ;
        RECT 65.825 138.655 67.575 140.950 ;
        RECT 68.215 138.655 69.025 139.655 ;
        RECT 71.395 138.655 73.145 141.440 ;
        RECT 73.785 138.655 74.595 139.655 ;
        RECT 75.235 138.655 76.985 140.950 ;
        RECT 77.625 138.655 78.435 139.655 ;
        RECT 79.075 138.655 80.825 140.950 ;
        RECT 81.465 138.655 82.275 139.655 ;
        RECT 82.915 138.655 84.665 140.950 ;
        RECT 85.305 138.655 86.115 139.655 ;
        RECT 86.755 138.655 88.505 140.950 ;
        RECT 89.145 138.655 89.955 139.655 ;
        RECT 90.595 138.655 92.345 140.950 ;
        RECT 92.985 138.655 93.795 139.655 ;
        RECT 94.435 138.655 96.185 140.950 ;
        RECT 96.825 138.655 97.635 139.655 ;
        RECT 98.275 138.655 100.025 140.950 ;
        RECT 100.665 138.655 101.475 139.655 ;
        RECT 103.845 138.655 105.595 141.440 ;
        RECT 106.235 138.655 107.045 139.655 ;
        RECT 107.685 138.655 109.435 140.950 ;
        RECT 110.075 138.655 110.885 139.655 ;
        RECT 111.525 138.655 113.275 140.950 ;
        RECT 113.915 138.655 114.725 139.655 ;
        RECT 115.365 138.655 117.115 140.950 ;
        RECT 117.755 138.655 118.565 139.655 ;
        RECT 119.205 138.655 120.955 140.950 ;
        RECT 121.595 138.655 122.405 139.655 ;
        RECT 123.045 138.655 124.795 140.950 ;
        RECT 125.435 138.655 126.245 139.655 ;
        RECT 126.885 138.655 128.635 140.950 ;
        RECT 129.275 138.655 130.085 139.655 ;
        RECT 130.725 138.655 132.475 140.950 ;
        RECT 133.115 138.655 133.925 139.655 ;
        RECT 136.340 138.845 136.710 157.355 ;
        RECT 137.360 153.720 137.730 157.355 ;
        RECT 137.355 153.340 137.735 153.720 ;
        RECT 137.360 150.720 137.730 153.340 ;
        RECT 137.355 150.340 137.735 150.720 ;
        RECT 137.360 147.720 137.730 150.340 ;
        RECT 137.355 147.340 137.735 147.720 ;
        RECT 137.360 144.720 137.730 147.340 ;
        RECT 137.355 144.340 137.735 144.720 ;
        RECT 137.360 141.720 137.730 144.340 ;
        RECT 137.355 141.340 137.735 141.720 ;
        RECT 136.340 138.465 136.720 138.845 ;
        RECT 136.340 137.395 136.710 138.465 ;
        RECT 6.965 136.205 7.775 137.205 ;
        RECT 0.130 134.810 1.820 135.040 ;
        RECT 3.190 134.910 4.650 135.140 ;
        RECT 0.130 132.800 0.730 134.810 ;
        RECT 2.150 134.350 3.150 134.675 ;
        RECT 0.960 133.790 3.820 134.120 ;
        RECT 0.130 132.570 1.820 132.800 ;
        RECT 0.130 130.560 0.730 132.570 ;
        RECT 2.535 132.435 2.800 133.790 ;
        RECT 4.050 132.900 4.650 134.910 ;
        RECT 8.415 134.375 10.165 137.205 ;
        RECT 10.805 136.205 11.615 137.205 ;
        RECT 12.255 134.910 14.005 137.205 ;
        RECT 14.645 136.205 15.455 137.205 ;
        RECT 16.095 134.910 17.845 137.205 ;
        RECT 18.485 136.205 19.295 137.205 ;
        RECT 19.935 134.910 21.685 137.205 ;
        RECT 22.325 136.205 23.135 137.205 ;
        RECT 23.775 134.910 25.525 137.205 ;
        RECT 26.165 136.205 26.975 137.205 ;
        RECT 27.615 134.910 29.365 137.205 ;
        RECT 30.005 136.205 30.815 137.205 ;
        RECT 31.455 134.910 33.205 137.205 ;
        RECT 33.845 136.205 34.655 137.205 ;
        RECT 35.295 134.910 37.045 137.205 ;
        RECT 39.415 136.205 40.225 137.205 ;
        RECT 40.865 134.375 42.615 137.205 ;
        RECT 43.255 136.205 44.065 137.205 ;
        RECT 44.705 134.910 46.455 137.205 ;
        RECT 47.095 136.205 47.905 137.205 ;
        RECT 48.545 134.910 50.295 137.205 ;
        RECT 50.935 136.205 51.745 137.205 ;
        RECT 52.385 134.910 54.135 137.205 ;
        RECT 54.775 136.205 55.585 137.205 ;
        RECT 56.225 134.910 57.975 137.205 ;
        RECT 58.615 136.205 59.425 137.205 ;
        RECT 60.065 134.910 61.815 137.205 ;
        RECT 62.455 136.205 63.265 137.205 ;
        RECT 63.905 134.910 65.655 137.205 ;
        RECT 66.295 136.205 67.105 137.205 ;
        RECT 67.745 134.910 69.495 137.205 ;
        RECT 71.865 136.205 72.675 137.205 ;
        RECT 73.315 134.375 75.065 137.205 ;
        RECT 75.705 136.205 76.515 137.205 ;
        RECT 77.155 134.910 78.905 137.205 ;
        RECT 79.545 136.205 80.355 137.205 ;
        RECT 80.995 134.910 82.745 137.205 ;
        RECT 83.385 136.205 84.195 137.205 ;
        RECT 84.835 134.910 86.585 137.205 ;
        RECT 87.225 136.205 88.035 137.205 ;
        RECT 88.675 134.910 90.425 137.205 ;
        RECT 91.065 136.205 91.875 137.205 ;
        RECT 92.515 134.910 94.265 137.205 ;
        RECT 94.905 136.205 95.715 137.205 ;
        RECT 96.355 134.910 98.105 137.205 ;
        RECT 98.745 136.205 99.555 137.205 ;
        RECT 100.195 134.910 101.945 137.205 ;
        RECT 104.315 136.205 105.125 137.205 ;
        RECT 105.765 134.375 107.515 137.205 ;
        RECT 108.155 136.205 108.965 137.205 ;
        RECT 109.605 134.910 111.355 137.205 ;
        RECT 111.995 136.205 112.805 137.205 ;
        RECT 113.445 134.910 115.195 137.205 ;
        RECT 115.835 136.205 116.645 137.205 ;
        RECT 117.285 134.910 119.035 137.205 ;
        RECT 119.675 136.205 120.485 137.205 ;
        RECT 121.125 134.910 122.875 137.205 ;
        RECT 123.515 136.205 124.325 137.205 ;
        RECT 124.965 134.910 126.715 137.205 ;
        RECT 127.355 136.205 128.165 137.205 ;
        RECT 128.805 134.910 130.555 137.205 ;
        RECT 131.195 136.205 132.005 137.205 ;
        RECT 132.645 134.910 134.395 137.205 ;
        RECT 136.340 137.015 136.720 137.395 ;
        RECT 6.690 134.005 37.210 134.375 ;
        RECT 39.140 134.005 69.660 134.375 ;
        RECT 71.590 134.005 102.110 134.375 ;
        RECT 104.040 134.005 134.560 134.375 ;
        RECT 5.840 133.740 6.460 133.925 ;
        RECT 37.440 133.740 38.060 133.925 ;
        RECT 5.840 133.510 38.060 133.740 ;
        RECT 5.840 133.325 6.460 133.510 ;
        RECT 37.440 133.325 38.060 133.510 ;
        RECT 38.290 133.740 38.910 133.925 ;
        RECT 69.890 133.740 70.510 133.925 ;
        RECT 38.290 133.510 70.510 133.740 ;
        RECT 38.290 133.325 38.910 133.510 ;
        RECT 69.890 133.325 70.510 133.510 ;
        RECT 70.740 133.740 71.360 133.925 ;
        RECT 102.340 133.740 102.960 133.925 ;
        RECT 70.740 133.510 102.960 133.740 ;
        RECT 70.740 133.325 71.360 133.510 ;
        RECT 102.340 133.325 102.960 133.510 ;
        RECT 103.190 133.740 103.810 133.925 ;
        RECT 134.790 133.740 135.410 133.925 ;
        RECT 103.190 133.510 135.410 133.740 ;
        RECT 103.190 133.325 103.810 133.510 ;
        RECT 134.790 133.325 135.410 133.510 ;
        RECT 3.190 132.670 4.650 132.900 ;
        RECT 6.690 132.875 37.210 133.255 ;
        RECT 39.140 132.875 69.660 133.255 ;
        RECT 71.590 132.875 102.110 133.255 ;
        RECT 104.040 132.875 134.560 133.255 ;
        RECT 2.150 132.110 3.150 132.435 ;
        RECT 0.960 131.550 3.820 131.880 ;
        RECT 4.050 130.660 4.650 132.670 ;
        RECT 6.690 132.165 37.210 132.535 ;
        RECT 39.140 132.165 69.660 132.535 ;
        RECT 71.590 132.165 102.110 132.535 ;
        RECT 104.040 132.165 134.560 132.535 ;
        RECT 12.320 132.155 13.940 132.165 ;
        RECT 44.770 132.155 46.390 132.165 ;
        RECT 77.220 132.155 78.840 132.165 ;
        RECT 109.670 132.155 111.290 132.165 ;
        RECT 5.840 131.900 6.460 132.085 ;
        RECT 37.440 131.900 38.060 132.085 ;
        RECT 5.840 131.670 38.060 131.900 ;
        RECT 5.840 131.485 6.460 131.670 ;
        RECT 37.440 131.485 38.060 131.670 ;
        RECT 38.290 131.900 38.910 132.085 ;
        RECT 69.890 131.900 70.510 132.085 ;
        RECT 38.290 131.670 70.510 131.900 ;
        RECT 38.290 131.485 38.910 131.670 ;
        RECT 69.890 131.485 70.510 131.670 ;
        RECT 70.740 131.900 71.360 132.085 ;
        RECT 102.340 131.900 102.960 132.085 ;
        RECT 70.740 131.670 102.960 131.900 ;
        RECT 70.740 131.485 71.360 131.670 ;
        RECT 102.340 131.485 102.960 131.670 ;
        RECT 103.190 131.900 103.810 132.085 ;
        RECT 134.790 131.900 135.410 132.085 ;
        RECT 103.190 131.670 135.410 131.900 ;
        RECT 103.190 131.485 103.810 131.670 ;
        RECT 134.790 131.485 135.410 131.670 ;
        RECT 6.690 131.035 37.210 131.415 ;
        RECT 39.140 131.035 69.660 131.415 ;
        RECT 71.590 131.035 102.110 131.415 ;
        RECT 104.040 131.035 134.560 131.415 ;
        RECT 0.130 130.330 1.820 130.560 ;
        RECT 3.190 130.430 4.650 130.660 ;
        RECT 0.130 128.275 0.730 130.330 ;
        RECT 2.150 129.870 3.150 130.195 ;
        RECT 0.960 129.310 3.820 129.640 ;
        RECT 2.300 129.185 2.680 129.310 ;
        RECT 4.050 128.275 4.650 130.430 ;
        RECT 6.690 130.320 37.210 130.690 ;
        RECT 39.140 130.320 69.660 130.690 ;
        RECT 71.590 130.320 102.110 130.690 ;
        RECT 104.040 130.320 134.560 130.690 ;
        RECT 16.160 130.310 17.780 130.320 ;
        RECT 48.610 130.310 50.230 130.320 ;
        RECT 81.060 130.310 82.680 130.320 ;
        RECT 113.510 130.310 115.130 130.320 ;
        RECT 5.840 130.055 6.460 130.240 ;
        RECT 37.440 130.055 38.060 130.240 ;
        RECT 5.840 129.825 38.060 130.055 ;
        RECT 5.840 129.640 6.460 129.825 ;
        RECT 37.440 129.640 38.060 129.825 ;
        RECT 38.290 130.055 38.910 130.240 ;
        RECT 69.890 130.055 70.510 130.240 ;
        RECT 38.290 129.825 70.510 130.055 ;
        RECT 38.290 129.640 38.910 129.825 ;
        RECT 69.890 129.640 70.510 129.825 ;
        RECT 70.740 130.055 71.360 130.240 ;
        RECT 102.340 130.055 102.960 130.240 ;
        RECT 70.740 129.825 102.960 130.055 ;
        RECT 70.740 129.640 71.360 129.825 ;
        RECT 102.340 129.640 102.960 129.825 ;
        RECT 103.190 130.055 103.810 130.240 ;
        RECT 134.790 130.055 135.410 130.240 ;
        RECT 103.190 129.825 135.410 130.055 ;
        RECT 103.190 129.640 103.810 129.825 ;
        RECT 134.790 129.640 135.410 129.825 ;
        RECT 6.690 129.190 37.210 129.570 ;
        RECT 39.140 129.190 69.660 129.570 ;
        RECT 71.590 129.190 102.110 129.570 ;
        RECT 104.040 129.190 134.560 129.570 ;
        RECT 6.700 128.400 37.200 128.840 ;
        RECT 39.150 128.400 69.650 128.840 ;
        RECT 71.600 128.400 102.100 128.840 ;
        RECT 104.050 128.400 134.550 128.840 ;
        RECT 0.130 127.935 2.420 128.275 ;
        RECT 3.165 127.935 4.650 128.275 ;
        RECT 0.130 127.155 0.730 127.935 ;
        RECT 4.050 127.155 4.650 127.935 ;
        RECT 6.690 127.680 37.210 128.050 ;
        RECT 39.140 127.680 69.660 128.050 ;
        RECT 71.590 127.680 102.110 128.050 ;
        RECT 104.040 127.680 134.560 128.050 ;
        RECT 20.000 127.670 21.620 127.680 ;
        RECT 52.450 127.670 54.070 127.680 ;
        RECT 84.900 127.670 86.520 127.680 ;
        RECT 117.350 127.670 118.970 127.680 ;
        RECT 0.130 126.815 2.420 127.155 ;
        RECT 3.165 126.815 4.650 127.155 ;
        RECT 5.840 127.415 6.460 127.600 ;
        RECT 37.440 127.415 38.060 127.600 ;
        RECT 5.840 127.185 38.060 127.415 ;
        RECT 5.840 127.000 6.460 127.185 ;
        RECT 37.440 127.000 38.060 127.185 ;
        RECT 38.290 127.415 38.910 127.600 ;
        RECT 69.890 127.415 70.510 127.600 ;
        RECT 38.290 127.185 70.510 127.415 ;
        RECT 38.290 127.000 38.910 127.185 ;
        RECT 69.890 127.000 70.510 127.185 ;
        RECT 70.740 127.415 71.360 127.600 ;
        RECT 102.340 127.415 102.960 127.600 ;
        RECT 70.740 127.185 102.960 127.415 ;
        RECT 70.740 127.000 71.360 127.185 ;
        RECT 102.340 127.000 102.960 127.185 ;
        RECT 103.190 127.415 103.810 127.600 ;
        RECT 134.790 127.415 135.410 127.600 ;
        RECT 103.190 127.185 135.410 127.415 ;
        RECT 103.190 127.000 103.810 127.185 ;
        RECT 134.790 127.000 135.410 127.185 ;
        RECT 0.130 126.180 0.730 126.815 ;
        RECT 0.130 125.950 1.860 126.180 ;
        RECT 2.160 125.950 3.820 126.180 ;
        RECT 0.130 123.940 0.730 125.950 ;
        RECT 2.160 124.915 2.390 125.950 ;
        RECT 2.795 124.660 3.025 125.705 ;
        RECT 4.050 124.660 4.650 126.815 ;
        RECT 6.690 126.550 37.210 126.930 ;
        RECT 39.140 126.550 69.660 126.930 ;
        RECT 71.590 126.550 102.110 126.930 ;
        RECT 104.040 126.550 134.560 126.930 ;
        RECT 6.690 125.840 37.210 126.210 ;
        RECT 39.140 125.840 69.660 126.210 ;
        RECT 71.590 125.840 102.110 126.210 ;
        RECT 104.040 125.840 134.560 126.210 ;
        RECT 23.840 125.830 25.460 125.840 ;
        RECT 56.290 125.830 57.910 125.840 ;
        RECT 88.740 125.830 90.360 125.840 ;
        RECT 121.190 125.830 122.810 125.840 ;
        RECT 5.840 125.575 6.460 125.760 ;
        RECT 37.440 125.575 38.060 125.760 ;
        RECT 5.840 125.345 38.060 125.575 ;
        RECT 5.840 125.160 6.460 125.345 ;
        RECT 37.440 125.160 38.060 125.345 ;
        RECT 38.290 125.575 38.910 125.760 ;
        RECT 69.890 125.575 70.510 125.760 ;
        RECT 38.290 125.345 70.510 125.575 ;
        RECT 38.290 125.160 38.910 125.345 ;
        RECT 69.890 125.160 70.510 125.345 ;
        RECT 70.740 125.575 71.360 125.760 ;
        RECT 102.340 125.575 102.960 125.760 ;
        RECT 70.740 125.345 102.960 125.575 ;
        RECT 70.740 125.160 71.360 125.345 ;
        RECT 102.340 125.160 102.960 125.345 ;
        RECT 103.190 125.575 103.810 125.760 ;
        RECT 134.790 125.575 135.410 125.760 ;
        RECT 103.190 125.345 135.410 125.575 ;
        RECT 103.190 125.160 103.810 125.345 ;
        RECT 134.790 125.160 135.410 125.345 ;
        RECT 6.690 124.710 37.210 125.090 ;
        RECT 39.140 124.710 69.660 125.090 ;
        RECT 71.590 124.710 102.110 125.090 ;
        RECT 104.040 124.710 134.560 125.090 ;
        RECT 0.960 124.430 3.025 124.660 ;
        RECT 3.255 124.430 4.650 124.660 ;
        RECT 0.130 123.710 1.860 123.940 ;
        RECT 2.160 123.710 3.820 123.940 ;
        RECT 0.130 121.700 0.730 123.710 ;
        RECT 2.160 122.675 2.390 123.710 ;
        RECT 2.795 122.420 3.025 123.465 ;
        RECT 4.050 122.420 4.650 124.430 ;
        RECT 6.690 123.995 37.210 124.365 ;
        RECT 39.140 123.995 69.660 124.365 ;
        RECT 71.590 123.995 102.110 124.365 ;
        RECT 104.040 123.995 134.560 124.365 ;
        RECT 27.680 123.985 29.300 123.995 ;
        RECT 60.130 123.985 61.750 123.995 ;
        RECT 92.580 123.985 94.200 123.995 ;
        RECT 125.030 123.985 126.650 123.995 ;
        RECT 5.840 123.730 6.460 123.915 ;
        RECT 37.440 123.730 38.060 123.915 ;
        RECT 5.840 123.500 38.060 123.730 ;
        RECT 5.840 123.315 6.460 123.500 ;
        RECT 37.440 123.315 38.060 123.500 ;
        RECT 38.290 123.730 38.910 123.915 ;
        RECT 69.890 123.730 70.510 123.915 ;
        RECT 38.290 123.500 70.510 123.730 ;
        RECT 38.290 123.315 38.910 123.500 ;
        RECT 69.890 123.315 70.510 123.500 ;
        RECT 70.740 123.730 71.360 123.915 ;
        RECT 102.340 123.730 102.960 123.915 ;
        RECT 70.740 123.500 102.960 123.730 ;
        RECT 70.740 123.315 71.360 123.500 ;
        RECT 102.340 123.315 102.960 123.500 ;
        RECT 103.190 123.730 103.810 123.915 ;
        RECT 134.790 123.730 135.410 123.915 ;
        RECT 103.190 123.500 135.410 123.730 ;
        RECT 103.190 123.315 103.810 123.500 ;
        RECT 134.790 123.315 135.410 123.500 ;
        RECT 6.690 122.865 37.210 123.245 ;
        RECT 39.140 122.865 69.660 123.245 ;
        RECT 71.590 122.865 102.110 123.245 ;
        RECT 104.040 122.865 134.560 123.245 ;
        RECT 0.960 122.190 3.025 122.420 ;
        RECT 3.255 122.190 4.650 122.420 ;
        RECT 0.130 121.470 1.860 121.700 ;
        RECT 2.160 121.470 3.820 121.700 ;
        RECT 0.130 119.295 0.730 121.470 ;
        RECT 2.160 120.435 2.390 121.470 ;
        RECT 2.795 120.180 3.025 121.225 ;
        RECT 4.050 120.180 4.650 122.190 ;
        RECT 6.700 122.075 37.200 122.515 ;
        RECT 39.150 122.075 69.650 122.515 ;
        RECT 71.600 122.075 102.100 122.515 ;
        RECT 104.050 122.075 134.550 122.515 ;
        RECT 6.690 121.355 37.210 121.725 ;
        RECT 39.140 121.355 69.660 121.725 ;
        RECT 71.590 121.355 102.110 121.725 ;
        RECT 104.040 121.355 134.560 121.725 ;
        RECT 31.520 121.345 33.140 121.355 ;
        RECT 63.970 121.345 65.590 121.355 ;
        RECT 96.420 121.345 98.040 121.355 ;
        RECT 128.870 121.345 130.490 121.355 ;
        RECT 5.840 121.090 6.460 121.275 ;
        RECT 37.440 121.090 38.060 121.275 ;
        RECT 5.840 120.860 38.060 121.090 ;
        RECT 5.840 120.675 6.460 120.860 ;
        RECT 37.440 120.675 38.060 120.860 ;
        RECT 38.290 121.090 38.910 121.275 ;
        RECT 69.890 121.090 70.510 121.275 ;
        RECT 38.290 120.860 70.510 121.090 ;
        RECT 38.290 120.675 38.910 120.860 ;
        RECT 69.890 120.675 70.510 120.860 ;
        RECT 70.740 121.090 71.360 121.275 ;
        RECT 102.340 121.090 102.960 121.275 ;
        RECT 70.740 120.860 102.960 121.090 ;
        RECT 70.740 120.675 71.360 120.860 ;
        RECT 102.340 120.675 102.960 120.860 ;
        RECT 103.190 121.090 103.810 121.275 ;
        RECT 134.790 121.090 135.410 121.275 ;
        RECT 103.190 120.860 135.410 121.090 ;
        RECT 103.190 120.675 103.810 120.860 ;
        RECT 134.790 120.675 135.410 120.860 ;
        RECT 6.690 120.225 37.210 120.605 ;
        RECT 39.140 120.225 69.660 120.605 ;
        RECT 71.590 120.225 102.110 120.605 ;
        RECT 104.040 120.225 134.560 120.605 ;
        RECT 0.960 119.950 3.025 120.180 ;
        RECT 3.255 119.950 4.650 120.180 ;
        RECT 4.050 119.295 4.650 119.950 ;
        RECT 6.690 119.515 37.210 119.885 ;
        RECT 39.140 119.515 69.660 119.885 ;
        RECT 71.590 119.515 102.110 119.885 ;
        RECT 104.040 119.515 134.560 119.885 ;
        RECT 35.360 119.505 36.980 119.515 ;
        RECT 67.810 119.505 69.430 119.515 ;
        RECT 100.260 119.505 101.880 119.515 ;
        RECT 132.710 119.505 134.330 119.515 ;
        RECT 0.130 118.955 2.430 119.295 ;
        RECT 3.160 118.955 4.650 119.295 ;
        RECT 0.130 117.990 0.730 118.955 ;
        RECT 4.050 117.990 4.650 118.955 ;
        RECT 5.840 119.250 6.460 119.435 ;
        RECT 37.440 119.250 38.060 119.435 ;
        RECT 5.840 119.020 38.060 119.250 ;
        RECT 5.840 118.835 6.460 119.020 ;
        RECT 37.440 118.835 38.060 119.020 ;
        RECT 38.290 119.250 38.910 119.435 ;
        RECT 69.890 119.250 70.510 119.435 ;
        RECT 38.290 119.020 70.510 119.250 ;
        RECT 38.290 118.835 38.910 119.020 ;
        RECT 69.890 118.835 70.510 119.020 ;
        RECT 70.740 119.250 71.360 119.435 ;
        RECT 102.340 119.250 102.960 119.435 ;
        RECT 70.740 119.020 102.960 119.250 ;
        RECT 70.740 118.835 71.360 119.020 ;
        RECT 102.340 118.835 102.960 119.020 ;
        RECT 103.190 119.250 103.810 119.435 ;
        RECT 134.790 119.250 135.410 119.435 ;
        RECT 103.190 119.020 135.410 119.250 ;
        RECT 136.340 119.085 136.710 137.015 ;
        RECT 137.360 135.720 137.730 141.340 ;
        RECT 138.380 138.845 138.750 157.355 ;
        RECT 139.400 153.720 139.770 157.355 ;
        RECT 139.395 153.340 139.775 153.720 ;
        RECT 139.400 150.720 139.770 153.340 ;
        RECT 139.395 150.340 139.775 150.720 ;
        RECT 139.400 147.720 139.770 150.340 ;
        RECT 139.395 147.340 139.775 147.720 ;
        RECT 139.400 144.720 139.770 147.340 ;
        RECT 139.395 144.340 139.775 144.720 ;
        RECT 139.400 141.720 139.770 144.340 ;
        RECT 139.395 141.340 139.775 141.720 ;
        RECT 138.380 138.465 138.760 138.845 ;
        RECT 138.380 137.395 138.750 138.465 ;
        RECT 138.380 137.015 138.760 137.395 ;
        RECT 137.355 135.340 137.735 135.720 ;
        RECT 137.360 132.720 137.730 135.340 ;
        RECT 137.355 132.340 137.735 132.720 ;
        RECT 137.360 129.720 137.730 132.340 ;
        RECT 137.355 129.340 137.735 129.720 ;
        RECT 137.360 126.720 137.730 129.340 ;
        RECT 137.355 126.340 137.735 126.720 ;
        RECT 137.360 123.720 137.730 126.340 ;
        RECT 137.355 123.340 137.735 123.720 ;
        RECT 137.360 120.720 137.730 123.340 ;
        RECT 137.355 120.340 137.735 120.720 ;
        RECT 137.360 119.085 137.730 120.340 ;
        RECT 138.380 119.085 138.750 137.015 ;
        RECT 139.400 135.720 139.770 141.340 ;
        RECT 139.395 135.340 139.775 135.720 ;
        RECT 139.400 132.720 139.770 135.340 ;
        RECT 139.395 132.340 139.775 132.720 ;
        RECT 139.400 129.720 139.770 132.340 ;
        RECT 139.395 129.340 139.775 129.720 ;
        RECT 139.400 126.720 139.770 129.340 ;
        RECT 139.395 126.340 139.775 126.720 ;
        RECT 139.400 123.720 139.770 126.340 ;
        RECT 139.395 123.340 139.775 123.720 ;
        RECT 139.400 120.720 139.770 123.340 ;
        RECT 139.395 120.340 139.775 120.720 ;
        RECT 139.400 119.085 139.770 120.340 ;
        RECT 140.420 119.085 140.800 157.355 ;
        RECT 141.150 119.095 141.590 157.345 ;
        RECT 103.190 118.835 103.810 119.020 ;
        RECT 134.790 118.835 135.410 119.020 ;
        RECT 6.690 118.385 37.210 118.765 ;
        RECT 39.140 118.385 69.660 118.765 ;
        RECT 71.590 118.385 102.110 118.765 ;
        RECT 104.040 118.385 134.560 118.765 ;
        RECT 0.130 117.650 2.430 117.990 ;
        RECT 3.160 117.650 4.650 117.990 ;
        RECT 6.690 117.665 37.210 118.045 ;
        RECT 39.140 117.665 69.660 118.045 ;
        RECT 71.590 117.665 102.110 118.045 ;
        RECT 104.040 117.665 134.560 118.045 ;
        RECT 0.130 117.035 0.730 117.650 ;
        RECT 0.130 116.805 1.860 117.035 ;
        RECT 2.160 116.805 3.820 117.035 ;
        RECT 0.130 114.795 0.730 116.805 ;
        RECT 2.160 115.770 2.390 116.805 ;
        RECT 2.795 115.515 3.025 116.560 ;
        RECT 4.050 115.515 4.650 117.650 ;
        RECT 5.840 117.410 6.460 117.595 ;
        RECT 37.440 117.410 38.060 117.595 ;
        RECT 5.840 117.180 38.060 117.410 ;
        RECT 5.840 116.995 6.460 117.180 ;
        RECT 37.440 116.995 38.060 117.180 ;
        RECT 38.290 117.410 38.910 117.595 ;
        RECT 69.890 117.410 70.510 117.595 ;
        RECT 38.290 117.180 70.510 117.410 ;
        RECT 38.290 116.995 38.910 117.180 ;
        RECT 69.890 116.995 70.510 117.180 ;
        RECT 70.740 117.410 71.360 117.595 ;
        RECT 102.340 117.410 102.960 117.595 ;
        RECT 70.740 117.180 102.960 117.410 ;
        RECT 70.740 116.995 71.360 117.180 ;
        RECT 102.340 116.995 102.960 117.180 ;
        RECT 103.190 117.410 103.810 117.595 ;
        RECT 134.790 117.410 135.410 117.595 ;
        RECT 103.190 117.180 135.410 117.410 ;
        RECT 103.190 116.995 103.810 117.180 ;
        RECT 134.790 116.995 135.410 117.180 ;
        RECT 33.440 116.915 35.060 116.925 ;
        RECT 65.890 116.915 67.510 116.925 ;
        RECT 98.340 116.915 99.960 116.925 ;
        RECT 130.790 116.915 132.410 116.925 ;
        RECT 6.690 116.545 37.210 116.915 ;
        RECT 39.140 116.545 69.660 116.915 ;
        RECT 71.590 116.545 102.110 116.915 ;
        RECT 104.040 116.545 134.560 116.915 ;
        RECT 6.690 115.825 37.210 116.205 ;
        RECT 39.140 115.825 69.660 116.205 ;
        RECT 71.590 115.825 102.110 116.205 ;
        RECT 104.040 115.825 134.560 116.205 ;
        RECT 0.960 115.285 3.025 115.515 ;
        RECT 3.255 115.285 4.650 115.515 ;
        RECT 0.130 114.565 1.860 114.795 ;
        RECT 2.160 114.565 3.820 114.795 ;
        RECT 0.130 112.555 0.730 114.565 ;
        RECT 2.160 113.530 2.390 114.565 ;
        RECT 2.795 113.275 3.025 114.320 ;
        RECT 4.050 113.275 4.650 115.285 ;
        RECT 5.840 115.570 6.460 115.755 ;
        RECT 37.440 115.570 38.060 115.755 ;
        RECT 5.840 115.340 38.060 115.570 ;
        RECT 5.840 115.155 6.460 115.340 ;
        RECT 37.440 115.155 38.060 115.340 ;
        RECT 38.290 115.570 38.910 115.755 ;
        RECT 69.890 115.570 70.510 115.755 ;
        RECT 38.290 115.340 70.510 115.570 ;
        RECT 38.290 115.155 38.910 115.340 ;
        RECT 69.890 115.155 70.510 115.340 ;
        RECT 70.740 115.570 71.360 115.755 ;
        RECT 102.340 115.570 102.960 115.755 ;
        RECT 70.740 115.340 102.960 115.570 ;
        RECT 70.740 115.155 71.360 115.340 ;
        RECT 102.340 115.155 102.960 115.340 ;
        RECT 103.190 115.570 103.810 115.755 ;
        RECT 134.790 115.570 135.410 115.755 ;
        RECT 103.190 115.340 135.410 115.570 ;
        RECT 103.190 115.155 103.810 115.340 ;
        RECT 134.790 115.155 135.410 115.340 ;
        RECT 29.600 115.075 31.220 115.085 ;
        RECT 62.050 115.075 63.670 115.085 ;
        RECT 94.500 115.075 96.120 115.085 ;
        RECT 126.950 115.075 128.570 115.085 ;
        RECT 6.690 114.705 37.210 115.075 ;
        RECT 39.140 114.705 69.660 115.075 ;
        RECT 71.590 114.705 102.110 115.075 ;
        RECT 104.040 114.705 134.560 115.075 ;
        RECT 6.700 113.910 37.200 114.350 ;
        RECT 39.150 113.910 69.650 114.350 ;
        RECT 71.600 113.910 102.100 114.350 ;
        RECT 104.050 113.910 134.550 114.350 ;
        RECT 0.960 113.045 3.025 113.275 ;
        RECT 3.255 113.045 4.650 113.275 ;
        RECT 6.690 113.180 37.210 113.560 ;
        RECT 39.140 113.180 69.660 113.560 ;
        RECT 71.590 113.180 102.110 113.560 ;
        RECT 104.040 113.180 134.560 113.560 ;
        RECT 0.130 112.325 1.860 112.555 ;
        RECT 2.160 112.325 3.820 112.555 ;
        RECT 0.130 110.315 0.730 112.325 ;
        RECT 2.160 111.290 2.390 112.325 ;
        RECT 2.795 111.035 3.025 112.080 ;
        RECT 4.050 111.035 4.650 113.045 ;
        RECT 5.840 112.925 6.460 113.110 ;
        RECT 37.440 112.925 38.060 113.110 ;
        RECT 5.840 112.695 38.060 112.925 ;
        RECT 5.840 112.510 6.460 112.695 ;
        RECT 37.440 112.510 38.060 112.695 ;
        RECT 38.290 112.925 38.910 113.110 ;
        RECT 69.890 112.925 70.510 113.110 ;
        RECT 38.290 112.695 70.510 112.925 ;
        RECT 38.290 112.510 38.910 112.695 ;
        RECT 69.890 112.510 70.510 112.695 ;
        RECT 70.740 112.925 71.360 113.110 ;
        RECT 102.340 112.925 102.960 113.110 ;
        RECT 70.740 112.695 102.960 112.925 ;
        RECT 70.740 112.510 71.360 112.695 ;
        RECT 102.340 112.510 102.960 112.695 ;
        RECT 103.190 112.925 103.810 113.110 ;
        RECT 134.790 112.925 135.410 113.110 ;
        RECT 103.190 112.695 135.410 112.925 ;
        RECT 103.190 112.510 103.810 112.695 ;
        RECT 134.790 112.510 135.410 112.695 ;
        RECT 25.760 112.430 27.380 112.440 ;
        RECT 58.210 112.430 59.830 112.440 ;
        RECT 90.660 112.430 92.280 112.440 ;
        RECT 123.110 112.430 124.730 112.440 ;
        RECT 6.690 112.060 37.210 112.430 ;
        RECT 39.140 112.060 69.660 112.430 ;
        RECT 71.590 112.060 102.110 112.430 ;
        RECT 104.040 112.060 134.560 112.430 ;
        RECT 6.690 111.340 37.210 111.720 ;
        RECT 39.140 111.340 69.660 111.720 ;
        RECT 71.590 111.340 102.110 111.720 ;
        RECT 104.040 111.340 134.560 111.720 ;
        RECT 0.960 110.805 3.025 111.035 ;
        RECT 3.255 110.805 4.650 111.035 ;
        RECT 0.130 110.085 1.860 110.315 ;
        RECT 2.160 110.085 3.820 110.315 ;
        RECT 0.130 108.075 0.730 110.085 ;
        RECT 2.160 109.050 2.390 110.085 ;
        RECT 2.795 108.795 3.025 109.840 ;
        RECT 4.050 108.795 4.650 110.805 ;
        RECT 5.840 111.085 6.460 111.270 ;
        RECT 37.440 111.085 38.060 111.270 ;
        RECT 5.840 110.855 38.060 111.085 ;
        RECT 5.840 110.670 6.460 110.855 ;
        RECT 37.440 110.670 38.060 110.855 ;
        RECT 38.290 111.085 38.910 111.270 ;
        RECT 69.890 111.085 70.510 111.270 ;
        RECT 38.290 110.855 70.510 111.085 ;
        RECT 38.290 110.670 38.910 110.855 ;
        RECT 69.890 110.670 70.510 110.855 ;
        RECT 70.740 111.085 71.360 111.270 ;
        RECT 102.340 111.085 102.960 111.270 ;
        RECT 70.740 110.855 102.960 111.085 ;
        RECT 70.740 110.670 71.360 110.855 ;
        RECT 102.340 110.670 102.960 110.855 ;
        RECT 103.190 111.085 103.810 111.270 ;
        RECT 134.790 111.085 135.410 111.270 ;
        RECT 103.190 110.855 135.410 111.085 ;
        RECT 103.190 110.670 103.810 110.855 ;
        RECT 134.790 110.670 135.410 110.855 ;
        RECT 21.920 110.590 23.540 110.600 ;
        RECT 54.370 110.590 55.990 110.600 ;
        RECT 86.820 110.590 88.440 110.600 ;
        RECT 119.270 110.590 120.890 110.600 ;
        RECT 6.690 110.220 37.210 110.590 ;
        RECT 39.140 110.220 69.660 110.590 ;
        RECT 71.590 110.220 102.110 110.590 ;
        RECT 104.040 110.220 134.560 110.590 ;
        RECT 6.690 109.500 37.210 109.880 ;
        RECT 39.140 109.500 69.660 109.880 ;
        RECT 71.590 109.500 102.110 109.880 ;
        RECT 104.040 109.500 134.560 109.880 ;
        RECT 5.840 109.245 6.460 109.430 ;
        RECT 37.440 109.245 38.060 109.430 ;
        RECT 5.840 109.015 38.060 109.245 ;
        RECT 5.840 108.830 6.460 109.015 ;
        RECT 37.440 108.830 38.060 109.015 ;
        RECT 38.290 109.245 38.910 109.430 ;
        RECT 69.890 109.245 70.510 109.430 ;
        RECT 38.290 109.015 70.510 109.245 ;
        RECT 38.290 108.830 38.910 109.015 ;
        RECT 69.890 108.830 70.510 109.015 ;
        RECT 70.740 109.245 71.360 109.430 ;
        RECT 102.340 109.245 102.960 109.430 ;
        RECT 70.740 109.015 102.960 109.245 ;
        RECT 70.740 108.830 71.360 109.015 ;
        RECT 102.340 108.830 102.960 109.015 ;
        RECT 103.190 109.245 103.810 109.430 ;
        RECT 134.790 109.245 135.410 109.430 ;
        RECT 103.190 109.015 135.410 109.245 ;
        RECT 103.190 108.830 103.810 109.015 ;
        RECT 134.790 108.830 135.410 109.015 ;
        RECT 0.960 108.565 3.025 108.795 ;
        RECT 3.255 108.565 4.650 108.795 ;
        RECT 18.080 108.750 19.700 108.760 ;
        RECT 50.530 108.750 52.150 108.760 ;
        RECT 82.980 108.750 84.600 108.760 ;
        RECT 115.430 108.750 117.050 108.760 ;
        RECT 0.130 107.845 1.860 108.075 ;
        RECT 2.160 107.845 3.820 108.075 ;
        RECT 0.130 105.690 0.730 107.845 ;
        RECT 2.160 106.810 2.390 107.845 ;
        RECT 2.795 106.555 3.025 107.600 ;
        RECT 4.050 106.555 4.650 108.565 ;
        RECT 6.690 108.380 37.210 108.750 ;
        RECT 39.140 108.380 69.660 108.750 ;
        RECT 71.590 108.380 102.110 108.750 ;
        RECT 104.040 108.380 134.560 108.750 ;
        RECT 6.700 107.585 37.200 108.025 ;
        RECT 39.150 107.585 69.650 108.025 ;
        RECT 71.600 107.585 102.100 108.025 ;
        RECT 104.050 107.585 134.550 108.025 ;
        RECT 6.690 106.855 37.210 107.235 ;
        RECT 39.140 106.855 69.660 107.235 ;
        RECT 71.590 106.855 102.110 107.235 ;
        RECT 104.040 106.855 134.560 107.235 ;
        RECT 0.960 106.325 3.025 106.555 ;
        RECT 3.255 106.325 4.650 106.555 ;
        RECT 4.050 105.690 4.650 106.325 ;
        RECT 5.840 106.600 6.460 106.785 ;
        RECT 37.440 106.600 38.060 106.785 ;
        RECT 5.840 106.370 38.060 106.600 ;
        RECT 5.840 106.185 6.460 106.370 ;
        RECT 37.440 106.185 38.060 106.370 ;
        RECT 38.290 106.600 38.910 106.785 ;
        RECT 69.890 106.600 70.510 106.785 ;
        RECT 38.290 106.370 70.510 106.600 ;
        RECT 38.290 106.185 38.910 106.370 ;
        RECT 69.890 106.185 70.510 106.370 ;
        RECT 70.740 106.600 71.360 106.785 ;
        RECT 102.340 106.600 102.960 106.785 ;
        RECT 70.740 106.370 102.960 106.600 ;
        RECT 70.740 106.185 71.360 106.370 ;
        RECT 102.340 106.185 102.960 106.370 ;
        RECT 103.190 106.600 103.810 106.785 ;
        RECT 134.790 106.600 135.410 106.785 ;
        RECT 103.190 106.370 135.410 106.600 ;
        RECT 103.190 106.185 103.810 106.370 ;
        RECT 134.790 106.185 135.410 106.370 ;
        RECT 14.240 106.105 15.860 106.115 ;
        RECT 46.690 106.105 48.310 106.115 ;
        RECT 79.140 106.105 80.760 106.115 ;
        RECT 111.590 106.105 113.210 106.115 ;
        RECT 6.690 105.735 37.210 106.105 ;
        RECT 39.140 105.735 69.660 106.105 ;
        RECT 71.590 105.735 102.110 106.105 ;
        RECT 104.040 105.735 134.560 106.105 ;
        RECT 0.130 105.350 2.420 105.690 ;
        RECT 3.165 105.350 4.650 105.690 ;
        RECT 0.130 104.715 0.730 105.350 ;
        RECT 0.130 104.485 1.860 104.715 ;
        RECT 2.160 104.485 3.820 104.715 ;
        RECT 0.130 102.475 0.730 104.485 ;
        RECT 2.160 103.450 2.390 104.485 ;
        RECT 2.795 103.195 3.025 104.240 ;
        RECT 4.050 103.195 4.650 105.350 ;
        RECT 6.690 105.015 37.210 105.395 ;
        RECT 39.140 105.015 69.660 105.395 ;
        RECT 71.590 105.015 102.110 105.395 ;
        RECT 104.040 105.015 134.560 105.395 ;
        RECT 5.840 104.760 6.460 104.945 ;
        RECT 37.440 104.760 38.060 104.945 ;
        RECT 5.840 104.530 38.060 104.760 ;
        RECT 5.840 104.345 6.460 104.530 ;
        RECT 37.440 104.345 38.060 104.530 ;
        RECT 38.290 104.760 38.910 104.945 ;
        RECT 69.890 104.760 70.510 104.945 ;
        RECT 38.290 104.530 70.510 104.760 ;
        RECT 38.290 104.345 38.910 104.530 ;
        RECT 69.890 104.345 70.510 104.530 ;
        RECT 70.740 104.760 71.360 104.945 ;
        RECT 102.340 104.760 102.960 104.945 ;
        RECT 70.740 104.530 102.960 104.760 ;
        RECT 70.740 104.345 71.360 104.530 ;
        RECT 102.340 104.345 102.960 104.530 ;
        RECT 103.190 104.760 103.810 104.945 ;
        RECT 134.790 104.760 135.410 104.945 ;
        RECT 103.190 104.530 135.410 104.760 ;
        RECT 103.190 104.345 103.810 104.530 ;
        RECT 134.790 104.345 135.410 104.530 ;
        RECT 10.400 104.265 12.020 104.275 ;
        RECT 42.850 104.265 44.470 104.275 ;
        RECT 75.300 104.265 76.920 104.275 ;
        RECT 107.750 104.265 109.370 104.275 ;
        RECT 6.690 103.895 37.210 104.265 ;
        RECT 39.140 103.895 69.660 104.265 ;
        RECT 71.590 103.895 102.110 104.265 ;
        RECT 104.040 103.895 134.560 104.265 ;
        RECT 0.960 102.965 3.025 103.195 ;
        RECT 3.255 102.965 4.650 103.195 ;
        RECT 6.690 103.175 37.210 103.555 ;
        RECT 39.140 103.175 69.660 103.555 ;
        RECT 71.590 103.175 102.110 103.555 ;
        RECT 104.040 103.175 134.560 103.555 ;
        RECT 0.130 102.245 1.860 102.475 ;
        RECT 2.160 102.245 3.820 102.475 ;
        RECT 0.130 100.090 0.730 102.245 ;
        RECT 2.160 101.210 2.390 102.245 ;
        RECT 2.795 100.955 3.025 102.000 ;
        RECT 4.050 100.955 4.650 102.965 ;
        RECT 5.840 102.920 6.460 103.105 ;
        RECT 37.440 102.920 38.060 103.105 ;
        RECT 5.840 102.690 38.060 102.920 ;
        RECT 5.840 102.505 6.460 102.690 ;
        RECT 37.440 102.505 38.060 102.690 ;
        RECT 38.290 102.920 38.910 103.105 ;
        RECT 69.890 102.920 70.510 103.105 ;
        RECT 38.290 102.690 70.510 102.920 ;
        RECT 38.290 102.505 38.910 102.690 ;
        RECT 69.890 102.505 70.510 102.690 ;
        RECT 70.740 102.920 71.360 103.105 ;
        RECT 102.340 102.920 102.960 103.105 ;
        RECT 70.740 102.690 102.960 102.920 ;
        RECT 70.740 102.505 71.360 102.690 ;
        RECT 102.340 102.505 102.960 102.690 ;
        RECT 103.190 102.920 103.810 103.105 ;
        RECT 134.790 102.920 135.410 103.105 ;
        RECT 103.190 102.690 135.410 102.920 ;
        RECT 103.190 102.505 103.810 102.690 ;
        RECT 134.790 102.505 135.410 102.690 ;
        RECT 6.690 102.055 37.210 102.425 ;
        RECT 39.140 102.055 69.660 102.425 ;
        RECT 71.590 102.055 102.110 102.425 ;
        RECT 104.040 102.055 134.560 102.425 ;
        RECT 0.960 100.725 3.025 100.955 ;
        RECT 3.255 100.725 4.650 100.955 ;
        RECT 4.050 100.090 4.650 100.725 ;
        RECT 0.130 99.750 2.420 100.090 ;
        RECT 3.165 99.750 4.650 100.090 ;
        RECT 0.130 99.115 0.730 99.750 ;
        RECT 0.130 98.885 1.710 99.115 ;
        RECT 0.130 96.845 0.730 98.885 ;
        RECT 2.140 98.655 2.500 98.740 ;
        RECT 1.010 98.425 2.500 98.655 ;
        RECT 1.010 98.275 1.370 98.425 ;
        RECT 0.960 97.640 1.910 98.045 ;
        RECT 0.130 96.615 1.420 96.845 ;
        RECT 0.130 95.655 0.730 96.615 ;
        RECT 1.650 96.295 1.910 97.640 ;
        RECT 2.140 96.990 2.500 98.425 ;
        RECT 2.730 97.090 3.080 98.290 ;
        RECT 3.440 97.680 3.820 99.325 ;
        RECT 2.520 96.295 2.870 96.355 ;
        RECT 3.440 96.295 3.780 96.900 ;
        RECT 1.650 96.035 3.780 96.295 ;
        RECT 2.520 95.975 2.870 96.035 ;
        RECT 4.050 95.755 4.650 99.750 ;
        RECT 6.495 99.270 8.245 102.055 ;
        RECT 8.885 99.270 9.695 100.270 ;
        RECT 10.335 99.270 12.085 101.565 ;
        RECT 12.725 99.270 13.535 100.270 ;
        RECT 14.175 99.270 15.925 101.565 ;
        RECT 16.565 99.270 17.375 100.270 ;
        RECT 18.015 99.270 19.765 101.565 ;
        RECT 20.405 99.270 21.215 100.270 ;
        RECT 21.855 99.270 23.605 101.565 ;
        RECT 24.245 99.270 25.055 100.270 ;
        RECT 25.695 99.270 27.445 101.565 ;
        RECT 28.085 99.270 28.895 100.270 ;
        RECT 29.535 99.270 31.285 101.565 ;
        RECT 31.925 99.270 32.735 100.270 ;
        RECT 33.375 99.270 35.125 101.565 ;
        RECT 35.765 99.270 36.575 100.270 ;
        RECT 38.945 99.270 40.695 102.055 ;
        RECT 41.335 99.270 42.145 100.270 ;
        RECT 42.785 99.270 44.535 101.565 ;
        RECT 45.175 99.270 45.985 100.270 ;
        RECT 46.625 99.270 48.375 101.565 ;
        RECT 49.015 99.270 49.825 100.270 ;
        RECT 50.465 99.270 52.215 101.565 ;
        RECT 52.855 99.270 53.665 100.270 ;
        RECT 54.305 99.270 56.055 101.565 ;
        RECT 56.695 99.270 57.505 100.270 ;
        RECT 58.145 99.270 59.895 101.565 ;
        RECT 60.535 99.270 61.345 100.270 ;
        RECT 61.985 99.270 63.735 101.565 ;
        RECT 64.375 99.270 65.185 100.270 ;
        RECT 65.825 99.270 67.575 101.565 ;
        RECT 68.215 99.270 69.025 100.270 ;
        RECT 71.395 99.270 73.145 102.055 ;
        RECT 73.785 99.270 74.595 100.270 ;
        RECT 75.235 99.270 76.985 101.565 ;
        RECT 77.625 99.270 78.435 100.270 ;
        RECT 79.075 99.270 80.825 101.565 ;
        RECT 81.465 99.270 82.275 100.270 ;
        RECT 82.915 99.270 84.665 101.565 ;
        RECT 85.305 99.270 86.115 100.270 ;
        RECT 86.755 99.270 88.505 101.565 ;
        RECT 89.145 99.270 89.955 100.270 ;
        RECT 90.595 99.270 92.345 101.565 ;
        RECT 92.985 99.270 93.795 100.270 ;
        RECT 94.435 99.270 96.185 101.565 ;
        RECT 96.825 99.270 97.635 100.270 ;
        RECT 98.275 99.270 100.025 101.565 ;
        RECT 100.665 99.270 101.475 100.270 ;
        RECT 103.845 99.270 105.595 102.055 ;
        RECT 106.235 99.270 107.045 100.270 ;
        RECT 107.685 99.270 109.435 101.565 ;
        RECT 110.075 99.270 110.885 100.270 ;
        RECT 111.525 99.270 113.275 101.565 ;
        RECT 113.915 99.270 114.725 100.270 ;
        RECT 115.365 99.270 117.115 101.565 ;
        RECT 117.755 99.270 118.565 100.270 ;
        RECT 119.205 99.270 120.955 101.565 ;
        RECT 121.595 99.270 122.405 100.270 ;
        RECT 123.045 99.270 124.795 101.565 ;
        RECT 125.435 99.270 126.245 100.270 ;
        RECT 126.885 99.270 128.635 101.565 ;
        RECT 129.275 99.270 130.085 100.270 ;
        RECT 130.725 99.270 132.475 101.565 ;
        RECT 133.115 99.270 133.925 100.270 ;
        RECT 136.340 99.460 136.710 117.970 ;
        RECT 137.360 114.335 137.730 117.970 ;
        RECT 137.355 113.955 137.735 114.335 ;
        RECT 137.360 111.335 137.730 113.955 ;
        RECT 137.355 110.955 137.735 111.335 ;
        RECT 137.360 108.335 137.730 110.955 ;
        RECT 137.355 107.955 137.735 108.335 ;
        RECT 137.360 105.335 137.730 107.955 ;
        RECT 137.355 104.955 137.735 105.335 ;
        RECT 137.360 102.335 137.730 104.955 ;
        RECT 137.355 101.955 137.735 102.335 ;
        RECT 136.340 99.080 136.720 99.460 ;
        RECT 136.340 98.010 136.710 99.080 ;
        RECT 6.965 96.820 7.775 97.820 ;
        RECT 0.130 95.425 1.820 95.655 ;
        RECT 3.190 95.525 4.650 95.755 ;
        RECT 0.130 93.415 0.730 95.425 ;
        RECT 2.150 94.965 3.150 95.290 ;
        RECT 0.960 94.405 3.820 94.735 ;
        RECT 0.130 93.185 1.820 93.415 ;
        RECT 0.130 91.175 0.730 93.185 ;
        RECT 2.535 93.050 2.800 94.405 ;
        RECT 4.050 93.515 4.650 95.525 ;
        RECT 8.415 94.990 10.165 97.820 ;
        RECT 10.805 96.820 11.615 97.820 ;
        RECT 12.255 95.525 14.005 97.820 ;
        RECT 14.645 96.820 15.455 97.820 ;
        RECT 16.095 95.525 17.845 97.820 ;
        RECT 18.485 96.820 19.295 97.820 ;
        RECT 19.935 95.525 21.685 97.820 ;
        RECT 22.325 96.820 23.135 97.820 ;
        RECT 23.775 95.525 25.525 97.820 ;
        RECT 26.165 96.820 26.975 97.820 ;
        RECT 27.615 95.525 29.365 97.820 ;
        RECT 30.005 96.820 30.815 97.820 ;
        RECT 31.455 95.525 33.205 97.820 ;
        RECT 33.845 96.820 34.655 97.820 ;
        RECT 35.295 95.525 37.045 97.820 ;
        RECT 39.415 96.820 40.225 97.820 ;
        RECT 40.865 94.990 42.615 97.820 ;
        RECT 43.255 96.820 44.065 97.820 ;
        RECT 44.705 95.525 46.455 97.820 ;
        RECT 47.095 96.820 47.905 97.820 ;
        RECT 48.545 95.525 50.295 97.820 ;
        RECT 50.935 96.820 51.745 97.820 ;
        RECT 52.385 95.525 54.135 97.820 ;
        RECT 54.775 96.820 55.585 97.820 ;
        RECT 56.225 95.525 57.975 97.820 ;
        RECT 58.615 96.820 59.425 97.820 ;
        RECT 60.065 95.525 61.815 97.820 ;
        RECT 62.455 96.820 63.265 97.820 ;
        RECT 63.905 95.525 65.655 97.820 ;
        RECT 66.295 96.820 67.105 97.820 ;
        RECT 67.745 95.525 69.495 97.820 ;
        RECT 71.865 96.820 72.675 97.820 ;
        RECT 73.315 94.990 75.065 97.820 ;
        RECT 75.705 96.820 76.515 97.820 ;
        RECT 77.155 95.525 78.905 97.820 ;
        RECT 79.545 96.820 80.355 97.820 ;
        RECT 80.995 95.525 82.745 97.820 ;
        RECT 83.385 96.820 84.195 97.820 ;
        RECT 84.835 95.525 86.585 97.820 ;
        RECT 87.225 96.820 88.035 97.820 ;
        RECT 88.675 95.525 90.425 97.820 ;
        RECT 91.065 96.820 91.875 97.820 ;
        RECT 92.515 95.525 94.265 97.820 ;
        RECT 94.905 96.820 95.715 97.820 ;
        RECT 96.355 95.525 98.105 97.820 ;
        RECT 98.745 96.820 99.555 97.820 ;
        RECT 100.195 95.525 101.945 97.820 ;
        RECT 104.315 96.820 105.125 97.820 ;
        RECT 105.765 94.990 107.515 97.820 ;
        RECT 108.155 96.820 108.965 97.820 ;
        RECT 109.605 95.525 111.355 97.820 ;
        RECT 111.995 96.820 112.805 97.820 ;
        RECT 113.445 95.525 115.195 97.820 ;
        RECT 115.835 96.820 116.645 97.820 ;
        RECT 117.285 95.525 119.035 97.820 ;
        RECT 119.675 96.820 120.485 97.820 ;
        RECT 121.125 95.525 122.875 97.820 ;
        RECT 123.515 96.820 124.325 97.820 ;
        RECT 124.965 95.525 126.715 97.820 ;
        RECT 127.355 96.820 128.165 97.820 ;
        RECT 128.805 95.525 130.555 97.820 ;
        RECT 131.195 96.820 132.005 97.820 ;
        RECT 132.645 95.525 134.395 97.820 ;
        RECT 136.340 97.630 136.720 98.010 ;
        RECT 6.690 94.620 37.210 94.990 ;
        RECT 39.140 94.620 69.660 94.990 ;
        RECT 71.590 94.620 102.110 94.990 ;
        RECT 104.040 94.620 134.560 94.990 ;
        RECT 5.840 94.355 6.460 94.540 ;
        RECT 37.440 94.355 38.060 94.540 ;
        RECT 5.840 94.125 38.060 94.355 ;
        RECT 5.840 93.940 6.460 94.125 ;
        RECT 37.440 93.940 38.060 94.125 ;
        RECT 38.290 94.355 38.910 94.540 ;
        RECT 69.890 94.355 70.510 94.540 ;
        RECT 38.290 94.125 70.510 94.355 ;
        RECT 38.290 93.940 38.910 94.125 ;
        RECT 69.890 93.940 70.510 94.125 ;
        RECT 70.740 94.355 71.360 94.540 ;
        RECT 102.340 94.355 102.960 94.540 ;
        RECT 70.740 94.125 102.960 94.355 ;
        RECT 70.740 93.940 71.360 94.125 ;
        RECT 102.340 93.940 102.960 94.125 ;
        RECT 103.190 94.355 103.810 94.540 ;
        RECT 134.790 94.355 135.410 94.540 ;
        RECT 103.190 94.125 135.410 94.355 ;
        RECT 103.190 93.940 103.810 94.125 ;
        RECT 134.790 93.940 135.410 94.125 ;
        RECT 3.190 93.285 4.650 93.515 ;
        RECT 6.690 93.490 37.210 93.870 ;
        RECT 39.140 93.490 69.660 93.870 ;
        RECT 71.590 93.490 102.110 93.870 ;
        RECT 104.040 93.490 134.560 93.870 ;
        RECT 2.150 92.725 3.150 93.050 ;
        RECT 0.960 92.165 3.820 92.495 ;
        RECT 4.050 91.275 4.650 93.285 ;
        RECT 6.690 92.780 37.210 93.150 ;
        RECT 39.140 92.780 69.660 93.150 ;
        RECT 71.590 92.780 102.110 93.150 ;
        RECT 104.040 92.780 134.560 93.150 ;
        RECT 12.320 92.770 13.940 92.780 ;
        RECT 44.770 92.770 46.390 92.780 ;
        RECT 77.220 92.770 78.840 92.780 ;
        RECT 109.670 92.770 111.290 92.780 ;
        RECT 5.840 92.515 6.460 92.700 ;
        RECT 37.440 92.515 38.060 92.700 ;
        RECT 5.840 92.285 38.060 92.515 ;
        RECT 5.840 92.100 6.460 92.285 ;
        RECT 37.440 92.100 38.060 92.285 ;
        RECT 38.290 92.515 38.910 92.700 ;
        RECT 69.890 92.515 70.510 92.700 ;
        RECT 38.290 92.285 70.510 92.515 ;
        RECT 38.290 92.100 38.910 92.285 ;
        RECT 69.890 92.100 70.510 92.285 ;
        RECT 70.740 92.515 71.360 92.700 ;
        RECT 102.340 92.515 102.960 92.700 ;
        RECT 70.740 92.285 102.960 92.515 ;
        RECT 70.740 92.100 71.360 92.285 ;
        RECT 102.340 92.100 102.960 92.285 ;
        RECT 103.190 92.515 103.810 92.700 ;
        RECT 134.790 92.515 135.410 92.700 ;
        RECT 103.190 92.285 135.410 92.515 ;
        RECT 103.190 92.100 103.810 92.285 ;
        RECT 134.790 92.100 135.410 92.285 ;
        RECT 6.690 91.650 37.210 92.030 ;
        RECT 39.140 91.650 69.660 92.030 ;
        RECT 71.590 91.650 102.110 92.030 ;
        RECT 104.040 91.650 134.560 92.030 ;
        RECT 0.130 90.945 1.820 91.175 ;
        RECT 3.190 91.045 4.650 91.275 ;
        RECT 0.130 88.890 0.730 90.945 ;
        RECT 2.150 90.485 3.150 90.810 ;
        RECT 0.960 89.925 3.820 90.255 ;
        RECT 2.300 89.800 2.680 89.925 ;
        RECT 4.050 88.890 4.650 91.045 ;
        RECT 6.690 90.935 37.210 91.305 ;
        RECT 39.140 90.935 69.660 91.305 ;
        RECT 71.590 90.935 102.110 91.305 ;
        RECT 104.040 90.935 134.560 91.305 ;
        RECT 16.160 90.925 17.780 90.935 ;
        RECT 48.610 90.925 50.230 90.935 ;
        RECT 81.060 90.925 82.680 90.935 ;
        RECT 113.510 90.925 115.130 90.935 ;
        RECT 5.840 90.670 6.460 90.855 ;
        RECT 37.440 90.670 38.060 90.855 ;
        RECT 5.840 90.440 38.060 90.670 ;
        RECT 5.840 90.255 6.460 90.440 ;
        RECT 37.440 90.255 38.060 90.440 ;
        RECT 38.290 90.670 38.910 90.855 ;
        RECT 69.890 90.670 70.510 90.855 ;
        RECT 38.290 90.440 70.510 90.670 ;
        RECT 38.290 90.255 38.910 90.440 ;
        RECT 69.890 90.255 70.510 90.440 ;
        RECT 70.740 90.670 71.360 90.855 ;
        RECT 102.340 90.670 102.960 90.855 ;
        RECT 70.740 90.440 102.960 90.670 ;
        RECT 70.740 90.255 71.360 90.440 ;
        RECT 102.340 90.255 102.960 90.440 ;
        RECT 103.190 90.670 103.810 90.855 ;
        RECT 134.790 90.670 135.410 90.855 ;
        RECT 103.190 90.440 135.410 90.670 ;
        RECT 103.190 90.255 103.810 90.440 ;
        RECT 134.790 90.255 135.410 90.440 ;
        RECT 6.690 89.805 37.210 90.185 ;
        RECT 39.140 89.805 69.660 90.185 ;
        RECT 71.590 89.805 102.110 90.185 ;
        RECT 104.040 89.805 134.560 90.185 ;
        RECT 6.700 89.015 37.200 89.455 ;
        RECT 39.150 89.015 69.650 89.455 ;
        RECT 71.600 89.015 102.100 89.455 ;
        RECT 104.050 89.015 134.550 89.455 ;
        RECT 0.130 88.550 2.420 88.890 ;
        RECT 3.165 88.550 4.650 88.890 ;
        RECT 0.130 87.770 0.730 88.550 ;
        RECT 4.050 87.770 4.650 88.550 ;
        RECT 6.690 88.295 37.210 88.665 ;
        RECT 39.140 88.295 69.660 88.665 ;
        RECT 71.590 88.295 102.110 88.665 ;
        RECT 104.040 88.295 134.560 88.665 ;
        RECT 20.000 88.285 21.620 88.295 ;
        RECT 52.450 88.285 54.070 88.295 ;
        RECT 84.900 88.285 86.520 88.295 ;
        RECT 117.350 88.285 118.970 88.295 ;
        RECT 0.130 87.430 2.420 87.770 ;
        RECT 3.165 87.430 4.650 87.770 ;
        RECT 5.840 88.030 6.460 88.215 ;
        RECT 37.440 88.030 38.060 88.215 ;
        RECT 5.840 87.800 38.060 88.030 ;
        RECT 5.840 87.615 6.460 87.800 ;
        RECT 37.440 87.615 38.060 87.800 ;
        RECT 38.290 88.030 38.910 88.215 ;
        RECT 69.890 88.030 70.510 88.215 ;
        RECT 38.290 87.800 70.510 88.030 ;
        RECT 38.290 87.615 38.910 87.800 ;
        RECT 69.890 87.615 70.510 87.800 ;
        RECT 70.740 88.030 71.360 88.215 ;
        RECT 102.340 88.030 102.960 88.215 ;
        RECT 70.740 87.800 102.960 88.030 ;
        RECT 70.740 87.615 71.360 87.800 ;
        RECT 102.340 87.615 102.960 87.800 ;
        RECT 103.190 88.030 103.810 88.215 ;
        RECT 134.790 88.030 135.410 88.215 ;
        RECT 103.190 87.800 135.410 88.030 ;
        RECT 103.190 87.615 103.810 87.800 ;
        RECT 134.790 87.615 135.410 87.800 ;
        RECT 0.130 86.795 0.730 87.430 ;
        RECT 0.130 86.565 1.860 86.795 ;
        RECT 2.160 86.565 3.820 86.795 ;
        RECT 0.130 84.555 0.730 86.565 ;
        RECT 2.160 85.530 2.390 86.565 ;
        RECT 2.795 85.275 3.025 86.320 ;
        RECT 4.050 85.275 4.650 87.430 ;
        RECT 6.690 87.165 37.210 87.545 ;
        RECT 39.140 87.165 69.660 87.545 ;
        RECT 71.590 87.165 102.110 87.545 ;
        RECT 104.040 87.165 134.560 87.545 ;
        RECT 6.690 86.455 37.210 86.825 ;
        RECT 39.140 86.455 69.660 86.825 ;
        RECT 71.590 86.455 102.110 86.825 ;
        RECT 104.040 86.455 134.560 86.825 ;
        RECT 23.840 86.445 25.460 86.455 ;
        RECT 56.290 86.445 57.910 86.455 ;
        RECT 88.740 86.445 90.360 86.455 ;
        RECT 121.190 86.445 122.810 86.455 ;
        RECT 5.840 86.190 6.460 86.375 ;
        RECT 37.440 86.190 38.060 86.375 ;
        RECT 5.840 85.960 38.060 86.190 ;
        RECT 5.840 85.775 6.460 85.960 ;
        RECT 37.440 85.775 38.060 85.960 ;
        RECT 38.290 86.190 38.910 86.375 ;
        RECT 69.890 86.190 70.510 86.375 ;
        RECT 38.290 85.960 70.510 86.190 ;
        RECT 38.290 85.775 38.910 85.960 ;
        RECT 69.890 85.775 70.510 85.960 ;
        RECT 70.740 86.190 71.360 86.375 ;
        RECT 102.340 86.190 102.960 86.375 ;
        RECT 70.740 85.960 102.960 86.190 ;
        RECT 70.740 85.775 71.360 85.960 ;
        RECT 102.340 85.775 102.960 85.960 ;
        RECT 103.190 86.190 103.810 86.375 ;
        RECT 134.790 86.190 135.410 86.375 ;
        RECT 103.190 85.960 135.410 86.190 ;
        RECT 103.190 85.775 103.810 85.960 ;
        RECT 134.790 85.775 135.410 85.960 ;
        RECT 6.690 85.325 37.210 85.705 ;
        RECT 39.140 85.325 69.660 85.705 ;
        RECT 71.590 85.325 102.110 85.705 ;
        RECT 104.040 85.325 134.560 85.705 ;
        RECT 0.960 85.045 3.025 85.275 ;
        RECT 3.255 85.045 4.650 85.275 ;
        RECT 0.130 84.325 1.860 84.555 ;
        RECT 2.160 84.325 3.820 84.555 ;
        RECT 0.130 82.315 0.730 84.325 ;
        RECT 2.160 83.290 2.390 84.325 ;
        RECT 2.795 83.035 3.025 84.080 ;
        RECT 4.050 83.035 4.650 85.045 ;
        RECT 6.690 84.610 37.210 84.980 ;
        RECT 39.140 84.610 69.660 84.980 ;
        RECT 71.590 84.610 102.110 84.980 ;
        RECT 104.040 84.610 134.560 84.980 ;
        RECT 27.680 84.600 29.300 84.610 ;
        RECT 60.130 84.600 61.750 84.610 ;
        RECT 92.580 84.600 94.200 84.610 ;
        RECT 125.030 84.600 126.650 84.610 ;
        RECT 5.840 84.345 6.460 84.530 ;
        RECT 37.440 84.345 38.060 84.530 ;
        RECT 5.840 84.115 38.060 84.345 ;
        RECT 5.840 83.930 6.460 84.115 ;
        RECT 37.440 83.930 38.060 84.115 ;
        RECT 38.290 84.345 38.910 84.530 ;
        RECT 69.890 84.345 70.510 84.530 ;
        RECT 38.290 84.115 70.510 84.345 ;
        RECT 38.290 83.930 38.910 84.115 ;
        RECT 69.890 83.930 70.510 84.115 ;
        RECT 70.740 84.345 71.360 84.530 ;
        RECT 102.340 84.345 102.960 84.530 ;
        RECT 70.740 84.115 102.960 84.345 ;
        RECT 70.740 83.930 71.360 84.115 ;
        RECT 102.340 83.930 102.960 84.115 ;
        RECT 103.190 84.345 103.810 84.530 ;
        RECT 134.790 84.345 135.410 84.530 ;
        RECT 103.190 84.115 135.410 84.345 ;
        RECT 103.190 83.930 103.810 84.115 ;
        RECT 134.790 83.930 135.410 84.115 ;
        RECT 6.690 83.480 37.210 83.860 ;
        RECT 39.140 83.480 69.660 83.860 ;
        RECT 71.590 83.480 102.110 83.860 ;
        RECT 104.040 83.480 134.560 83.860 ;
        RECT 0.960 82.805 3.025 83.035 ;
        RECT 3.255 82.805 4.650 83.035 ;
        RECT 0.130 82.085 1.860 82.315 ;
        RECT 2.160 82.085 3.820 82.315 ;
        RECT 0.130 79.910 0.730 82.085 ;
        RECT 2.160 81.050 2.390 82.085 ;
        RECT 2.795 80.795 3.025 81.840 ;
        RECT 4.050 80.795 4.650 82.805 ;
        RECT 6.700 82.690 37.200 83.130 ;
        RECT 39.150 82.690 69.650 83.130 ;
        RECT 71.600 82.690 102.100 83.130 ;
        RECT 104.050 82.690 134.550 83.130 ;
        RECT 6.690 81.970 37.210 82.340 ;
        RECT 39.140 81.970 69.660 82.340 ;
        RECT 71.590 81.970 102.110 82.340 ;
        RECT 104.040 81.970 134.560 82.340 ;
        RECT 31.520 81.960 33.140 81.970 ;
        RECT 63.970 81.960 65.590 81.970 ;
        RECT 96.420 81.960 98.040 81.970 ;
        RECT 128.870 81.960 130.490 81.970 ;
        RECT 5.840 81.705 6.460 81.890 ;
        RECT 37.440 81.705 38.060 81.890 ;
        RECT 5.840 81.475 38.060 81.705 ;
        RECT 5.840 81.290 6.460 81.475 ;
        RECT 37.440 81.290 38.060 81.475 ;
        RECT 38.290 81.705 38.910 81.890 ;
        RECT 69.890 81.705 70.510 81.890 ;
        RECT 38.290 81.475 70.510 81.705 ;
        RECT 38.290 81.290 38.910 81.475 ;
        RECT 69.890 81.290 70.510 81.475 ;
        RECT 70.740 81.705 71.360 81.890 ;
        RECT 102.340 81.705 102.960 81.890 ;
        RECT 70.740 81.475 102.960 81.705 ;
        RECT 70.740 81.290 71.360 81.475 ;
        RECT 102.340 81.290 102.960 81.475 ;
        RECT 103.190 81.705 103.810 81.890 ;
        RECT 134.790 81.705 135.410 81.890 ;
        RECT 103.190 81.475 135.410 81.705 ;
        RECT 103.190 81.290 103.810 81.475 ;
        RECT 134.790 81.290 135.410 81.475 ;
        RECT 6.690 80.840 37.210 81.220 ;
        RECT 39.140 80.840 69.660 81.220 ;
        RECT 71.590 80.840 102.110 81.220 ;
        RECT 104.040 80.840 134.560 81.220 ;
        RECT 0.960 80.565 3.025 80.795 ;
        RECT 3.255 80.565 4.650 80.795 ;
        RECT 4.050 79.910 4.650 80.565 ;
        RECT 6.690 80.130 37.210 80.500 ;
        RECT 39.140 80.130 69.660 80.500 ;
        RECT 71.590 80.130 102.110 80.500 ;
        RECT 104.040 80.130 134.560 80.500 ;
        RECT 35.360 80.120 36.980 80.130 ;
        RECT 67.810 80.120 69.430 80.130 ;
        RECT 100.260 80.120 101.880 80.130 ;
        RECT 132.710 80.120 134.330 80.130 ;
        RECT 0.130 79.570 2.430 79.910 ;
        RECT 3.160 79.570 4.650 79.910 ;
        RECT 0.130 78.605 0.730 79.570 ;
        RECT 4.050 78.605 4.650 79.570 ;
        RECT 5.840 79.865 6.460 80.050 ;
        RECT 37.440 79.865 38.060 80.050 ;
        RECT 5.840 79.635 38.060 79.865 ;
        RECT 5.840 79.450 6.460 79.635 ;
        RECT 37.440 79.450 38.060 79.635 ;
        RECT 38.290 79.865 38.910 80.050 ;
        RECT 69.890 79.865 70.510 80.050 ;
        RECT 38.290 79.635 70.510 79.865 ;
        RECT 38.290 79.450 38.910 79.635 ;
        RECT 69.890 79.450 70.510 79.635 ;
        RECT 70.740 79.865 71.360 80.050 ;
        RECT 102.340 79.865 102.960 80.050 ;
        RECT 70.740 79.635 102.960 79.865 ;
        RECT 70.740 79.450 71.360 79.635 ;
        RECT 102.340 79.450 102.960 79.635 ;
        RECT 103.190 79.865 103.810 80.050 ;
        RECT 134.790 79.865 135.410 80.050 ;
        RECT 103.190 79.635 135.410 79.865 ;
        RECT 136.340 79.700 136.710 97.630 ;
        RECT 137.360 96.335 137.730 101.955 ;
        RECT 138.380 99.460 138.750 117.970 ;
        RECT 139.400 114.335 139.770 117.970 ;
        RECT 139.395 113.955 139.775 114.335 ;
        RECT 139.400 111.335 139.770 113.955 ;
        RECT 139.395 110.955 139.775 111.335 ;
        RECT 139.400 108.335 139.770 110.955 ;
        RECT 139.395 107.955 139.775 108.335 ;
        RECT 139.400 105.335 139.770 107.955 ;
        RECT 139.395 104.955 139.775 105.335 ;
        RECT 139.400 102.335 139.770 104.955 ;
        RECT 139.395 101.955 139.775 102.335 ;
        RECT 138.380 99.080 138.760 99.460 ;
        RECT 138.380 98.010 138.750 99.080 ;
        RECT 138.380 97.630 138.760 98.010 ;
        RECT 137.355 95.955 137.735 96.335 ;
        RECT 137.360 93.335 137.730 95.955 ;
        RECT 137.355 92.955 137.735 93.335 ;
        RECT 137.360 90.335 137.730 92.955 ;
        RECT 137.355 89.955 137.735 90.335 ;
        RECT 137.360 87.335 137.730 89.955 ;
        RECT 137.355 86.955 137.735 87.335 ;
        RECT 137.360 84.335 137.730 86.955 ;
        RECT 137.355 83.955 137.735 84.335 ;
        RECT 137.360 81.335 137.730 83.955 ;
        RECT 137.355 80.955 137.735 81.335 ;
        RECT 137.360 79.700 137.730 80.955 ;
        RECT 138.380 79.700 138.750 97.630 ;
        RECT 139.400 96.335 139.770 101.955 ;
        RECT 139.395 95.955 139.775 96.335 ;
        RECT 139.400 93.335 139.770 95.955 ;
        RECT 139.395 92.955 139.775 93.335 ;
        RECT 139.400 90.335 139.770 92.955 ;
        RECT 139.395 89.955 139.775 90.335 ;
        RECT 139.400 87.335 139.770 89.955 ;
        RECT 139.395 86.955 139.775 87.335 ;
        RECT 139.400 84.335 139.770 86.955 ;
        RECT 139.395 83.955 139.775 84.335 ;
        RECT 139.400 81.335 139.770 83.955 ;
        RECT 139.395 80.955 139.775 81.335 ;
        RECT 139.400 79.700 139.770 80.955 ;
        RECT 140.420 79.700 140.800 117.970 ;
        RECT 141.150 79.710 141.590 117.960 ;
        RECT 103.190 79.450 103.810 79.635 ;
        RECT 134.790 79.450 135.410 79.635 ;
        RECT 6.690 79.000 37.210 79.380 ;
        RECT 39.140 79.000 69.660 79.380 ;
        RECT 71.590 79.000 102.110 79.380 ;
        RECT 104.040 79.000 134.560 79.380 ;
        RECT 0.130 78.265 2.430 78.605 ;
        RECT 3.160 78.265 4.650 78.605 ;
        RECT 6.690 78.280 37.210 78.660 ;
        RECT 39.140 78.280 69.660 78.660 ;
        RECT 71.590 78.280 102.110 78.660 ;
        RECT 104.040 78.280 134.560 78.660 ;
        RECT 0.130 77.650 0.730 78.265 ;
        RECT 0.130 77.420 1.860 77.650 ;
        RECT 2.160 77.420 3.820 77.650 ;
        RECT 0.130 75.410 0.730 77.420 ;
        RECT 2.160 76.385 2.390 77.420 ;
        RECT 2.795 76.130 3.025 77.175 ;
        RECT 4.050 76.130 4.650 78.265 ;
        RECT 5.840 78.025 6.460 78.210 ;
        RECT 37.440 78.025 38.060 78.210 ;
        RECT 5.840 77.795 38.060 78.025 ;
        RECT 5.840 77.610 6.460 77.795 ;
        RECT 37.440 77.610 38.060 77.795 ;
        RECT 38.290 78.025 38.910 78.210 ;
        RECT 69.890 78.025 70.510 78.210 ;
        RECT 38.290 77.795 70.510 78.025 ;
        RECT 38.290 77.610 38.910 77.795 ;
        RECT 69.890 77.610 70.510 77.795 ;
        RECT 70.740 78.025 71.360 78.210 ;
        RECT 102.340 78.025 102.960 78.210 ;
        RECT 70.740 77.795 102.960 78.025 ;
        RECT 70.740 77.610 71.360 77.795 ;
        RECT 102.340 77.610 102.960 77.795 ;
        RECT 103.190 78.025 103.810 78.210 ;
        RECT 134.790 78.025 135.410 78.210 ;
        RECT 103.190 77.795 135.410 78.025 ;
        RECT 103.190 77.610 103.810 77.795 ;
        RECT 134.790 77.610 135.410 77.795 ;
        RECT 33.440 77.530 35.060 77.540 ;
        RECT 65.890 77.530 67.510 77.540 ;
        RECT 98.340 77.530 99.960 77.540 ;
        RECT 130.790 77.530 132.410 77.540 ;
        RECT 6.690 77.160 37.210 77.530 ;
        RECT 39.140 77.160 69.660 77.530 ;
        RECT 71.590 77.160 102.110 77.530 ;
        RECT 104.040 77.160 134.560 77.530 ;
        RECT 6.690 76.440 37.210 76.820 ;
        RECT 39.140 76.440 69.660 76.820 ;
        RECT 71.590 76.440 102.110 76.820 ;
        RECT 104.040 76.440 134.560 76.820 ;
        RECT 0.960 75.900 3.025 76.130 ;
        RECT 3.255 75.900 4.650 76.130 ;
        RECT 0.130 75.180 1.860 75.410 ;
        RECT 2.160 75.180 3.820 75.410 ;
        RECT 0.130 73.170 0.730 75.180 ;
        RECT 2.160 74.145 2.390 75.180 ;
        RECT 2.795 73.890 3.025 74.935 ;
        RECT 4.050 73.890 4.650 75.900 ;
        RECT 5.840 76.185 6.460 76.370 ;
        RECT 37.440 76.185 38.060 76.370 ;
        RECT 5.840 75.955 38.060 76.185 ;
        RECT 5.840 75.770 6.460 75.955 ;
        RECT 37.440 75.770 38.060 75.955 ;
        RECT 38.290 76.185 38.910 76.370 ;
        RECT 69.890 76.185 70.510 76.370 ;
        RECT 38.290 75.955 70.510 76.185 ;
        RECT 38.290 75.770 38.910 75.955 ;
        RECT 69.890 75.770 70.510 75.955 ;
        RECT 70.740 76.185 71.360 76.370 ;
        RECT 102.340 76.185 102.960 76.370 ;
        RECT 70.740 75.955 102.960 76.185 ;
        RECT 70.740 75.770 71.360 75.955 ;
        RECT 102.340 75.770 102.960 75.955 ;
        RECT 103.190 76.185 103.810 76.370 ;
        RECT 134.790 76.185 135.410 76.370 ;
        RECT 103.190 75.955 135.410 76.185 ;
        RECT 103.190 75.770 103.810 75.955 ;
        RECT 134.790 75.770 135.410 75.955 ;
        RECT 29.600 75.690 31.220 75.700 ;
        RECT 62.050 75.690 63.670 75.700 ;
        RECT 94.500 75.690 96.120 75.700 ;
        RECT 126.950 75.690 128.570 75.700 ;
        RECT 6.690 75.320 37.210 75.690 ;
        RECT 39.140 75.320 69.660 75.690 ;
        RECT 71.590 75.320 102.110 75.690 ;
        RECT 104.040 75.320 134.560 75.690 ;
        RECT 6.700 74.525 37.200 74.965 ;
        RECT 39.150 74.525 69.650 74.965 ;
        RECT 71.600 74.525 102.100 74.965 ;
        RECT 104.050 74.525 134.550 74.965 ;
        RECT 0.960 73.660 3.025 73.890 ;
        RECT 3.255 73.660 4.650 73.890 ;
        RECT 6.690 73.795 37.210 74.175 ;
        RECT 39.140 73.795 69.660 74.175 ;
        RECT 71.590 73.795 102.110 74.175 ;
        RECT 104.040 73.795 134.560 74.175 ;
        RECT 0.130 72.940 1.860 73.170 ;
        RECT 2.160 72.940 3.820 73.170 ;
        RECT 0.130 70.930 0.730 72.940 ;
        RECT 2.160 71.905 2.390 72.940 ;
        RECT 2.795 71.650 3.025 72.695 ;
        RECT 4.050 71.650 4.650 73.660 ;
        RECT 5.840 73.540 6.460 73.725 ;
        RECT 37.440 73.540 38.060 73.725 ;
        RECT 5.840 73.310 38.060 73.540 ;
        RECT 5.840 73.125 6.460 73.310 ;
        RECT 37.440 73.125 38.060 73.310 ;
        RECT 38.290 73.540 38.910 73.725 ;
        RECT 69.890 73.540 70.510 73.725 ;
        RECT 38.290 73.310 70.510 73.540 ;
        RECT 38.290 73.125 38.910 73.310 ;
        RECT 69.890 73.125 70.510 73.310 ;
        RECT 70.740 73.540 71.360 73.725 ;
        RECT 102.340 73.540 102.960 73.725 ;
        RECT 70.740 73.310 102.960 73.540 ;
        RECT 70.740 73.125 71.360 73.310 ;
        RECT 102.340 73.125 102.960 73.310 ;
        RECT 103.190 73.540 103.810 73.725 ;
        RECT 134.790 73.540 135.410 73.725 ;
        RECT 103.190 73.310 135.410 73.540 ;
        RECT 103.190 73.125 103.810 73.310 ;
        RECT 134.790 73.125 135.410 73.310 ;
        RECT 25.760 73.045 27.380 73.055 ;
        RECT 58.210 73.045 59.830 73.055 ;
        RECT 90.660 73.045 92.280 73.055 ;
        RECT 123.110 73.045 124.730 73.055 ;
        RECT 6.690 72.675 37.210 73.045 ;
        RECT 39.140 72.675 69.660 73.045 ;
        RECT 71.590 72.675 102.110 73.045 ;
        RECT 104.040 72.675 134.560 73.045 ;
        RECT 6.690 71.955 37.210 72.335 ;
        RECT 39.140 71.955 69.660 72.335 ;
        RECT 71.590 71.955 102.110 72.335 ;
        RECT 104.040 71.955 134.560 72.335 ;
        RECT 0.960 71.420 3.025 71.650 ;
        RECT 3.255 71.420 4.650 71.650 ;
        RECT 0.130 70.700 1.860 70.930 ;
        RECT 2.160 70.700 3.820 70.930 ;
        RECT 0.130 68.690 0.730 70.700 ;
        RECT 2.160 69.665 2.390 70.700 ;
        RECT 2.795 69.410 3.025 70.455 ;
        RECT 4.050 69.410 4.650 71.420 ;
        RECT 5.840 71.700 6.460 71.885 ;
        RECT 37.440 71.700 38.060 71.885 ;
        RECT 5.840 71.470 38.060 71.700 ;
        RECT 5.840 71.285 6.460 71.470 ;
        RECT 37.440 71.285 38.060 71.470 ;
        RECT 38.290 71.700 38.910 71.885 ;
        RECT 69.890 71.700 70.510 71.885 ;
        RECT 38.290 71.470 70.510 71.700 ;
        RECT 38.290 71.285 38.910 71.470 ;
        RECT 69.890 71.285 70.510 71.470 ;
        RECT 70.740 71.700 71.360 71.885 ;
        RECT 102.340 71.700 102.960 71.885 ;
        RECT 70.740 71.470 102.960 71.700 ;
        RECT 70.740 71.285 71.360 71.470 ;
        RECT 102.340 71.285 102.960 71.470 ;
        RECT 103.190 71.700 103.810 71.885 ;
        RECT 134.790 71.700 135.410 71.885 ;
        RECT 103.190 71.470 135.410 71.700 ;
        RECT 103.190 71.285 103.810 71.470 ;
        RECT 134.790 71.285 135.410 71.470 ;
        RECT 21.920 71.205 23.540 71.215 ;
        RECT 54.370 71.205 55.990 71.215 ;
        RECT 86.820 71.205 88.440 71.215 ;
        RECT 119.270 71.205 120.890 71.215 ;
        RECT 6.690 70.835 37.210 71.205 ;
        RECT 39.140 70.835 69.660 71.205 ;
        RECT 71.590 70.835 102.110 71.205 ;
        RECT 104.040 70.835 134.560 71.205 ;
        RECT 6.690 70.115 37.210 70.495 ;
        RECT 39.140 70.115 69.660 70.495 ;
        RECT 71.590 70.115 102.110 70.495 ;
        RECT 104.040 70.115 134.560 70.495 ;
        RECT 5.840 69.860 6.460 70.045 ;
        RECT 37.440 69.860 38.060 70.045 ;
        RECT 5.840 69.630 38.060 69.860 ;
        RECT 5.840 69.445 6.460 69.630 ;
        RECT 37.440 69.445 38.060 69.630 ;
        RECT 38.290 69.860 38.910 70.045 ;
        RECT 69.890 69.860 70.510 70.045 ;
        RECT 38.290 69.630 70.510 69.860 ;
        RECT 38.290 69.445 38.910 69.630 ;
        RECT 69.890 69.445 70.510 69.630 ;
        RECT 70.740 69.860 71.360 70.045 ;
        RECT 102.340 69.860 102.960 70.045 ;
        RECT 70.740 69.630 102.960 69.860 ;
        RECT 70.740 69.445 71.360 69.630 ;
        RECT 102.340 69.445 102.960 69.630 ;
        RECT 103.190 69.860 103.810 70.045 ;
        RECT 134.790 69.860 135.410 70.045 ;
        RECT 103.190 69.630 135.410 69.860 ;
        RECT 103.190 69.445 103.810 69.630 ;
        RECT 134.790 69.445 135.410 69.630 ;
        RECT 0.960 69.180 3.025 69.410 ;
        RECT 3.255 69.180 4.650 69.410 ;
        RECT 18.080 69.365 19.700 69.375 ;
        RECT 50.530 69.365 52.150 69.375 ;
        RECT 82.980 69.365 84.600 69.375 ;
        RECT 115.430 69.365 117.050 69.375 ;
        RECT 0.130 68.460 1.860 68.690 ;
        RECT 2.160 68.460 3.820 68.690 ;
        RECT 0.130 66.305 0.730 68.460 ;
        RECT 2.160 67.425 2.390 68.460 ;
        RECT 2.795 67.170 3.025 68.215 ;
        RECT 4.050 67.170 4.650 69.180 ;
        RECT 6.690 68.995 37.210 69.365 ;
        RECT 39.140 68.995 69.660 69.365 ;
        RECT 71.590 68.995 102.110 69.365 ;
        RECT 104.040 68.995 134.560 69.365 ;
        RECT 6.700 68.200 37.200 68.640 ;
        RECT 39.150 68.200 69.650 68.640 ;
        RECT 71.600 68.200 102.100 68.640 ;
        RECT 104.050 68.200 134.550 68.640 ;
        RECT 6.690 67.470 37.210 67.850 ;
        RECT 39.140 67.470 69.660 67.850 ;
        RECT 71.590 67.470 102.110 67.850 ;
        RECT 104.040 67.470 134.560 67.850 ;
        RECT 0.960 66.940 3.025 67.170 ;
        RECT 3.255 66.940 4.650 67.170 ;
        RECT 4.050 66.305 4.650 66.940 ;
        RECT 5.840 67.215 6.460 67.400 ;
        RECT 37.440 67.215 38.060 67.400 ;
        RECT 5.840 66.985 38.060 67.215 ;
        RECT 5.840 66.800 6.460 66.985 ;
        RECT 37.440 66.800 38.060 66.985 ;
        RECT 38.290 67.215 38.910 67.400 ;
        RECT 69.890 67.215 70.510 67.400 ;
        RECT 38.290 66.985 70.510 67.215 ;
        RECT 38.290 66.800 38.910 66.985 ;
        RECT 69.890 66.800 70.510 66.985 ;
        RECT 70.740 67.215 71.360 67.400 ;
        RECT 102.340 67.215 102.960 67.400 ;
        RECT 70.740 66.985 102.960 67.215 ;
        RECT 70.740 66.800 71.360 66.985 ;
        RECT 102.340 66.800 102.960 66.985 ;
        RECT 103.190 67.215 103.810 67.400 ;
        RECT 134.790 67.215 135.410 67.400 ;
        RECT 103.190 66.985 135.410 67.215 ;
        RECT 103.190 66.800 103.810 66.985 ;
        RECT 134.790 66.800 135.410 66.985 ;
        RECT 14.240 66.720 15.860 66.730 ;
        RECT 46.690 66.720 48.310 66.730 ;
        RECT 79.140 66.720 80.760 66.730 ;
        RECT 111.590 66.720 113.210 66.730 ;
        RECT 6.690 66.350 37.210 66.720 ;
        RECT 39.140 66.350 69.660 66.720 ;
        RECT 71.590 66.350 102.110 66.720 ;
        RECT 104.040 66.350 134.560 66.720 ;
        RECT 0.130 65.965 2.420 66.305 ;
        RECT 3.165 65.965 4.650 66.305 ;
        RECT 0.130 65.330 0.730 65.965 ;
        RECT 0.130 65.100 1.860 65.330 ;
        RECT 2.160 65.100 3.820 65.330 ;
        RECT 0.130 63.090 0.730 65.100 ;
        RECT 2.160 64.065 2.390 65.100 ;
        RECT 2.795 63.810 3.025 64.855 ;
        RECT 4.050 63.810 4.650 65.965 ;
        RECT 6.690 65.630 37.210 66.010 ;
        RECT 39.140 65.630 69.660 66.010 ;
        RECT 71.590 65.630 102.110 66.010 ;
        RECT 104.040 65.630 134.560 66.010 ;
        RECT 5.840 65.375 6.460 65.560 ;
        RECT 37.440 65.375 38.060 65.560 ;
        RECT 5.840 65.145 38.060 65.375 ;
        RECT 5.840 64.960 6.460 65.145 ;
        RECT 37.440 64.960 38.060 65.145 ;
        RECT 38.290 65.375 38.910 65.560 ;
        RECT 69.890 65.375 70.510 65.560 ;
        RECT 38.290 65.145 70.510 65.375 ;
        RECT 38.290 64.960 38.910 65.145 ;
        RECT 69.890 64.960 70.510 65.145 ;
        RECT 70.740 65.375 71.360 65.560 ;
        RECT 102.340 65.375 102.960 65.560 ;
        RECT 70.740 65.145 102.960 65.375 ;
        RECT 70.740 64.960 71.360 65.145 ;
        RECT 102.340 64.960 102.960 65.145 ;
        RECT 103.190 65.375 103.810 65.560 ;
        RECT 134.790 65.375 135.410 65.560 ;
        RECT 103.190 65.145 135.410 65.375 ;
        RECT 103.190 64.960 103.810 65.145 ;
        RECT 134.790 64.960 135.410 65.145 ;
        RECT 10.400 64.880 12.020 64.890 ;
        RECT 42.850 64.880 44.470 64.890 ;
        RECT 75.300 64.880 76.920 64.890 ;
        RECT 107.750 64.880 109.370 64.890 ;
        RECT 6.690 64.510 37.210 64.880 ;
        RECT 39.140 64.510 69.660 64.880 ;
        RECT 71.590 64.510 102.110 64.880 ;
        RECT 104.040 64.510 134.560 64.880 ;
        RECT 0.960 63.580 3.025 63.810 ;
        RECT 3.255 63.580 4.650 63.810 ;
        RECT 6.690 63.790 37.210 64.170 ;
        RECT 39.140 63.790 69.660 64.170 ;
        RECT 71.590 63.790 102.110 64.170 ;
        RECT 104.040 63.790 134.560 64.170 ;
        RECT 0.130 62.860 1.860 63.090 ;
        RECT 2.160 62.860 3.820 63.090 ;
        RECT 0.130 60.705 0.730 62.860 ;
        RECT 2.160 61.825 2.390 62.860 ;
        RECT 2.795 61.570 3.025 62.615 ;
        RECT 4.050 61.570 4.650 63.580 ;
        RECT 5.840 63.535 6.460 63.720 ;
        RECT 37.440 63.535 38.060 63.720 ;
        RECT 5.840 63.305 38.060 63.535 ;
        RECT 5.840 63.120 6.460 63.305 ;
        RECT 37.440 63.120 38.060 63.305 ;
        RECT 38.290 63.535 38.910 63.720 ;
        RECT 69.890 63.535 70.510 63.720 ;
        RECT 38.290 63.305 70.510 63.535 ;
        RECT 38.290 63.120 38.910 63.305 ;
        RECT 69.890 63.120 70.510 63.305 ;
        RECT 70.740 63.535 71.360 63.720 ;
        RECT 102.340 63.535 102.960 63.720 ;
        RECT 70.740 63.305 102.960 63.535 ;
        RECT 70.740 63.120 71.360 63.305 ;
        RECT 102.340 63.120 102.960 63.305 ;
        RECT 103.190 63.535 103.810 63.720 ;
        RECT 134.790 63.535 135.410 63.720 ;
        RECT 103.190 63.305 135.410 63.535 ;
        RECT 103.190 63.120 103.810 63.305 ;
        RECT 134.790 63.120 135.410 63.305 ;
        RECT 6.690 62.670 37.210 63.040 ;
        RECT 39.140 62.670 69.660 63.040 ;
        RECT 71.590 62.670 102.110 63.040 ;
        RECT 104.040 62.670 134.560 63.040 ;
        RECT 0.960 61.340 3.025 61.570 ;
        RECT 3.255 61.340 4.650 61.570 ;
        RECT 4.050 60.705 4.650 61.340 ;
        RECT 0.130 60.365 2.420 60.705 ;
        RECT 3.165 60.365 4.650 60.705 ;
        RECT 0.130 59.730 0.730 60.365 ;
        RECT 0.130 59.500 1.710 59.730 ;
        RECT 0.130 57.460 0.730 59.500 ;
        RECT 2.140 59.270 2.500 59.355 ;
        RECT 1.010 59.040 2.500 59.270 ;
        RECT 1.010 58.890 1.370 59.040 ;
        RECT 0.960 58.255 1.910 58.660 ;
        RECT 0.130 57.230 1.420 57.460 ;
        RECT 0.130 56.270 0.730 57.230 ;
        RECT 1.650 56.910 1.910 58.255 ;
        RECT 2.140 57.605 2.500 59.040 ;
        RECT 2.730 57.705 3.080 58.905 ;
        RECT 3.440 58.295 3.820 59.940 ;
        RECT 2.520 56.910 2.870 56.970 ;
        RECT 3.440 56.910 3.780 57.515 ;
        RECT 1.650 56.650 3.780 56.910 ;
        RECT 2.520 56.590 2.870 56.650 ;
        RECT 4.050 56.370 4.650 60.365 ;
        RECT 6.495 59.885 8.245 62.670 ;
        RECT 8.885 59.885 9.695 60.885 ;
        RECT 10.335 59.885 12.085 62.180 ;
        RECT 12.725 59.885 13.535 60.885 ;
        RECT 14.175 59.885 15.925 62.180 ;
        RECT 16.565 59.885 17.375 60.885 ;
        RECT 18.015 59.885 19.765 62.180 ;
        RECT 20.405 59.885 21.215 60.885 ;
        RECT 21.855 59.885 23.605 62.180 ;
        RECT 24.245 59.885 25.055 60.885 ;
        RECT 25.695 59.885 27.445 62.180 ;
        RECT 28.085 59.885 28.895 60.885 ;
        RECT 29.535 59.885 31.285 62.180 ;
        RECT 31.925 59.885 32.735 60.885 ;
        RECT 33.375 59.885 35.125 62.180 ;
        RECT 35.765 59.885 36.575 60.885 ;
        RECT 38.945 59.885 40.695 62.670 ;
        RECT 41.335 59.885 42.145 60.885 ;
        RECT 42.785 59.885 44.535 62.180 ;
        RECT 45.175 59.885 45.985 60.885 ;
        RECT 46.625 59.885 48.375 62.180 ;
        RECT 49.015 59.885 49.825 60.885 ;
        RECT 50.465 59.885 52.215 62.180 ;
        RECT 52.855 59.885 53.665 60.885 ;
        RECT 54.305 59.885 56.055 62.180 ;
        RECT 56.695 59.885 57.505 60.885 ;
        RECT 58.145 59.885 59.895 62.180 ;
        RECT 60.535 59.885 61.345 60.885 ;
        RECT 61.985 59.885 63.735 62.180 ;
        RECT 64.375 59.885 65.185 60.885 ;
        RECT 65.825 59.885 67.575 62.180 ;
        RECT 68.215 59.885 69.025 60.885 ;
        RECT 71.395 59.885 73.145 62.670 ;
        RECT 73.785 59.885 74.595 60.885 ;
        RECT 75.235 59.885 76.985 62.180 ;
        RECT 77.625 59.885 78.435 60.885 ;
        RECT 79.075 59.885 80.825 62.180 ;
        RECT 81.465 59.885 82.275 60.885 ;
        RECT 82.915 59.885 84.665 62.180 ;
        RECT 85.305 59.885 86.115 60.885 ;
        RECT 86.755 59.885 88.505 62.180 ;
        RECT 89.145 59.885 89.955 60.885 ;
        RECT 90.595 59.885 92.345 62.180 ;
        RECT 92.985 59.885 93.795 60.885 ;
        RECT 94.435 59.885 96.185 62.180 ;
        RECT 96.825 59.885 97.635 60.885 ;
        RECT 98.275 59.885 100.025 62.180 ;
        RECT 100.665 59.885 101.475 60.885 ;
        RECT 103.845 59.885 105.595 62.670 ;
        RECT 106.235 59.885 107.045 60.885 ;
        RECT 107.685 59.885 109.435 62.180 ;
        RECT 110.075 59.885 110.885 60.885 ;
        RECT 111.525 59.885 113.275 62.180 ;
        RECT 113.915 59.885 114.725 60.885 ;
        RECT 115.365 59.885 117.115 62.180 ;
        RECT 117.755 59.885 118.565 60.885 ;
        RECT 119.205 59.885 120.955 62.180 ;
        RECT 121.595 59.885 122.405 60.885 ;
        RECT 123.045 59.885 124.795 62.180 ;
        RECT 125.435 59.885 126.245 60.885 ;
        RECT 126.885 59.885 128.635 62.180 ;
        RECT 129.275 59.885 130.085 60.885 ;
        RECT 130.725 59.885 132.475 62.180 ;
        RECT 133.115 59.885 133.925 60.885 ;
        RECT 136.340 60.075 136.710 78.585 ;
        RECT 137.360 74.950 137.730 78.585 ;
        RECT 137.355 74.570 137.735 74.950 ;
        RECT 137.360 71.950 137.730 74.570 ;
        RECT 137.355 71.570 137.735 71.950 ;
        RECT 137.360 68.950 137.730 71.570 ;
        RECT 137.355 68.570 137.735 68.950 ;
        RECT 137.360 65.950 137.730 68.570 ;
        RECT 137.355 65.570 137.735 65.950 ;
        RECT 137.360 62.950 137.730 65.570 ;
        RECT 137.355 62.570 137.735 62.950 ;
        RECT 136.340 59.695 136.720 60.075 ;
        RECT 136.340 58.625 136.710 59.695 ;
        RECT 6.965 57.435 7.775 58.435 ;
        RECT 0.130 56.040 1.820 56.270 ;
        RECT 3.190 56.140 4.650 56.370 ;
        RECT 0.130 54.030 0.730 56.040 ;
        RECT 2.150 55.580 3.150 55.905 ;
        RECT 0.960 55.020 3.820 55.350 ;
        RECT 0.130 53.800 1.820 54.030 ;
        RECT 0.130 51.790 0.730 53.800 ;
        RECT 2.535 53.665 2.800 55.020 ;
        RECT 4.050 54.130 4.650 56.140 ;
        RECT 8.415 55.605 10.165 58.435 ;
        RECT 10.805 57.435 11.615 58.435 ;
        RECT 12.255 56.140 14.005 58.435 ;
        RECT 14.645 57.435 15.455 58.435 ;
        RECT 16.095 56.140 17.845 58.435 ;
        RECT 18.485 57.435 19.295 58.435 ;
        RECT 19.935 56.140 21.685 58.435 ;
        RECT 22.325 57.435 23.135 58.435 ;
        RECT 23.775 56.140 25.525 58.435 ;
        RECT 26.165 57.435 26.975 58.435 ;
        RECT 27.615 56.140 29.365 58.435 ;
        RECT 30.005 57.435 30.815 58.435 ;
        RECT 31.455 56.140 33.205 58.435 ;
        RECT 33.845 57.435 34.655 58.435 ;
        RECT 35.295 56.140 37.045 58.435 ;
        RECT 39.415 57.435 40.225 58.435 ;
        RECT 40.865 55.605 42.615 58.435 ;
        RECT 43.255 57.435 44.065 58.435 ;
        RECT 44.705 56.140 46.455 58.435 ;
        RECT 47.095 57.435 47.905 58.435 ;
        RECT 48.545 56.140 50.295 58.435 ;
        RECT 50.935 57.435 51.745 58.435 ;
        RECT 52.385 56.140 54.135 58.435 ;
        RECT 54.775 57.435 55.585 58.435 ;
        RECT 56.225 56.140 57.975 58.435 ;
        RECT 58.615 57.435 59.425 58.435 ;
        RECT 60.065 56.140 61.815 58.435 ;
        RECT 62.455 57.435 63.265 58.435 ;
        RECT 63.905 56.140 65.655 58.435 ;
        RECT 66.295 57.435 67.105 58.435 ;
        RECT 67.745 56.140 69.495 58.435 ;
        RECT 71.865 57.435 72.675 58.435 ;
        RECT 73.315 55.605 75.065 58.435 ;
        RECT 75.705 57.435 76.515 58.435 ;
        RECT 77.155 56.140 78.905 58.435 ;
        RECT 79.545 57.435 80.355 58.435 ;
        RECT 80.995 56.140 82.745 58.435 ;
        RECT 83.385 57.435 84.195 58.435 ;
        RECT 84.835 56.140 86.585 58.435 ;
        RECT 87.225 57.435 88.035 58.435 ;
        RECT 88.675 56.140 90.425 58.435 ;
        RECT 91.065 57.435 91.875 58.435 ;
        RECT 92.515 56.140 94.265 58.435 ;
        RECT 94.905 57.435 95.715 58.435 ;
        RECT 96.355 56.140 98.105 58.435 ;
        RECT 98.745 57.435 99.555 58.435 ;
        RECT 100.195 56.140 101.945 58.435 ;
        RECT 104.315 57.435 105.125 58.435 ;
        RECT 105.765 55.605 107.515 58.435 ;
        RECT 108.155 57.435 108.965 58.435 ;
        RECT 109.605 56.140 111.355 58.435 ;
        RECT 111.995 57.435 112.805 58.435 ;
        RECT 113.445 56.140 115.195 58.435 ;
        RECT 115.835 57.435 116.645 58.435 ;
        RECT 117.285 56.140 119.035 58.435 ;
        RECT 119.675 57.435 120.485 58.435 ;
        RECT 121.125 56.140 122.875 58.435 ;
        RECT 123.515 57.435 124.325 58.435 ;
        RECT 124.965 56.140 126.715 58.435 ;
        RECT 127.355 57.435 128.165 58.435 ;
        RECT 128.805 56.140 130.555 58.435 ;
        RECT 131.195 57.435 132.005 58.435 ;
        RECT 132.645 56.140 134.395 58.435 ;
        RECT 136.340 58.245 136.720 58.625 ;
        RECT 6.690 55.235 37.210 55.605 ;
        RECT 39.140 55.235 69.660 55.605 ;
        RECT 71.590 55.235 102.110 55.605 ;
        RECT 104.040 55.235 134.560 55.605 ;
        RECT 5.840 54.970 6.460 55.155 ;
        RECT 37.440 54.970 38.060 55.155 ;
        RECT 5.840 54.740 38.060 54.970 ;
        RECT 5.840 54.555 6.460 54.740 ;
        RECT 37.440 54.555 38.060 54.740 ;
        RECT 38.290 54.970 38.910 55.155 ;
        RECT 69.890 54.970 70.510 55.155 ;
        RECT 38.290 54.740 70.510 54.970 ;
        RECT 38.290 54.555 38.910 54.740 ;
        RECT 69.890 54.555 70.510 54.740 ;
        RECT 70.740 54.970 71.360 55.155 ;
        RECT 102.340 54.970 102.960 55.155 ;
        RECT 70.740 54.740 102.960 54.970 ;
        RECT 70.740 54.555 71.360 54.740 ;
        RECT 102.340 54.555 102.960 54.740 ;
        RECT 103.190 54.970 103.810 55.155 ;
        RECT 134.790 54.970 135.410 55.155 ;
        RECT 103.190 54.740 135.410 54.970 ;
        RECT 103.190 54.555 103.810 54.740 ;
        RECT 134.790 54.555 135.410 54.740 ;
        RECT 3.190 53.900 4.650 54.130 ;
        RECT 6.690 54.105 37.210 54.485 ;
        RECT 39.140 54.105 69.660 54.485 ;
        RECT 71.590 54.105 102.110 54.485 ;
        RECT 104.040 54.105 134.560 54.485 ;
        RECT 2.150 53.340 3.150 53.665 ;
        RECT 0.960 52.780 3.820 53.110 ;
        RECT 4.050 51.890 4.650 53.900 ;
        RECT 6.690 53.395 37.210 53.765 ;
        RECT 39.140 53.395 69.660 53.765 ;
        RECT 71.590 53.395 102.110 53.765 ;
        RECT 104.040 53.395 134.560 53.765 ;
        RECT 12.320 53.385 13.940 53.395 ;
        RECT 44.770 53.385 46.390 53.395 ;
        RECT 77.220 53.385 78.840 53.395 ;
        RECT 109.670 53.385 111.290 53.395 ;
        RECT 5.840 53.130 6.460 53.315 ;
        RECT 37.440 53.130 38.060 53.315 ;
        RECT 5.840 52.900 38.060 53.130 ;
        RECT 5.840 52.715 6.460 52.900 ;
        RECT 37.440 52.715 38.060 52.900 ;
        RECT 38.290 53.130 38.910 53.315 ;
        RECT 69.890 53.130 70.510 53.315 ;
        RECT 38.290 52.900 70.510 53.130 ;
        RECT 38.290 52.715 38.910 52.900 ;
        RECT 69.890 52.715 70.510 52.900 ;
        RECT 70.740 53.130 71.360 53.315 ;
        RECT 102.340 53.130 102.960 53.315 ;
        RECT 70.740 52.900 102.960 53.130 ;
        RECT 70.740 52.715 71.360 52.900 ;
        RECT 102.340 52.715 102.960 52.900 ;
        RECT 103.190 53.130 103.810 53.315 ;
        RECT 134.790 53.130 135.410 53.315 ;
        RECT 103.190 52.900 135.410 53.130 ;
        RECT 103.190 52.715 103.810 52.900 ;
        RECT 134.790 52.715 135.410 52.900 ;
        RECT 6.690 52.265 37.210 52.645 ;
        RECT 39.140 52.265 69.660 52.645 ;
        RECT 71.590 52.265 102.110 52.645 ;
        RECT 104.040 52.265 134.560 52.645 ;
        RECT 0.130 51.560 1.820 51.790 ;
        RECT 3.190 51.660 4.650 51.890 ;
        RECT 0.130 49.505 0.730 51.560 ;
        RECT 2.150 51.100 3.150 51.425 ;
        RECT 0.960 50.540 3.820 50.870 ;
        RECT 2.300 50.415 2.680 50.540 ;
        RECT 4.050 49.505 4.650 51.660 ;
        RECT 6.690 51.550 37.210 51.920 ;
        RECT 39.140 51.550 69.660 51.920 ;
        RECT 71.590 51.550 102.110 51.920 ;
        RECT 104.040 51.550 134.560 51.920 ;
        RECT 16.160 51.540 17.780 51.550 ;
        RECT 48.610 51.540 50.230 51.550 ;
        RECT 81.060 51.540 82.680 51.550 ;
        RECT 113.510 51.540 115.130 51.550 ;
        RECT 5.840 51.285 6.460 51.470 ;
        RECT 37.440 51.285 38.060 51.470 ;
        RECT 5.840 51.055 38.060 51.285 ;
        RECT 5.840 50.870 6.460 51.055 ;
        RECT 37.440 50.870 38.060 51.055 ;
        RECT 38.290 51.285 38.910 51.470 ;
        RECT 69.890 51.285 70.510 51.470 ;
        RECT 38.290 51.055 70.510 51.285 ;
        RECT 38.290 50.870 38.910 51.055 ;
        RECT 69.890 50.870 70.510 51.055 ;
        RECT 70.740 51.285 71.360 51.470 ;
        RECT 102.340 51.285 102.960 51.470 ;
        RECT 70.740 51.055 102.960 51.285 ;
        RECT 70.740 50.870 71.360 51.055 ;
        RECT 102.340 50.870 102.960 51.055 ;
        RECT 103.190 51.285 103.810 51.470 ;
        RECT 134.790 51.285 135.410 51.470 ;
        RECT 103.190 51.055 135.410 51.285 ;
        RECT 103.190 50.870 103.810 51.055 ;
        RECT 134.790 50.870 135.410 51.055 ;
        RECT 6.690 50.420 37.210 50.800 ;
        RECT 39.140 50.420 69.660 50.800 ;
        RECT 71.590 50.420 102.110 50.800 ;
        RECT 104.040 50.420 134.560 50.800 ;
        RECT 6.700 49.630 37.200 50.070 ;
        RECT 39.150 49.630 69.650 50.070 ;
        RECT 71.600 49.630 102.100 50.070 ;
        RECT 104.050 49.630 134.550 50.070 ;
        RECT 0.130 49.165 2.420 49.505 ;
        RECT 3.165 49.165 4.650 49.505 ;
        RECT 0.130 48.385 0.730 49.165 ;
        RECT 4.050 48.385 4.650 49.165 ;
        RECT 6.690 48.910 37.210 49.280 ;
        RECT 39.140 48.910 69.660 49.280 ;
        RECT 71.590 48.910 102.110 49.280 ;
        RECT 104.040 48.910 134.560 49.280 ;
        RECT 20.000 48.900 21.620 48.910 ;
        RECT 52.450 48.900 54.070 48.910 ;
        RECT 84.900 48.900 86.520 48.910 ;
        RECT 117.350 48.900 118.970 48.910 ;
        RECT 0.130 48.045 2.420 48.385 ;
        RECT 3.165 48.045 4.650 48.385 ;
        RECT 5.840 48.645 6.460 48.830 ;
        RECT 37.440 48.645 38.060 48.830 ;
        RECT 5.840 48.415 38.060 48.645 ;
        RECT 5.840 48.230 6.460 48.415 ;
        RECT 37.440 48.230 38.060 48.415 ;
        RECT 38.290 48.645 38.910 48.830 ;
        RECT 69.890 48.645 70.510 48.830 ;
        RECT 38.290 48.415 70.510 48.645 ;
        RECT 38.290 48.230 38.910 48.415 ;
        RECT 69.890 48.230 70.510 48.415 ;
        RECT 70.740 48.645 71.360 48.830 ;
        RECT 102.340 48.645 102.960 48.830 ;
        RECT 70.740 48.415 102.960 48.645 ;
        RECT 70.740 48.230 71.360 48.415 ;
        RECT 102.340 48.230 102.960 48.415 ;
        RECT 103.190 48.645 103.810 48.830 ;
        RECT 134.790 48.645 135.410 48.830 ;
        RECT 103.190 48.415 135.410 48.645 ;
        RECT 103.190 48.230 103.810 48.415 ;
        RECT 134.790 48.230 135.410 48.415 ;
        RECT 0.130 47.410 0.730 48.045 ;
        RECT 0.130 47.180 1.860 47.410 ;
        RECT 2.160 47.180 3.820 47.410 ;
        RECT 0.130 45.170 0.730 47.180 ;
        RECT 2.160 46.145 2.390 47.180 ;
        RECT 2.795 45.890 3.025 46.935 ;
        RECT 4.050 45.890 4.650 48.045 ;
        RECT 6.690 47.780 37.210 48.160 ;
        RECT 39.140 47.780 69.660 48.160 ;
        RECT 71.590 47.780 102.110 48.160 ;
        RECT 104.040 47.780 134.560 48.160 ;
        RECT 6.690 47.070 37.210 47.440 ;
        RECT 39.140 47.070 69.660 47.440 ;
        RECT 71.590 47.070 102.110 47.440 ;
        RECT 104.040 47.070 134.560 47.440 ;
        RECT 23.840 47.060 25.460 47.070 ;
        RECT 56.290 47.060 57.910 47.070 ;
        RECT 88.740 47.060 90.360 47.070 ;
        RECT 121.190 47.060 122.810 47.070 ;
        RECT 5.840 46.805 6.460 46.990 ;
        RECT 37.440 46.805 38.060 46.990 ;
        RECT 5.840 46.575 38.060 46.805 ;
        RECT 5.840 46.390 6.460 46.575 ;
        RECT 37.440 46.390 38.060 46.575 ;
        RECT 38.290 46.805 38.910 46.990 ;
        RECT 69.890 46.805 70.510 46.990 ;
        RECT 38.290 46.575 70.510 46.805 ;
        RECT 38.290 46.390 38.910 46.575 ;
        RECT 69.890 46.390 70.510 46.575 ;
        RECT 70.740 46.805 71.360 46.990 ;
        RECT 102.340 46.805 102.960 46.990 ;
        RECT 70.740 46.575 102.960 46.805 ;
        RECT 70.740 46.390 71.360 46.575 ;
        RECT 102.340 46.390 102.960 46.575 ;
        RECT 103.190 46.805 103.810 46.990 ;
        RECT 134.790 46.805 135.410 46.990 ;
        RECT 103.190 46.575 135.410 46.805 ;
        RECT 103.190 46.390 103.810 46.575 ;
        RECT 134.790 46.390 135.410 46.575 ;
        RECT 6.690 45.940 37.210 46.320 ;
        RECT 39.140 45.940 69.660 46.320 ;
        RECT 71.590 45.940 102.110 46.320 ;
        RECT 104.040 45.940 134.560 46.320 ;
        RECT 0.960 45.660 3.025 45.890 ;
        RECT 3.255 45.660 4.650 45.890 ;
        RECT 0.130 44.940 1.860 45.170 ;
        RECT 2.160 44.940 3.820 45.170 ;
        RECT 0.130 42.930 0.730 44.940 ;
        RECT 2.160 43.905 2.390 44.940 ;
        RECT 2.795 43.650 3.025 44.695 ;
        RECT 4.050 43.650 4.650 45.660 ;
        RECT 6.690 45.225 37.210 45.595 ;
        RECT 39.140 45.225 69.660 45.595 ;
        RECT 71.590 45.225 102.110 45.595 ;
        RECT 104.040 45.225 134.560 45.595 ;
        RECT 27.680 45.215 29.300 45.225 ;
        RECT 60.130 45.215 61.750 45.225 ;
        RECT 92.580 45.215 94.200 45.225 ;
        RECT 125.030 45.215 126.650 45.225 ;
        RECT 5.840 44.960 6.460 45.145 ;
        RECT 37.440 44.960 38.060 45.145 ;
        RECT 5.840 44.730 38.060 44.960 ;
        RECT 5.840 44.545 6.460 44.730 ;
        RECT 37.440 44.545 38.060 44.730 ;
        RECT 38.290 44.960 38.910 45.145 ;
        RECT 69.890 44.960 70.510 45.145 ;
        RECT 38.290 44.730 70.510 44.960 ;
        RECT 38.290 44.545 38.910 44.730 ;
        RECT 69.890 44.545 70.510 44.730 ;
        RECT 70.740 44.960 71.360 45.145 ;
        RECT 102.340 44.960 102.960 45.145 ;
        RECT 70.740 44.730 102.960 44.960 ;
        RECT 70.740 44.545 71.360 44.730 ;
        RECT 102.340 44.545 102.960 44.730 ;
        RECT 103.190 44.960 103.810 45.145 ;
        RECT 134.790 44.960 135.410 45.145 ;
        RECT 103.190 44.730 135.410 44.960 ;
        RECT 103.190 44.545 103.810 44.730 ;
        RECT 134.790 44.545 135.410 44.730 ;
        RECT 6.690 44.095 37.210 44.475 ;
        RECT 39.140 44.095 69.660 44.475 ;
        RECT 71.590 44.095 102.110 44.475 ;
        RECT 104.040 44.095 134.560 44.475 ;
        RECT 0.960 43.420 3.025 43.650 ;
        RECT 3.255 43.420 4.650 43.650 ;
        RECT 0.130 42.700 1.860 42.930 ;
        RECT 2.160 42.700 3.820 42.930 ;
        RECT 0.130 40.525 0.730 42.700 ;
        RECT 2.160 41.665 2.390 42.700 ;
        RECT 2.795 41.410 3.025 42.455 ;
        RECT 4.050 41.410 4.650 43.420 ;
        RECT 6.700 43.305 37.200 43.745 ;
        RECT 39.150 43.305 69.650 43.745 ;
        RECT 71.600 43.305 102.100 43.745 ;
        RECT 104.050 43.305 134.550 43.745 ;
        RECT 6.690 42.585 37.210 42.955 ;
        RECT 39.140 42.585 69.660 42.955 ;
        RECT 71.590 42.585 102.110 42.955 ;
        RECT 104.040 42.585 134.560 42.955 ;
        RECT 31.520 42.575 33.140 42.585 ;
        RECT 63.970 42.575 65.590 42.585 ;
        RECT 96.420 42.575 98.040 42.585 ;
        RECT 128.870 42.575 130.490 42.585 ;
        RECT 5.840 42.320 6.460 42.505 ;
        RECT 37.440 42.320 38.060 42.505 ;
        RECT 5.840 42.090 38.060 42.320 ;
        RECT 5.840 41.905 6.460 42.090 ;
        RECT 37.440 41.905 38.060 42.090 ;
        RECT 38.290 42.320 38.910 42.505 ;
        RECT 69.890 42.320 70.510 42.505 ;
        RECT 38.290 42.090 70.510 42.320 ;
        RECT 38.290 41.905 38.910 42.090 ;
        RECT 69.890 41.905 70.510 42.090 ;
        RECT 70.740 42.320 71.360 42.505 ;
        RECT 102.340 42.320 102.960 42.505 ;
        RECT 70.740 42.090 102.960 42.320 ;
        RECT 70.740 41.905 71.360 42.090 ;
        RECT 102.340 41.905 102.960 42.090 ;
        RECT 103.190 42.320 103.810 42.505 ;
        RECT 134.790 42.320 135.410 42.505 ;
        RECT 103.190 42.090 135.410 42.320 ;
        RECT 103.190 41.905 103.810 42.090 ;
        RECT 134.790 41.905 135.410 42.090 ;
        RECT 6.690 41.455 37.210 41.835 ;
        RECT 39.140 41.455 69.660 41.835 ;
        RECT 71.590 41.455 102.110 41.835 ;
        RECT 104.040 41.455 134.560 41.835 ;
        RECT 0.960 41.180 3.025 41.410 ;
        RECT 3.255 41.180 4.650 41.410 ;
        RECT 4.050 40.525 4.650 41.180 ;
        RECT 6.690 40.745 37.210 41.115 ;
        RECT 39.140 40.745 69.660 41.115 ;
        RECT 71.590 40.745 102.110 41.115 ;
        RECT 104.040 40.745 134.560 41.115 ;
        RECT 35.360 40.735 36.980 40.745 ;
        RECT 67.810 40.735 69.430 40.745 ;
        RECT 100.260 40.735 101.880 40.745 ;
        RECT 132.710 40.735 134.330 40.745 ;
        RECT 0.130 40.185 2.430 40.525 ;
        RECT 3.160 40.185 4.650 40.525 ;
        RECT 0.130 39.220 0.730 40.185 ;
        RECT 4.050 39.220 4.650 40.185 ;
        RECT 5.840 40.480 6.460 40.665 ;
        RECT 37.440 40.480 38.060 40.665 ;
        RECT 5.840 40.250 38.060 40.480 ;
        RECT 5.840 40.065 6.460 40.250 ;
        RECT 37.440 40.065 38.060 40.250 ;
        RECT 38.290 40.480 38.910 40.665 ;
        RECT 69.890 40.480 70.510 40.665 ;
        RECT 38.290 40.250 70.510 40.480 ;
        RECT 38.290 40.065 38.910 40.250 ;
        RECT 69.890 40.065 70.510 40.250 ;
        RECT 70.740 40.480 71.360 40.665 ;
        RECT 102.340 40.480 102.960 40.665 ;
        RECT 70.740 40.250 102.960 40.480 ;
        RECT 70.740 40.065 71.360 40.250 ;
        RECT 102.340 40.065 102.960 40.250 ;
        RECT 103.190 40.480 103.810 40.665 ;
        RECT 134.790 40.480 135.410 40.665 ;
        RECT 103.190 40.250 135.410 40.480 ;
        RECT 136.340 40.315 136.710 58.245 ;
        RECT 137.360 56.950 137.730 62.570 ;
        RECT 138.380 60.075 138.750 78.585 ;
        RECT 139.400 74.950 139.770 78.585 ;
        RECT 139.395 74.570 139.775 74.950 ;
        RECT 139.400 71.950 139.770 74.570 ;
        RECT 139.395 71.570 139.775 71.950 ;
        RECT 139.400 68.950 139.770 71.570 ;
        RECT 139.395 68.570 139.775 68.950 ;
        RECT 139.400 65.950 139.770 68.570 ;
        RECT 139.395 65.570 139.775 65.950 ;
        RECT 139.400 62.950 139.770 65.570 ;
        RECT 139.395 62.570 139.775 62.950 ;
        RECT 138.380 59.695 138.760 60.075 ;
        RECT 138.380 58.625 138.750 59.695 ;
        RECT 138.380 58.245 138.760 58.625 ;
        RECT 137.355 56.570 137.735 56.950 ;
        RECT 137.360 53.950 137.730 56.570 ;
        RECT 137.355 53.570 137.735 53.950 ;
        RECT 137.360 50.950 137.730 53.570 ;
        RECT 137.355 50.570 137.735 50.950 ;
        RECT 137.360 47.950 137.730 50.570 ;
        RECT 137.355 47.570 137.735 47.950 ;
        RECT 137.360 44.950 137.730 47.570 ;
        RECT 137.355 44.570 137.735 44.950 ;
        RECT 137.360 41.950 137.730 44.570 ;
        RECT 137.355 41.570 137.735 41.950 ;
        RECT 137.360 40.315 137.730 41.570 ;
        RECT 138.380 40.315 138.750 58.245 ;
        RECT 139.400 56.950 139.770 62.570 ;
        RECT 139.395 56.570 139.775 56.950 ;
        RECT 139.400 53.950 139.770 56.570 ;
        RECT 139.395 53.570 139.775 53.950 ;
        RECT 139.400 50.950 139.770 53.570 ;
        RECT 139.395 50.570 139.775 50.950 ;
        RECT 139.400 47.950 139.770 50.570 ;
        RECT 139.395 47.570 139.775 47.950 ;
        RECT 139.400 44.950 139.770 47.570 ;
        RECT 139.395 44.570 139.775 44.950 ;
        RECT 139.400 41.950 139.770 44.570 ;
        RECT 139.395 41.570 139.775 41.950 ;
        RECT 139.400 40.315 139.770 41.570 ;
        RECT 140.420 40.315 140.800 78.585 ;
        RECT 141.150 40.325 141.590 78.575 ;
        RECT 103.190 40.065 103.810 40.250 ;
        RECT 134.790 40.065 135.410 40.250 ;
        RECT 6.690 39.615 37.210 39.995 ;
        RECT 39.140 39.615 69.660 39.995 ;
        RECT 71.590 39.615 102.110 39.995 ;
        RECT 104.040 39.615 134.560 39.995 ;
        RECT 0.130 38.880 2.430 39.220 ;
        RECT 3.160 38.880 4.650 39.220 ;
        RECT 6.690 38.895 37.210 39.275 ;
        RECT 39.140 38.895 69.660 39.275 ;
        RECT 71.590 38.895 102.110 39.275 ;
        RECT 104.040 38.895 134.560 39.275 ;
        RECT 0.130 38.265 0.730 38.880 ;
        RECT 0.130 38.035 1.860 38.265 ;
        RECT 2.160 38.035 3.820 38.265 ;
        RECT 0.130 36.025 0.730 38.035 ;
        RECT 2.160 37.000 2.390 38.035 ;
        RECT 2.795 36.745 3.025 37.790 ;
        RECT 4.050 36.745 4.650 38.880 ;
        RECT 5.840 38.640 6.460 38.825 ;
        RECT 37.440 38.640 38.060 38.825 ;
        RECT 5.840 38.410 38.060 38.640 ;
        RECT 5.840 38.225 6.460 38.410 ;
        RECT 37.440 38.225 38.060 38.410 ;
        RECT 38.290 38.640 38.910 38.825 ;
        RECT 69.890 38.640 70.510 38.825 ;
        RECT 38.290 38.410 70.510 38.640 ;
        RECT 38.290 38.225 38.910 38.410 ;
        RECT 69.890 38.225 70.510 38.410 ;
        RECT 70.740 38.640 71.360 38.825 ;
        RECT 102.340 38.640 102.960 38.825 ;
        RECT 70.740 38.410 102.960 38.640 ;
        RECT 70.740 38.225 71.360 38.410 ;
        RECT 102.340 38.225 102.960 38.410 ;
        RECT 103.190 38.640 103.810 38.825 ;
        RECT 134.790 38.640 135.410 38.825 ;
        RECT 103.190 38.410 135.410 38.640 ;
        RECT 103.190 38.225 103.810 38.410 ;
        RECT 134.790 38.225 135.410 38.410 ;
        RECT 33.440 38.145 35.060 38.155 ;
        RECT 65.890 38.145 67.510 38.155 ;
        RECT 98.340 38.145 99.960 38.155 ;
        RECT 130.790 38.145 132.410 38.155 ;
        RECT 6.690 37.775 37.210 38.145 ;
        RECT 39.140 37.775 69.660 38.145 ;
        RECT 71.590 37.775 102.110 38.145 ;
        RECT 104.040 37.775 134.560 38.145 ;
        RECT 6.690 37.055 37.210 37.435 ;
        RECT 39.140 37.055 69.660 37.435 ;
        RECT 71.590 37.055 102.110 37.435 ;
        RECT 104.040 37.055 134.560 37.435 ;
        RECT 0.960 36.515 3.025 36.745 ;
        RECT 3.255 36.515 4.650 36.745 ;
        RECT 0.130 35.795 1.860 36.025 ;
        RECT 2.160 35.795 3.820 36.025 ;
        RECT 0.130 33.785 0.730 35.795 ;
        RECT 2.160 34.760 2.390 35.795 ;
        RECT 2.795 34.505 3.025 35.550 ;
        RECT 4.050 34.505 4.650 36.515 ;
        RECT 5.840 36.800 6.460 36.985 ;
        RECT 37.440 36.800 38.060 36.985 ;
        RECT 5.840 36.570 38.060 36.800 ;
        RECT 5.840 36.385 6.460 36.570 ;
        RECT 37.440 36.385 38.060 36.570 ;
        RECT 38.290 36.800 38.910 36.985 ;
        RECT 69.890 36.800 70.510 36.985 ;
        RECT 38.290 36.570 70.510 36.800 ;
        RECT 38.290 36.385 38.910 36.570 ;
        RECT 69.890 36.385 70.510 36.570 ;
        RECT 70.740 36.800 71.360 36.985 ;
        RECT 102.340 36.800 102.960 36.985 ;
        RECT 70.740 36.570 102.960 36.800 ;
        RECT 70.740 36.385 71.360 36.570 ;
        RECT 102.340 36.385 102.960 36.570 ;
        RECT 103.190 36.800 103.810 36.985 ;
        RECT 134.790 36.800 135.410 36.985 ;
        RECT 103.190 36.570 135.410 36.800 ;
        RECT 103.190 36.385 103.810 36.570 ;
        RECT 134.790 36.385 135.410 36.570 ;
        RECT 29.600 36.305 31.220 36.315 ;
        RECT 62.050 36.305 63.670 36.315 ;
        RECT 94.500 36.305 96.120 36.315 ;
        RECT 126.950 36.305 128.570 36.315 ;
        RECT 6.690 35.935 37.210 36.305 ;
        RECT 39.140 35.935 69.660 36.305 ;
        RECT 71.590 35.935 102.110 36.305 ;
        RECT 104.040 35.935 134.560 36.305 ;
        RECT 6.700 35.140 37.200 35.580 ;
        RECT 39.150 35.140 69.650 35.580 ;
        RECT 71.600 35.140 102.100 35.580 ;
        RECT 104.050 35.140 134.550 35.580 ;
        RECT 0.960 34.275 3.025 34.505 ;
        RECT 3.255 34.275 4.650 34.505 ;
        RECT 6.690 34.410 37.210 34.790 ;
        RECT 39.140 34.410 69.660 34.790 ;
        RECT 71.590 34.410 102.110 34.790 ;
        RECT 104.040 34.410 134.560 34.790 ;
        RECT 0.130 33.555 1.860 33.785 ;
        RECT 2.160 33.555 3.820 33.785 ;
        RECT 0.130 31.545 0.730 33.555 ;
        RECT 2.160 32.520 2.390 33.555 ;
        RECT 2.795 32.265 3.025 33.310 ;
        RECT 4.050 32.265 4.650 34.275 ;
        RECT 5.840 34.155 6.460 34.340 ;
        RECT 37.440 34.155 38.060 34.340 ;
        RECT 5.840 33.925 38.060 34.155 ;
        RECT 5.840 33.740 6.460 33.925 ;
        RECT 37.440 33.740 38.060 33.925 ;
        RECT 38.290 34.155 38.910 34.340 ;
        RECT 69.890 34.155 70.510 34.340 ;
        RECT 38.290 33.925 70.510 34.155 ;
        RECT 38.290 33.740 38.910 33.925 ;
        RECT 69.890 33.740 70.510 33.925 ;
        RECT 70.740 34.155 71.360 34.340 ;
        RECT 102.340 34.155 102.960 34.340 ;
        RECT 70.740 33.925 102.960 34.155 ;
        RECT 70.740 33.740 71.360 33.925 ;
        RECT 102.340 33.740 102.960 33.925 ;
        RECT 103.190 34.155 103.810 34.340 ;
        RECT 134.790 34.155 135.410 34.340 ;
        RECT 103.190 33.925 135.410 34.155 ;
        RECT 103.190 33.740 103.810 33.925 ;
        RECT 134.790 33.740 135.410 33.925 ;
        RECT 25.760 33.660 27.380 33.670 ;
        RECT 58.210 33.660 59.830 33.670 ;
        RECT 90.660 33.660 92.280 33.670 ;
        RECT 123.110 33.660 124.730 33.670 ;
        RECT 6.690 33.290 37.210 33.660 ;
        RECT 39.140 33.290 69.660 33.660 ;
        RECT 71.590 33.290 102.110 33.660 ;
        RECT 104.040 33.290 134.560 33.660 ;
        RECT 6.690 32.570 37.210 32.950 ;
        RECT 39.140 32.570 69.660 32.950 ;
        RECT 71.590 32.570 102.110 32.950 ;
        RECT 104.040 32.570 134.560 32.950 ;
        RECT 0.960 32.035 3.025 32.265 ;
        RECT 3.255 32.035 4.650 32.265 ;
        RECT 0.130 31.315 1.860 31.545 ;
        RECT 2.160 31.315 3.820 31.545 ;
        RECT 0.130 29.305 0.730 31.315 ;
        RECT 2.160 30.280 2.390 31.315 ;
        RECT 2.795 30.025 3.025 31.070 ;
        RECT 4.050 30.025 4.650 32.035 ;
        RECT 5.840 32.315 6.460 32.500 ;
        RECT 37.440 32.315 38.060 32.500 ;
        RECT 5.840 32.085 38.060 32.315 ;
        RECT 5.840 31.900 6.460 32.085 ;
        RECT 37.440 31.900 38.060 32.085 ;
        RECT 38.290 32.315 38.910 32.500 ;
        RECT 69.890 32.315 70.510 32.500 ;
        RECT 38.290 32.085 70.510 32.315 ;
        RECT 38.290 31.900 38.910 32.085 ;
        RECT 69.890 31.900 70.510 32.085 ;
        RECT 70.740 32.315 71.360 32.500 ;
        RECT 102.340 32.315 102.960 32.500 ;
        RECT 70.740 32.085 102.960 32.315 ;
        RECT 70.740 31.900 71.360 32.085 ;
        RECT 102.340 31.900 102.960 32.085 ;
        RECT 103.190 32.315 103.810 32.500 ;
        RECT 134.790 32.315 135.410 32.500 ;
        RECT 103.190 32.085 135.410 32.315 ;
        RECT 103.190 31.900 103.810 32.085 ;
        RECT 134.790 31.900 135.410 32.085 ;
        RECT 21.920 31.820 23.540 31.830 ;
        RECT 54.370 31.820 55.990 31.830 ;
        RECT 86.820 31.820 88.440 31.830 ;
        RECT 119.270 31.820 120.890 31.830 ;
        RECT 6.690 31.450 37.210 31.820 ;
        RECT 39.140 31.450 69.660 31.820 ;
        RECT 71.590 31.450 102.110 31.820 ;
        RECT 104.040 31.450 134.560 31.820 ;
        RECT 6.690 30.730 37.210 31.110 ;
        RECT 39.140 30.730 69.660 31.110 ;
        RECT 71.590 30.730 102.110 31.110 ;
        RECT 104.040 30.730 134.560 31.110 ;
        RECT 5.840 30.475 6.460 30.660 ;
        RECT 37.440 30.475 38.060 30.660 ;
        RECT 5.840 30.245 38.060 30.475 ;
        RECT 5.840 30.060 6.460 30.245 ;
        RECT 37.440 30.060 38.060 30.245 ;
        RECT 38.290 30.475 38.910 30.660 ;
        RECT 69.890 30.475 70.510 30.660 ;
        RECT 38.290 30.245 70.510 30.475 ;
        RECT 38.290 30.060 38.910 30.245 ;
        RECT 69.890 30.060 70.510 30.245 ;
        RECT 70.740 30.475 71.360 30.660 ;
        RECT 102.340 30.475 102.960 30.660 ;
        RECT 70.740 30.245 102.960 30.475 ;
        RECT 70.740 30.060 71.360 30.245 ;
        RECT 102.340 30.060 102.960 30.245 ;
        RECT 103.190 30.475 103.810 30.660 ;
        RECT 134.790 30.475 135.410 30.660 ;
        RECT 103.190 30.245 135.410 30.475 ;
        RECT 103.190 30.060 103.810 30.245 ;
        RECT 134.790 30.060 135.410 30.245 ;
        RECT 0.960 29.795 3.025 30.025 ;
        RECT 3.255 29.795 4.650 30.025 ;
        RECT 18.080 29.980 19.700 29.990 ;
        RECT 50.530 29.980 52.150 29.990 ;
        RECT 82.980 29.980 84.600 29.990 ;
        RECT 115.430 29.980 117.050 29.990 ;
        RECT 0.130 29.075 1.860 29.305 ;
        RECT 2.160 29.075 3.820 29.305 ;
        RECT 0.130 26.920 0.730 29.075 ;
        RECT 2.160 28.040 2.390 29.075 ;
        RECT 2.795 27.785 3.025 28.830 ;
        RECT 4.050 27.785 4.650 29.795 ;
        RECT 6.690 29.610 37.210 29.980 ;
        RECT 39.140 29.610 69.660 29.980 ;
        RECT 71.590 29.610 102.110 29.980 ;
        RECT 104.040 29.610 134.560 29.980 ;
        RECT 6.700 28.815 37.200 29.255 ;
        RECT 39.150 28.815 69.650 29.255 ;
        RECT 71.600 28.815 102.100 29.255 ;
        RECT 104.050 28.815 134.550 29.255 ;
        RECT 6.690 28.085 37.210 28.465 ;
        RECT 39.140 28.085 69.660 28.465 ;
        RECT 71.590 28.085 102.110 28.465 ;
        RECT 104.040 28.085 134.560 28.465 ;
        RECT 0.960 27.555 3.025 27.785 ;
        RECT 3.255 27.555 4.650 27.785 ;
        RECT 4.050 26.920 4.650 27.555 ;
        RECT 5.840 27.830 6.460 28.015 ;
        RECT 37.440 27.830 38.060 28.015 ;
        RECT 5.840 27.600 38.060 27.830 ;
        RECT 5.840 27.415 6.460 27.600 ;
        RECT 37.440 27.415 38.060 27.600 ;
        RECT 38.290 27.830 38.910 28.015 ;
        RECT 69.890 27.830 70.510 28.015 ;
        RECT 38.290 27.600 70.510 27.830 ;
        RECT 38.290 27.415 38.910 27.600 ;
        RECT 69.890 27.415 70.510 27.600 ;
        RECT 70.740 27.830 71.360 28.015 ;
        RECT 102.340 27.830 102.960 28.015 ;
        RECT 70.740 27.600 102.960 27.830 ;
        RECT 70.740 27.415 71.360 27.600 ;
        RECT 102.340 27.415 102.960 27.600 ;
        RECT 103.190 27.830 103.810 28.015 ;
        RECT 134.790 27.830 135.410 28.015 ;
        RECT 103.190 27.600 135.410 27.830 ;
        RECT 103.190 27.415 103.810 27.600 ;
        RECT 134.790 27.415 135.410 27.600 ;
        RECT 14.240 27.335 15.860 27.345 ;
        RECT 46.690 27.335 48.310 27.345 ;
        RECT 79.140 27.335 80.760 27.345 ;
        RECT 111.590 27.335 113.210 27.345 ;
        RECT 6.690 26.965 37.210 27.335 ;
        RECT 39.140 26.965 69.660 27.335 ;
        RECT 71.590 26.965 102.110 27.335 ;
        RECT 104.040 26.965 134.560 27.335 ;
        RECT 0.130 26.580 2.420 26.920 ;
        RECT 3.165 26.580 4.650 26.920 ;
        RECT 0.130 25.945 0.730 26.580 ;
        RECT 0.130 25.715 1.860 25.945 ;
        RECT 2.160 25.715 3.820 25.945 ;
        RECT 0.130 23.705 0.730 25.715 ;
        RECT 2.160 24.680 2.390 25.715 ;
        RECT 2.795 24.425 3.025 25.470 ;
        RECT 4.050 24.425 4.650 26.580 ;
        RECT 6.690 26.245 37.210 26.625 ;
        RECT 39.140 26.245 69.660 26.625 ;
        RECT 71.590 26.245 102.110 26.625 ;
        RECT 104.040 26.245 134.560 26.625 ;
        RECT 5.840 25.990 6.460 26.175 ;
        RECT 37.440 25.990 38.060 26.175 ;
        RECT 5.840 25.760 38.060 25.990 ;
        RECT 5.840 25.575 6.460 25.760 ;
        RECT 37.440 25.575 38.060 25.760 ;
        RECT 38.290 25.990 38.910 26.175 ;
        RECT 69.890 25.990 70.510 26.175 ;
        RECT 38.290 25.760 70.510 25.990 ;
        RECT 38.290 25.575 38.910 25.760 ;
        RECT 69.890 25.575 70.510 25.760 ;
        RECT 70.740 25.990 71.360 26.175 ;
        RECT 102.340 25.990 102.960 26.175 ;
        RECT 70.740 25.760 102.960 25.990 ;
        RECT 70.740 25.575 71.360 25.760 ;
        RECT 102.340 25.575 102.960 25.760 ;
        RECT 103.190 25.990 103.810 26.175 ;
        RECT 134.790 25.990 135.410 26.175 ;
        RECT 103.190 25.760 135.410 25.990 ;
        RECT 103.190 25.575 103.810 25.760 ;
        RECT 134.790 25.575 135.410 25.760 ;
        RECT 10.400 25.495 12.020 25.505 ;
        RECT 42.850 25.495 44.470 25.505 ;
        RECT 75.300 25.495 76.920 25.505 ;
        RECT 107.750 25.495 109.370 25.505 ;
        RECT 6.690 25.125 37.210 25.495 ;
        RECT 39.140 25.125 69.660 25.495 ;
        RECT 71.590 25.125 102.110 25.495 ;
        RECT 104.040 25.125 134.560 25.495 ;
        RECT 0.960 24.195 3.025 24.425 ;
        RECT 3.255 24.195 4.650 24.425 ;
        RECT 6.690 24.405 37.210 24.785 ;
        RECT 39.140 24.405 69.660 24.785 ;
        RECT 71.590 24.405 102.110 24.785 ;
        RECT 104.040 24.405 134.560 24.785 ;
        RECT 0.130 23.475 1.860 23.705 ;
        RECT 2.160 23.475 3.820 23.705 ;
        RECT 0.130 21.320 0.730 23.475 ;
        RECT 2.160 22.440 2.390 23.475 ;
        RECT 2.795 22.185 3.025 23.230 ;
        RECT 4.050 22.185 4.650 24.195 ;
        RECT 5.840 24.150 6.460 24.335 ;
        RECT 37.440 24.150 38.060 24.335 ;
        RECT 5.840 23.920 38.060 24.150 ;
        RECT 5.840 23.735 6.460 23.920 ;
        RECT 37.440 23.735 38.060 23.920 ;
        RECT 38.290 24.150 38.910 24.335 ;
        RECT 69.890 24.150 70.510 24.335 ;
        RECT 38.290 23.920 70.510 24.150 ;
        RECT 38.290 23.735 38.910 23.920 ;
        RECT 69.890 23.735 70.510 23.920 ;
        RECT 70.740 24.150 71.360 24.335 ;
        RECT 102.340 24.150 102.960 24.335 ;
        RECT 70.740 23.920 102.960 24.150 ;
        RECT 70.740 23.735 71.360 23.920 ;
        RECT 102.340 23.735 102.960 23.920 ;
        RECT 103.190 24.150 103.810 24.335 ;
        RECT 134.790 24.150 135.410 24.335 ;
        RECT 103.190 23.920 135.410 24.150 ;
        RECT 103.190 23.735 103.810 23.920 ;
        RECT 134.790 23.735 135.410 23.920 ;
        RECT 6.690 23.285 37.210 23.655 ;
        RECT 39.140 23.285 69.660 23.655 ;
        RECT 71.590 23.285 102.110 23.655 ;
        RECT 104.040 23.285 134.560 23.655 ;
        RECT 0.960 21.955 3.025 22.185 ;
        RECT 3.255 21.955 4.650 22.185 ;
        RECT 4.050 21.320 4.650 21.955 ;
        RECT 0.130 20.980 2.420 21.320 ;
        RECT 3.165 20.980 4.650 21.320 ;
        RECT 0.130 20.345 0.730 20.980 ;
        RECT 0.130 20.115 1.710 20.345 ;
        RECT 0.130 18.075 0.730 20.115 ;
        RECT 2.140 19.885 2.500 19.970 ;
        RECT 1.010 19.655 2.500 19.885 ;
        RECT 1.010 19.505 1.370 19.655 ;
        RECT 0.960 18.870 1.910 19.275 ;
        RECT 0.130 17.845 1.420 18.075 ;
        RECT 0.130 16.885 0.730 17.845 ;
        RECT 1.650 17.525 1.910 18.870 ;
        RECT 2.140 18.220 2.500 19.655 ;
        RECT 2.730 18.320 3.080 19.520 ;
        RECT 3.440 18.910 3.820 20.555 ;
        RECT 2.520 17.525 2.870 17.585 ;
        RECT 3.440 17.525 3.780 18.130 ;
        RECT 1.650 17.265 3.780 17.525 ;
        RECT 2.520 17.205 2.870 17.265 ;
        RECT 4.050 16.985 4.650 20.980 ;
        RECT 6.495 20.500 8.245 23.285 ;
        RECT 8.885 20.500 9.695 21.500 ;
        RECT 10.335 20.500 12.085 22.795 ;
        RECT 12.725 20.500 13.535 21.500 ;
        RECT 14.175 20.500 15.925 22.795 ;
        RECT 16.565 20.500 17.375 21.500 ;
        RECT 18.015 20.500 19.765 22.795 ;
        RECT 20.405 20.500 21.215 21.500 ;
        RECT 21.855 20.500 23.605 22.795 ;
        RECT 24.245 20.500 25.055 21.500 ;
        RECT 25.695 20.500 27.445 22.795 ;
        RECT 28.085 20.500 28.895 21.500 ;
        RECT 29.535 20.500 31.285 22.795 ;
        RECT 31.925 20.500 32.735 21.500 ;
        RECT 33.375 20.500 35.125 22.795 ;
        RECT 35.765 20.500 36.575 21.500 ;
        RECT 38.945 20.500 40.695 23.285 ;
        RECT 41.335 20.500 42.145 21.500 ;
        RECT 42.785 20.500 44.535 22.795 ;
        RECT 45.175 20.500 45.985 21.500 ;
        RECT 46.625 20.500 48.375 22.795 ;
        RECT 49.015 20.500 49.825 21.500 ;
        RECT 50.465 20.500 52.215 22.795 ;
        RECT 52.855 20.500 53.665 21.500 ;
        RECT 54.305 20.500 56.055 22.795 ;
        RECT 56.695 20.500 57.505 21.500 ;
        RECT 58.145 20.500 59.895 22.795 ;
        RECT 60.535 20.500 61.345 21.500 ;
        RECT 61.985 20.500 63.735 22.795 ;
        RECT 64.375 20.500 65.185 21.500 ;
        RECT 65.825 20.500 67.575 22.795 ;
        RECT 68.215 20.500 69.025 21.500 ;
        RECT 71.395 20.500 73.145 23.285 ;
        RECT 73.785 20.500 74.595 21.500 ;
        RECT 75.235 20.500 76.985 22.795 ;
        RECT 77.625 20.500 78.435 21.500 ;
        RECT 79.075 20.500 80.825 22.795 ;
        RECT 81.465 20.500 82.275 21.500 ;
        RECT 82.915 20.500 84.665 22.795 ;
        RECT 85.305 20.500 86.115 21.500 ;
        RECT 86.755 20.500 88.505 22.795 ;
        RECT 89.145 20.500 89.955 21.500 ;
        RECT 90.595 20.500 92.345 22.795 ;
        RECT 92.985 20.500 93.795 21.500 ;
        RECT 94.435 20.500 96.185 22.795 ;
        RECT 96.825 20.500 97.635 21.500 ;
        RECT 98.275 20.500 100.025 22.795 ;
        RECT 100.665 20.500 101.475 21.500 ;
        RECT 103.845 20.500 105.595 23.285 ;
        RECT 106.235 20.500 107.045 21.500 ;
        RECT 107.685 20.500 109.435 22.795 ;
        RECT 110.075 20.500 110.885 21.500 ;
        RECT 111.525 20.500 113.275 22.795 ;
        RECT 113.915 20.500 114.725 21.500 ;
        RECT 115.365 20.500 117.115 22.795 ;
        RECT 117.755 20.500 118.565 21.500 ;
        RECT 119.205 20.500 120.955 22.795 ;
        RECT 121.595 20.500 122.405 21.500 ;
        RECT 123.045 20.500 124.795 22.795 ;
        RECT 125.435 20.500 126.245 21.500 ;
        RECT 126.885 20.500 128.635 22.795 ;
        RECT 129.275 20.500 130.085 21.500 ;
        RECT 130.725 20.500 132.475 22.795 ;
        RECT 133.115 20.500 133.925 21.500 ;
        RECT 136.340 20.690 136.710 39.200 ;
        RECT 137.360 35.565 137.730 39.200 ;
        RECT 137.355 35.185 137.735 35.565 ;
        RECT 137.360 32.565 137.730 35.185 ;
        RECT 137.355 32.185 137.735 32.565 ;
        RECT 137.360 29.565 137.730 32.185 ;
        RECT 137.355 29.185 137.735 29.565 ;
        RECT 137.360 26.565 137.730 29.185 ;
        RECT 137.355 26.185 137.735 26.565 ;
        RECT 137.360 23.565 137.730 26.185 ;
        RECT 137.355 23.185 137.735 23.565 ;
        RECT 136.340 20.310 136.720 20.690 ;
        RECT 136.340 19.240 136.710 20.310 ;
        RECT 6.965 18.050 7.775 19.050 ;
        RECT 0.130 16.655 1.820 16.885 ;
        RECT 3.190 16.755 4.650 16.985 ;
        RECT 0.130 14.645 0.730 16.655 ;
        RECT 2.150 16.195 3.150 16.520 ;
        RECT 0.960 15.635 3.820 15.965 ;
        RECT 0.130 14.415 1.820 14.645 ;
        RECT 0.130 12.405 0.730 14.415 ;
        RECT 2.535 14.280 2.800 15.635 ;
        RECT 4.050 14.745 4.650 16.755 ;
        RECT 8.415 16.220 10.165 19.050 ;
        RECT 10.805 18.050 11.615 19.050 ;
        RECT 12.255 16.755 14.005 19.050 ;
        RECT 14.645 18.050 15.455 19.050 ;
        RECT 16.095 16.755 17.845 19.050 ;
        RECT 18.485 18.050 19.295 19.050 ;
        RECT 19.935 16.755 21.685 19.050 ;
        RECT 22.325 18.050 23.135 19.050 ;
        RECT 23.775 16.755 25.525 19.050 ;
        RECT 26.165 18.050 26.975 19.050 ;
        RECT 27.615 16.755 29.365 19.050 ;
        RECT 30.005 18.050 30.815 19.050 ;
        RECT 31.455 16.755 33.205 19.050 ;
        RECT 33.845 18.050 34.655 19.050 ;
        RECT 35.295 16.755 37.045 19.050 ;
        RECT 39.415 18.050 40.225 19.050 ;
        RECT 40.865 16.220 42.615 19.050 ;
        RECT 43.255 18.050 44.065 19.050 ;
        RECT 44.705 16.755 46.455 19.050 ;
        RECT 47.095 18.050 47.905 19.050 ;
        RECT 48.545 16.755 50.295 19.050 ;
        RECT 50.935 18.050 51.745 19.050 ;
        RECT 52.385 16.755 54.135 19.050 ;
        RECT 54.775 18.050 55.585 19.050 ;
        RECT 56.225 16.755 57.975 19.050 ;
        RECT 58.615 18.050 59.425 19.050 ;
        RECT 60.065 16.755 61.815 19.050 ;
        RECT 62.455 18.050 63.265 19.050 ;
        RECT 63.905 16.755 65.655 19.050 ;
        RECT 66.295 18.050 67.105 19.050 ;
        RECT 67.745 16.755 69.495 19.050 ;
        RECT 71.865 18.050 72.675 19.050 ;
        RECT 73.315 16.220 75.065 19.050 ;
        RECT 75.705 18.050 76.515 19.050 ;
        RECT 77.155 16.755 78.905 19.050 ;
        RECT 79.545 18.050 80.355 19.050 ;
        RECT 80.995 16.755 82.745 19.050 ;
        RECT 83.385 18.050 84.195 19.050 ;
        RECT 84.835 16.755 86.585 19.050 ;
        RECT 87.225 18.050 88.035 19.050 ;
        RECT 88.675 16.755 90.425 19.050 ;
        RECT 91.065 18.050 91.875 19.050 ;
        RECT 92.515 16.755 94.265 19.050 ;
        RECT 94.905 18.050 95.715 19.050 ;
        RECT 96.355 16.755 98.105 19.050 ;
        RECT 98.745 18.050 99.555 19.050 ;
        RECT 100.195 16.755 101.945 19.050 ;
        RECT 104.315 18.050 105.125 19.050 ;
        RECT 105.765 16.220 107.515 19.050 ;
        RECT 108.155 18.050 108.965 19.050 ;
        RECT 109.605 16.755 111.355 19.050 ;
        RECT 111.995 18.050 112.805 19.050 ;
        RECT 113.445 16.755 115.195 19.050 ;
        RECT 115.835 18.050 116.645 19.050 ;
        RECT 117.285 16.755 119.035 19.050 ;
        RECT 119.675 18.050 120.485 19.050 ;
        RECT 121.125 16.755 122.875 19.050 ;
        RECT 123.515 18.050 124.325 19.050 ;
        RECT 124.965 16.755 126.715 19.050 ;
        RECT 127.355 18.050 128.165 19.050 ;
        RECT 128.805 16.755 130.555 19.050 ;
        RECT 131.195 18.050 132.005 19.050 ;
        RECT 132.645 16.755 134.395 19.050 ;
        RECT 136.340 18.860 136.720 19.240 ;
        RECT 6.690 15.850 37.210 16.220 ;
        RECT 39.140 15.850 69.660 16.220 ;
        RECT 71.590 15.850 102.110 16.220 ;
        RECT 104.040 15.850 134.560 16.220 ;
        RECT 5.840 15.585 6.460 15.770 ;
        RECT 37.440 15.585 38.060 15.770 ;
        RECT 5.840 15.355 38.060 15.585 ;
        RECT 5.840 15.170 6.460 15.355 ;
        RECT 37.440 15.170 38.060 15.355 ;
        RECT 38.290 15.585 38.910 15.770 ;
        RECT 69.890 15.585 70.510 15.770 ;
        RECT 38.290 15.355 70.510 15.585 ;
        RECT 38.290 15.170 38.910 15.355 ;
        RECT 69.890 15.170 70.510 15.355 ;
        RECT 70.740 15.585 71.360 15.770 ;
        RECT 102.340 15.585 102.960 15.770 ;
        RECT 70.740 15.355 102.960 15.585 ;
        RECT 70.740 15.170 71.360 15.355 ;
        RECT 102.340 15.170 102.960 15.355 ;
        RECT 103.190 15.585 103.810 15.770 ;
        RECT 134.790 15.585 135.410 15.770 ;
        RECT 103.190 15.355 135.410 15.585 ;
        RECT 103.190 15.170 103.810 15.355 ;
        RECT 134.790 15.170 135.410 15.355 ;
        RECT 3.190 14.515 4.650 14.745 ;
        RECT 6.690 14.720 37.210 15.100 ;
        RECT 39.140 14.720 69.660 15.100 ;
        RECT 71.590 14.720 102.110 15.100 ;
        RECT 104.040 14.720 134.560 15.100 ;
        RECT 2.150 13.955 3.150 14.280 ;
        RECT 0.960 13.395 3.820 13.725 ;
        RECT 4.050 12.505 4.650 14.515 ;
        RECT 6.690 14.010 37.210 14.380 ;
        RECT 39.140 14.010 69.660 14.380 ;
        RECT 71.590 14.010 102.110 14.380 ;
        RECT 104.040 14.010 134.560 14.380 ;
        RECT 12.320 14.000 13.940 14.010 ;
        RECT 44.770 14.000 46.390 14.010 ;
        RECT 77.220 14.000 78.840 14.010 ;
        RECT 109.670 14.000 111.290 14.010 ;
        RECT 5.840 13.745 6.460 13.930 ;
        RECT 37.440 13.745 38.060 13.930 ;
        RECT 5.840 13.515 38.060 13.745 ;
        RECT 5.840 13.330 6.460 13.515 ;
        RECT 37.440 13.330 38.060 13.515 ;
        RECT 38.290 13.745 38.910 13.930 ;
        RECT 69.890 13.745 70.510 13.930 ;
        RECT 38.290 13.515 70.510 13.745 ;
        RECT 38.290 13.330 38.910 13.515 ;
        RECT 69.890 13.330 70.510 13.515 ;
        RECT 70.740 13.745 71.360 13.930 ;
        RECT 102.340 13.745 102.960 13.930 ;
        RECT 70.740 13.515 102.960 13.745 ;
        RECT 70.740 13.330 71.360 13.515 ;
        RECT 102.340 13.330 102.960 13.515 ;
        RECT 103.190 13.745 103.810 13.930 ;
        RECT 134.790 13.745 135.410 13.930 ;
        RECT 103.190 13.515 135.410 13.745 ;
        RECT 103.190 13.330 103.810 13.515 ;
        RECT 134.790 13.330 135.410 13.515 ;
        RECT 6.690 12.880 37.210 13.260 ;
        RECT 39.140 12.880 69.660 13.260 ;
        RECT 71.590 12.880 102.110 13.260 ;
        RECT 104.040 12.880 134.560 13.260 ;
        RECT 0.130 12.175 1.820 12.405 ;
        RECT 3.190 12.275 4.650 12.505 ;
        RECT 0.130 10.120 0.730 12.175 ;
        RECT 2.150 11.715 3.150 12.040 ;
        RECT 0.960 11.155 3.820 11.485 ;
        RECT 2.300 11.030 2.680 11.155 ;
        RECT 4.050 10.120 4.650 12.275 ;
        RECT 6.690 12.165 37.210 12.535 ;
        RECT 39.140 12.165 69.660 12.535 ;
        RECT 71.590 12.165 102.110 12.535 ;
        RECT 104.040 12.165 134.560 12.535 ;
        RECT 16.160 12.155 17.780 12.165 ;
        RECT 48.610 12.155 50.230 12.165 ;
        RECT 81.060 12.155 82.680 12.165 ;
        RECT 113.510 12.155 115.130 12.165 ;
        RECT 5.840 11.900 6.460 12.085 ;
        RECT 37.440 11.900 38.060 12.085 ;
        RECT 5.840 11.670 38.060 11.900 ;
        RECT 5.840 11.485 6.460 11.670 ;
        RECT 37.440 11.485 38.060 11.670 ;
        RECT 38.290 11.900 38.910 12.085 ;
        RECT 69.890 11.900 70.510 12.085 ;
        RECT 38.290 11.670 70.510 11.900 ;
        RECT 38.290 11.485 38.910 11.670 ;
        RECT 69.890 11.485 70.510 11.670 ;
        RECT 70.740 11.900 71.360 12.085 ;
        RECT 102.340 11.900 102.960 12.085 ;
        RECT 70.740 11.670 102.960 11.900 ;
        RECT 70.740 11.485 71.360 11.670 ;
        RECT 102.340 11.485 102.960 11.670 ;
        RECT 103.190 11.900 103.810 12.085 ;
        RECT 134.790 11.900 135.410 12.085 ;
        RECT 103.190 11.670 135.410 11.900 ;
        RECT 103.190 11.485 103.810 11.670 ;
        RECT 134.790 11.485 135.410 11.670 ;
        RECT 6.690 11.035 37.210 11.415 ;
        RECT 39.140 11.035 69.660 11.415 ;
        RECT 71.590 11.035 102.110 11.415 ;
        RECT 104.040 11.035 134.560 11.415 ;
        RECT 6.700 10.245 37.200 10.685 ;
        RECT 39.150 10.245 69.650 10.685 ;
        RECT 71.600 10.245 102.100 10.685 ;
        RECT 104.050 10.245 134.550 10.685 ;
        RECT 0.130 9.780 2.420 10.120 ;
        RECT 3.165 9.780 4.650 10.120 ;
        RECT 0.130 9.000 0.730 9.780 ;
        RECT 4.050 9.000 4.650 9.780 ;
        RECT 6.690 9.525 37.210 9.895 ;
        RECT 39.140 9.525 69.660 9.895 ;
        RECT 71.590 9.525 102.110 9.895 ;
        RECT 104.040 9.525 134.560 9.895 ;
        RECT 20.000 9.515 21.620 9.525 ;
        RECT 52.450 9.515 54.070 9.525 ;
        RECT 84.900 9.515 86.520 9.525 ;
        RECT 117.350 9.515 118.970 9.525 ;
        RECT 0.130 8.660 2.420 9.000 ;
        RECT 3.165 8.660 4.650 9.000 ;
        RECT 5.840 9.260 6.460 9.445 ;
        RECT 37.440 9.260 38.060 9.445 ;
        RECT 5.840 9.030 38.060 9.260 ;
        RECT 5.840 8.845 6.460 9.030 ;
        RECT 37.440 8.845 38.060 9.030 ;
        RECT 38.290 9.260 38.910 9.445 ;
        RECT 69.890 9.260 70.510 9.445 ;
        RECT 38.290 9.030 70.510 9.260 ;
        RECT 38.290 8.845 38.910 9.030 ;
        RECT 69.890 8.845 70.510 9.030 ;
        RECT 70.740 9.260 71.360 9.445 ;
        RECT 102.340 9.260 102.960 9.445 ;
        RECT 70.740 9.030 102.960 9.260 ;
        RECT 70.740 8.845 71.360 9.030 ;
        RECT 102.340 8.845 102.960 9.030 ;
        RECT 103.190 9.260 103.810 9.445 ;
        RECT 134.790 9.260 135.410 9.445 ;
        RECT 103.190 9.030 135.410 9.260 ;
        RECT 103.190 8.845 103.810 9.030 ;
        RECT 134.790 8.845 135.410 9.030 ;
        RECT 0.130 8.025 0.730 8.660 ;
        RECT 0.130 7.795 1.860 8.025 ;
        RECT 2.160 7.795 3.820 8.025 ;
        RECT 0.130 5.785 0.730 7.795 ;
        RECT 2.160 6.760 2.390 7.795 ;
        RECT 2.795 6.505 3.025 7.550 ;
        RECT 4.050 6.505 4.650 8.660 ;
        RECT 6.690 8.395 37.210 8.775 ;
        RECT 39.140 8.395 69.660 8.775 ;
        RECT 71.590 8.395 102.110 8.775 ;
        RECT 104.040 8.395 134.560 8.775 ;
        RECT 6.690 7.685 37.210 8.055 ;
        RECT 39.140 7.685 69.660 8.055 ;
        RECT 71.590 7.685 102.110 8.055 ;
        RECT 104.040 7.685 134.560 8.055 ;
        RECT 23.840 7.675 25.460 7.685 ;
        RECT 56.290 7.675 57.910 7.685 ;
        RECT 88.740 7.675 90.360 7.685 ;
        RECT 121.190 7.675 122.810 7.685 ;
        RECT 5.840 7.420 6.460 7.605 ;
        RECT 37.440 7.420 38.060 7.605 ;
        RECT 5.840 7.190 38.060 7.420 ;
        RECT 5.840 7.005 6.460 7.190 ;
        RECT 37.440 7.005 38.060 7.190 ;
        RECT 38.290 7.420 38.910 7.605 ;
        RECT 69.890 7.420 70.510 7.605 ;
        RECT 38.290 7.190 70.510 7.420 ;
        RECT 38.290 7.005 38.910 7.190 ;
        RECT 69.890 7.005 70.510 7.190 ;
        RECT 70.740 7.420 71.360 7.605 ;
        RECT 102.340 7.420 102.960 7.605 ;
        RECT 70.740 7.190 102.960 7.420 ;
        RECT 70.740 7.005 71.360 7.190 ;
        RECT 102.340 7.005 102.960 7.190 ;
        RECT 103.190 7.420 103.810 7.605 ;
        RECT 134.790 7.420 135.410 7.605 ;
        RECT 103.190 7.190 135.410 7.420 ;
        RECT 103.190 7.005 103.810 7.190 ;
        RECT 134.790 7.005 135.410 7.190 ;
        RECT 6.690 6.555 37.210 6.935 ;
        RECT 39.140 6.555 69.660 6.935 ;
        RECT 71.590 6.555 102.110 6.935 ;
        RECT 104.040 6.555 134.560 6.935 ;
        RECT 0.960 6.275 3.025 6.505 ;
        RECT 3.255 6.275 4.650 6.505 ;
        RECT 0.130 5.555 1.860 5.785 ;
        RECT 2.160 5.555 3.820 5.785 ;
        RECT 0.130 3.545 0.730 5.555 ;
        RECT 2.160 4.520 2.390 5.555 ;
        RECT 2.795 4.265 3.025 5.310 ;
        RECT 4.050 4.265 4.650 6.275 ;
        RECT 6.690 5.840 37.210 6.210 ;
        RECT 39.140 5.840 69.660 6.210 ;
        RECT 71.590 5.840 102.110 6.210 ;
        RECT 104.040 5.840 134.560 6.210 ;
        RECT 27.680 5.830 29.300 5.840 ;
        RECT 60.130 5.830 61.750 5.840 ;
        RECT 92.580 5.830 94.200 5.840 ;
        RECT 125.030 5.830 126.650 5.840 ;
        RECT 5.840 5.575 6.460 5.760 ;
        RECT 37.440 5.575 38.060 5.760 ;
        RECT 5.840 5.345 38.060 5.575 ;
        RECT 5.840 5.160 6.460 5.345 ;
        RECT 37.440 5.160 38.060 5.345 ;
        RECT 38.290 5.575 38.910 5.760 ;
        RECT 69.890 5.575 70.510 5.760 ;
        RECT 38.290 5.345 70.510 5.575 ;
        RECT 38.290 5.160 38.910 5.345 ;
        RECT 69.890 5.160 70.510 5.345 ;
        RECT 70.740 5.575 71.360 5.760 ;
        RECT 102.340 5.575 102.960 5.760 ;
        RECT 70.740 5.345 102.960 5.575 ;
        RECT 70.740 5.160 71.360 5.345 ;
        RECT 102.340 5.160 102.960 5.345 ;
        RECT 103.190 5.575 103.810 5.760 ;
        RECT 134.790 5.575 135.410 5.760 ;
        RECT 103.190 5.345 135.410 5.575 ;
        RECT 103.190 5.160 103.810 5.345 ;
        RECT 134.790 5.160 135.410 5.345 ;
        RECT 6.690 4.710 37.210 5.090 ;
        RECT 39.140 4.710 69.660 5.090 ;
        RECT 71.590 4.710 102.110 5.090 ;
        RECT 104.040 4.710 134.560 5.090 ;
        RECT 0.960 4.035 3.025 4.265 ;
        RECT 3.255 4.035 4.650 4.265 ;
        RECT 0.130 3.315 1.860 3.545 ;
        RECT 2.160 3.315 3.820 3.545 ;
        RECT 0.130 1.140 0.730 3.315 ;
        RECT 2.160 2.280 2.390 3.315 ;
        RECT 2.795 2.025 3.025 3.070 ;
        RECT 4.050 2.025 4.650 4.035 ;
        RECT 6.700 3.920 37.200 4.360 ;
        RECT 39.150 3.920 69.650 4.360 ;
        RECT 71.600 3.920 102.100 4.360 ;
        RECT 104.050 3.920 134.550 4.360 ;
        RECT 6.690 3.200 37.210 3.570 ;
        RECT 39.140 3.200 69.660 3.570 ;
        RECT 71.590 3.200 102.110 3.570 ;
        RECT 104.040 3.200 134.560 3.570 ;
        RECT 31.520 3.190 33.140 3.200 ;
        RECT 63.970 3.190 65.590 3.200 ;
        RECT 96.420 3.190 98.040 3.200 ;
        RECT 128.870 3.190 130.490 3.200 ;
        RECT 5.840 2.935 6.460 3.120 ;
        RECT 37.440 2.935 38.060 3.120 ;
        RECT 5.840 2.705 38.060 2.935 ;
        RECT 5.840 2.520 6.460 2.705 ;
        RECT 37.440 2.520 38.060 2.705 ;
        RECT 38.290 2.935 38.910 3.120 ;
        RECT 69.890 2.935 70.510 3.120 ;
        RECT 38.290 2.705 70.510 2.935 ;
        RECT 38.290 2.520 38.910 2.705 ;
        RECT 69.890 2.520 70.510 2.705 ;
        RECT 70.740 2.935 71.360 3.120 ;
        RECT 102.340 2.935 102.960 3.120 ;
        RECT 70.740 2.705 102.960 2.935 ;
        RECT 70.740 2.520 71.360 2.705 ;
        RECT 102.340 2.520 102.960 2.705 ;
        RECT 103.190 2.935 103.810 3.120 ;
        RECT 134.790 2.935 135.410 3.120 ;
        RECT 103.190 2.705 135.410 2.935 ;
        RECT 103.190 2.520 103.810 2.705 ;
        RECT 134.790 2.520 135.410 2.705 ;
        RECT 6.690 2.070 37.210 2.450 ;
        RECT 39.140 2.070 69.660 2.450 ;
        RECT 71.590 2.070 102.110 2.450 ;
        RECT 104.040 2.070 134.560 2.450 ;
        RECT 0.960 1.795 3.025 2.025 ;
        RECT 3.255 1.795 4.650 2.025 ;
        RECT 4.050 1.140 4.650 1.795 ;
        RECT 6.690 1.360 37.210 1.730 ;
        RECT 39.140 1.360 69.660 1.730 ;
        RECT 71.590 1.360 102.110 1.730 ;
        RECT 104.040 1.360 134.560 1.730 ;
        RECT 35.360 1.350 36.980 1.360 ;
        RECT 67.810 1.350 69.430 1.360 ;
        RECT 100.260 1.350 101.880 1.360 ;
        RECT 132.710 1.350 134.330 1.360 ;
        RECT 0.130 0.800 2.430 1.140 ;
        RECT 3.160 0.800 4.650 1.140 ;
        RECT 0.130 0.000 0.730 0.800 ;
        RECT 4.050 0.000 4.650 0.800 ;
        RECT 5.840 1.095 6.460 1.280 ;
        RECT 37.440 1.095 38.060 1.280 ;
        RECT 5.840 0.865 38.060 1.095 ;
        RECT 5.840 0.680 6.460 0.865 ;
        RECT 37.440 0.680 38.060 0.865 ;
        RECT 38.290 1.095 38.910 1.280 ;
        RECT 69.890 1.095 70.510 1.280 ;
        RECT 38.290 0.865 70.510 1.095 ;
        RECT 38.290 0.680 38.910 0.865 ;
        RECT 69.890 0.680 70.510 0.865 ;
        RECT 70.740 1.095 71.360 1.280 ;
        RECT 102.340 1.095 102.960 1.280 ;
        RECT 70.740 0.865 102.960 1.095 ;
        RECT 70.740 0.680 71.360 0.865 ;
        RECT 102.340 0.680 102.960 0.865 ;
        RECT 103.190 1.095 103.810 1.280 ;
        RECT 134.790 1.095 135.410 1.280 ;
        RECT 103.190 0.865 135.410 1.095 ;
        RECT 136.340 0.930 136.710 18.860 ;
        RECT 137.360 17.565 137.730 23.185 ;
        RECT 138.380 20.690 138.750 39.200 ;
        RECT 139.400 35.565 139.770 39.200 ;
        RECT 139.395 35.185 139.775 35.565 ;
        RECT 139.400 32.565 139.770 35.185 ;
        RECT 139.395 32.185 139.775 32.565 ;
        RECT 139.400 29.565 139.770 32.185 ;
        RECT 139.395 29.185 139.775 29.565 ;
        RECT 139.400 26.565 139.770 29.185 ;
        RECT 139.395 26.185 139.775 26.565 ;
        RECT 139.400 23.565 139.770 26.185 ;
        RECT 139.395 23.185 139.775 23.565 ;
        RECT 138.380 20.310 138.760 20.690 ;
        RECT 138.380 19.240 138.750 20.310 ;
        RECT 138.380 18.860 138.760 19.240 ;
        RECT 137.355 17.185 137.735 17.565 ;
        RECT 137.360 14.565 137.730 17.185 ;
        RECT 137.355 14.185 137.735 14.565 ;
        RECT 137.360 11.565 137.730 14.185 ;
        RECT 137.355 11.185 137.735 11.565 ;
        RECT 137.360 8.565 137.730 11.185 ;
        RECT 137.355 8.185 137.735 8.565 ;
        RECT 137.360 5.565 137.730 8.185 ;
        RECT 137.355 5.185 137.735 5.565 ;
        RECT 137.360 2.565 137.730 5.185 ;
        RECT 137.355 2.185 137.735 2.565 ;
        RECT 137.360 0.930 137.730 2.185 ;
        RECT 138.380 0.930 138.750 18.860 ;
        RECT 139.400 17.565 139.770 23.185 ;
        RECT 139.395 17.185 139.775 17.565 ;
        RECT 139.400 14.565 139.770 17.185 ;
        RECT 139.395 14.185 139.775 14.565 ;
        RECT 139.400 11.565 139.770 14.185 ;
        RECT 139.395 11.185 139.775 11.565 ;
        RECT 139.400 8.565 139.770 11.185 ;
        RECT 139.395 8.185 139.775 8.565 ;
        RECT 139.400 5.565 139.770 8.185 ;
        RECT 139.395 5.185 139.775 5.565 ;
        RECT 139.400 2.565 139.770 5.185 ;
        RECT 139.395 2.185 139.775 2.565 ;
        RECT 139.400 0.930 139.770 2.185 ;
        RECT 140.420 0.930 140.800 39.200 ;
        RECT 141.150 0.940 141.590 39.190 ;
        RECT 103.190 0.680 103.810 0.865 ;
        RECT 134.790 0.680 135.410 0.865 ;
        RECT 6.690 0.230 37.210 0.610 ;
        RECT 39.140 0.230 69.660 0.610 ;
        RECT 71.590 0.230 102.110 0.610 ;
        RECT 104.040 0.230 134.560 0.610 ;
      LAYER Metal2 ;
        RECT 6.700 314.590 9.560 314.970 ;
        RECT 39.150 314.590 42.010 314.970 ;
        RECT 71.600 314.590 74.460 314.970 ;
        RECT 104.050 314.590 106.910 314.970 ;
        RECT 37.560 314.030 37.940 314.410 ;
        RECT 70.010 314.030 70.390 314.410 ;
        RECT 102.460 314.030 102.840 314.410 ;
        RECT 134.910 314.030 135.290 314.410 ;
        RECT 0.240 312.380 0.620 312.760 ;
        RECT 4.160 312.380 4.540 312.760 ;
        RECT 6.700 312.750 9.560 313.130 ;
        RECT 6.700 310.865 9.560 311.245 ;
        RECT 6.700 310.105 9.560 310.485 ;
        RECT 0.240 309.380 0.620 309.760 ;
        RECT 4.160 309.380 4.540 309.760 ;
        RECT 6.700 308.265 9.560 308.645 ;
        RECT 0.240 306.380 0.620 306.760 ;
        RECT 4.160 306.380 4.540 306.760 ;
        RECT 6.700 306.425 9.560 306.805 ;
        RECT 6.700 304.540 9.560 304.920 ;
        RECT 6.700 303.780 9.560 304.160 ;
        RECT 0.240 303.380 0.620 303.760 ;
        RECT 4.160 303.380 4.540 303.760 ;
        RECT 6.700 301.940 9.560 302.320 ;
        RECT 0.240 300.380 0.620 300.760 ;
        RECT 4.160 300.380 4.540 300.760 ;
        RECT 6.700 300.100 9.560 300.480 ;
        RECT 0.240 297.380 0.620 297.760 ;
        RECT 4.160 297.380 4.540 297.760 ;
        RECT 10.335 297.390 12.085 301.200 ;
        RECT 14.175 297.390 15.925 303.040 ;
        RECT 18.015 297.390 19.765 305.685 ;
        RECT 21.855 297.390 23.605 307.525 ;
        RECT 25.695 297.390 27.445 309.365 ;
        RECT 29.535 297.390 31.285 312.010 ;
        RECT 33.375 297.390 35.125 313.850 ;
        RECT 39.150 312.750 42.010 313.130 ;
        RECT 37.560 312.190 37.940 312.570 ;
        RECT 39.150 310.865 42.010 311.245 ;
        RECT 39.150 310.105 42.010 310.485 ;
        RECT 37.560 309.545 37.940 309.925 ;
        RECT 39.150 308.265 42.010 308.645 ;
        RECT 37.560 307.705 37.940 308.085 ;
        RECT 39.150 306.425 42.010 306.805 ;
        RECT 37.560 305.865 37.940 306.245 ;
        RECT 39.150 304.540 42.010 304.920 ;
        RECT 39.150 303.780 42.010 304.160 ;
        RECT 37.560 303.220 37.940 303.600 ;
        RECT 39.150 301.940 42.010 302.320 ;
        RECT 37.560 301.380 37.940 301.760 ;
        RECT 39.150 300.100 42.010 300.480 ;
        RECT 37.560 299.540 37.940 299.920 ;
        RECT 42.785 297.390 44.535 301.200 ;
        RECT 46.625 297.390 48.375 303.040 ;
        RECT 50.465 297.390 52.215 305.685 ;
        RECT 54.305 297.390 56.055 307.525 ;
        RECT 58.145 297.390 59.895 309.365 ;
        RECT 61.985 297.390 63.735 312.010 ;
        RECT 65.825 297.390 67.575 313.850 ;
        RECT 71.600 312.750 74.460 313.130 ;
        RECT 70.010 312.190 70.390 312.570 ;
        RECT 71.600 310.865 74.460 311.245 ;
        RECT 71.600 310.105 74.460 310.485 ;
        RECT 70.010 309.545 70.390 309.925 ;
        RECT 71.600 308.265 74.460 308.645 ;
        RECT 70.010 307.705 70.390 308.085 ;
        RECT 71.600 306.425 74.460 306.805 ;
        RECT 70.010 305.865 70.390 306.245 ;
        RECT 71.600 304.540 74.460 304.920 ;
        RECT 71.600 303.780 74.460 304.160 ;
        RECT 70.010 303.220 70.390 303.600 ;
        RECT 71.600 301.940 74.460 302.320 ;
        RECT 70.010 301.380 70.390 301.760 ;
        RECT 71.600 300.100 74.460 300.480 ;
        RECT 70.010 299.540 70.390 299.920 ;
        RECT 75.235 297.390 76.985 301.200 ;
        RECT 79.075 297.390 80.825 303.040 ;
        RECT 82.915 297.390 84.665 305.685 ;
        RECT 86.755 297.390 88.505 307.525 ;
        RECT 90.595 297.390 92.345 309.365 ;
        RECT 94.435 297.390 96.185 312.010 ;
        RECT 98.275 297.390 100.025 313.850 ;
        RECT 104.050 312.750 106.910 313.130 ;
        RECT 102.460 312.190 102.840 312.570 ;
        RECT 104.050 310.865 106.910 311.245 ;
        RECT 104.050 310.105 106.910 310.485 ;
        RECT 102.460 309.545 102.840 309.925 ;
        RECT 104.050 308.265 106.910 308.645 ;
        RECT 102.460 307.705 102.840 308.085 ;
        RECT 104.050 306.425 106.910 306.805 ;
        RECT 102.460 305.865 102.840 306.245 ;
        RECT 104.050 304.540 106.910 304.920 ;
        RECT 104.050 303.780 106.910 304.160 ;
        RECT 102.460 303.220 102.840 303.600 ;
        RECT 104.050 301.940 106.910 302.320 ;
        RECT 102.460 301.380 102.840 301.760 ;
        RECT 104.050 300.100 106.910 300.480 ;
        RECT 102.460 299.540 102.840 299.920 ;
        RECT 107.685 297.390 109.435 301.200 ;
        RECT 111.525 297.390 113.275 303.040 ;
        RECT 115.365 297.390 117.115 305.685 ;
        RECT 119.205 297.390 120.955 307.525 ;
        RECT 123.045 297.390 124.795 309.365 ;
        RECT 126.885 297.390 128.635 312.010 ;
        RECT 130.725 297.390 132.475 313.850 ;
        RECT 134.910 312.190 135.290 312.570 ;
        RECT 137.355 310.880 137.735 311.260 ;
        RECT 139.395 310.880 139.775 311.260 ;
        RECT 141.180 310.880 141.560 311.260 ;
        RECT 134.910 309.545 135.290 309.925 ;
        RECT 134.910 307.705 135.290 308.085 ;
        RECT 137.355 307.880 137.735 308.260 ;
        RECT 139.395 307.880 139.775 308.260 ;
        RECT 141.180 307.880 141.560 308.260 ;
        RECT 134.910 305.865 135.290 306.245 ;
        RECT 137.355 304.880 137.735 305.260 ;
        RECT 139.395 304.880 139.775 305.260 ;
        RECT 141.180 304.880 141.560 305.260 ;
        RECT 134.910 303.220 135.290 303.600 ;
        RECT 137.355 301.880 137.735 302.260 ;
        RECT 139.395 301.880 139.775 302.260 ;
        RECT 141.180 301.880 141.560 302.260 ;
        RECT 134.910 301.380 135.290 301.760 ;
        RECT 134.910 299.540 135.290 299.920 ;
        RECT 137.355 298.880 137.735 299.260 ;
        RECT 139.395 298.880 139.775 299.260 ;
        RECT 141.180 298.880 141.560 299.260 ;
        RECT 9.100 297.005 9.480 297.195 ;
        RECT 12.940 297.005 13.320 297.195 ;
        RECT 16.780 297.005 17.160 297.195 ;
        RECT 20.620 297.005 21.000 297.195 ;
        RECT 24.460 297.005 24.840 297.195 ;
        RECT 28.300 297.005 28.680 297.195 ;
        RECT 32.140 297.005 32.520 297.195 ;
        RECT 35.980 297.005 36.360 297.195 ;
        RECT 41.550 297.005 41.930 297.195 ;
        RECT 45.390 297.005 45.770 297.195 ;
        RECT 49.230 297.005 49.610 297.195 ;
        RECT 53.070 297.005 53.450 297.195 ;
        RECT 56.910 297.005 57.290 297.195 ;
        RECT 60.750 297.005 61.130 297.195 ;
        RECT 64.590 297.005 64.970 297.195 ;
        RECT 68.430 297.005 68.810 297.195 ;
        RECT 74.000 297.005 74.380 297.195 ;
        RECT 77.840 297.005 78.220 297.195 ;
        RECT 81.680 297.005 82.060 297.195 ;
        RECT 85.520 297.005 85.900 297.195 ;
        RECT 89.360 297.005 89.740 297.195 ;
        RECT 93.200 297.005 93.580 297.195 ;
        RECT 97.040 297.005 97.420 297.195 ;
        RECT 100.880 297.005 101.260 297.195 ;
        RECT 106.450 297.005 106.830 297.195 ;
        RECT 110.290 297.005 110.670 297.195 ;
        RECT 114.130 297.005 114.510 297.195 ;
        RECT 117.970 297.005 118.350 297.195 ;
        RECT 121.810 297.005 122.190 297.195 ;
        RECT 125.650 297.005 126.030 297.195 ;
        RECT 129.490 297.005 129.870 297.195 ;
        RECT 133.330 297.005 133.710 297.195 ;
        RECT 3.430 296.195 141.830 297.005 ;
        RECT 0.240 294.380 0.620 294.760 ;
        RECT 3.430 294.745 4.240 296.195 ;
        RECT 136.340 296.005 136.720 296.195 ;
        RECT 138.380 296.005 138.760 296.195 ;
        RECT 140.420 296.005 140.800 296.195 ;
        RECT 136.340 294.745 136.720 294.935 ;
        RECT 138.380 294.745 138.760 294.935 ;
        RECT 140.420 294.745 140.800 294.935 ;
        RECT 3.430 293.935 141.830 294.745 ;
        RECT 7.180 293.745 7.560 293.935 ;
        RECT 11.020 293.745 11.400 293.935 ;
        RECT 14.860 293.745 15.240 293.935 ;
        RECT 18.700 293.745 19.080 293.935 ;
        RECT 22.540 293.745 22.920 293.935 ;
        RECT 26.380 293.745 26.760 293.935 ;
        RECT 30.220 293.745 30.600 293.935 ;
        RECT 34.060 293.745 34.440 293.935 ;
        RECT 39.630 293.745 40.010 293.935 ;
        RECT 43.470 293.745 43.850 293.935 ;
        RECT 47.310 293.745 47.690 293.935 ;
        RECT 51.150 293.745 51.530 293.935 ;
        RECT 54.990 293.745 55.370 293.935 ;
        RECT 58.830 293.745 59.210 293.935 ;
        RECT 62.670 293.745 63.050 293.935 ;
        RECT 66.510 293.745 66.890 293.935 ;
        RECT 72.080 293.745 72.460 293.935 ;
        RECT 75.920 293.745 76.300 293.935 ;
        RECT 79.760 293.745 80.140 293.935 ;
        RECT 83.600 293.745 83.980 293.935 ;
        RECT 87.440 293.745 87.820 293.935 ;
        RECT 91.280 293.745 91.660 293.935 ;
        RECT 95.120 293.745 95.500 293.935 ;
        RECT 98.960 293.745 99.340 293.935 ;
        RECT 104.530 293.745 104.910 293.935 ;
        RECT 108.370 293.745 108.750 293.935 ;
        RECT 112.210 293.745 112.590 293.935 ;
        RECT 116.050 293.745 116.430 293.935 ;
        RECT 119.890 293.745 120.270 293.935 ;
        RECT 123.730 293.745 124.110 293.935 ;
        RECT 127.570 293.745 127.950 293.935 ;
        RECT 131.410 293.745 131.790 293.935 ;
        RECT 0.240 291.380 0.620 291.760 ;
        RECT 2.520 289.090 2.870 293.280 ;
        RECT 0.240 288.380 0.620 288.760 ;
        RECT 3.150 287.735 3.500 291.650 ;
        RECT 4.160 291.380 4.540 291.760 ;
        RECT 6.700 290.415 9.560 290.795 ;
        RECT 12.255 289.695 14.005 293.550 ;
        RECT 4.160 288.380 4.540 288.760 ;
        RECT 6.700 288.575 9.560 288.955 ;
        RECT 16.095 287.850 17.845 293.550 ;
        RECT 2.745 287.410 3.500 287.735 ;
        RECT 2.300 286.725 2.680 287.105 ;
        RECT 6.700 286.730 9.560 287.110 ;
        RECT 6.700 285.970 9.560 286.350 ;
        RECT 0.240 285.380 0.620 285.760 ;
        RECT 4.160 285.380 4.540 285.760 ;
        RECT 19.935 285.210 21.685 293.550 ;
        RECT 6.700 284.090 9.560 284.470 ;
        RECT 23.775 283.370 25.525 293.550 ;
        RECT 0.240 282.380 0.620 282.760 ;
        RECT 4.160 282.380 4.540 282.760 ;
        RECT 6.700 282.250 9.560 282.630 ;
        RECT 27.615 281.525 29.365 293.550 ;
        RECT 6.700 280.405 9.560 280.785 ;
        RECT 0.240 279.380 0.620 279.760 ;
        RECT 4.160 279.380 4.540 279.760 ;
        RECT 6.700 279.645 9.560 280.025 ;
        RECT 31.455 278.885 33.205 293.550 ;
        RECT 6.700 277.765 9.560 278.145 ;
        RECT 35.295 277.045 37.045 293.550 ;
        RECT 37.560 290.975 37.940 291.355 ;
        RECT 39.150 290.415 42.010 290.795 ;
        RECT 44.705 289.695 46.455 293.550 ;
        RECT 37.560 289.135 37.940 289.515 ;
        RECT 39.150 288.575 42.010 288.955 ;
        RECT 48.545 287.850 50.295 293.550 ;
        RECT 37.560 287.290 37.940 287.670 ;
        RECT 39.150 286.730 42.010 287.110 ;
        RECT 39.150 285.970 42.010 286.350 ;
        RECT 52.385 285.210 54.135 293.550 ;
        RECT 37.560 284.650 37.940 285.030 ;
        RECT 39.150 284.090 42.010 284.470 ;
        RECT 56.225 283.370 57.975 293.550 ;
        RECT 37.560 282.810 37.940 283.190 ;
        RECT 39.150 282.250 42.010 282.630 ;
        RECT 60.065 281.525 61.815 293.550 ;
        RECT 37.560 280.965 37.940 281.345 ;
        RECT 39.150 280.405 42.010 280.785 ;
        RECT 39.150 279.645 42.010 280.025 ;
        RECT 63.905 278.885 65.655 293.550 ;
        RECT 37.560 278.325 37.940 278.705 ;
        RECT 39.150 277.765 42.010 278.145 ;
        RECT 67.745 277.045 69.495 293.550 ;
        RECT 70.010 290.975 70.390 291.355 ;
        RECT 71.600 290.415 74.460 290.795 ;
        RECT 77.155 289.695 78.905 293.550 ;
        RECT 70.010 289.135 70.390 289.515 ;
        RECT 71.600 288.575 74.460 288.955 ;
        RECT 80.995 287.850 82.745 293.550 ;
        RECT 70.010 287.290 70.390 287.670 ;
        RECT 71.600 286.730 74.460 287.110 ;
        RECT 71.600 285.970 74.460 286.350 ;
        RECT 84.835 285.210 86.585 293.550 ;
        RECT 70.010 284.650 70.390 285.030 ;
        RECT 71.600 284.090 74.460 284.470 ;
        RECT 88.675 283.370 90.425 293.550 ;
        RECT 70.010 282.810 70.390 283.190 ;
        RECT 71.600 282.250 74.460 282.630 ;
        RECT 92.515 281.525 94.265 293.550 ;
        RECT 70.010 280.965 70.390 281.345 ;
        RECT 71.600 280.405 74.460 280.785 ;
        RECT 71.600 279.645 74.460 280.025 ;
        RECT 96.355 278.885 98.105 293.550 ;
        RECT 70.010 278.325 70.390 278.705 ;
        RECT 71.600 277.765 74.460 278.145 ;
        RECT 100.195 277.045 101.945 293.550 ;
        RECT 102.460 290.975 102.840 291.355 ;
        RECT 104.050 290.415 106.910 290.795 ;
        RECT 109.605 289.695 111.355 293.550 ;
        RECT 102.460 289.135 102.840 289.515 ;
        RECT 104.050 288.575 106.910 288.955 ;
        RECT 113.445 287.850 115.195 293.550 ;
        RECT 102.460 287.290 102.840 287.670 ;
        RECT 104.050 286.730 106.910 287.110 ;
        RECT 104.050 285.970 106.910 286.350 ;
        RECT 117.285 285.210 119.035 293.550 ;
        RECT 102.460 284.650 102.840 285.030 ;
        RECT 104.050 284.090 106.910 284.470 ;
        RECT 121.125 283.370 122.875 293.550 ;
        RECT 102.460 282.810 102.840 283.190 ;
        RECT 104.050 282.250 106.910 282.630 ;
        RECT 124.965 281.525 126.715 293.550 ;
        RECT 102.460 280.965 102.840 281.345 ;
        RECT 104.050 280.405 106.910 280.785 ;
        RECT 104.050 279.645 106.910 280.025 ;
        RECT 128.805 278.885 130.555 293.550 ;
        RECT 102.460 278.325 102.840 278.705 ;
        RECT 104.050 277.765 106.910 278.145 ;
        RECT 132.645 277.045 134.395 293.550 ;
        RECT 137.355 292.880 137.735 293.260 ;
        RECT 139.395 292.880 139.775 293.260 ;
        RECT 141.180 292.880 141.560 293.260 ;
        RECT 134.910 290.975 135.290 291.355 ;
        RECT 137.355 289.880 137.735 290.260 ;
        RECT 139.395 289.880 139.775 290.260 ;
        RECT 141.180 289.880 141.560 290.260 ;
        RECT 134.910 289.135 135.290 289.515 ;
        RECT 134.910 287.290 135.290 287.670 ;
        RECT 137.355 286.880 137.735 287.260 ;
        RECT 139.395 286.880 139.775 287.260 ;
        RECT 141.180 286.880 141.560 287.260 ;
        RECT 134.910 284.650 135.290 285.030 ;
        RECT 137.355 283.880 137.735 284.260 ;
        RECT 139.395 283.880 139.775 284.260 ;
        RECT 141.180 283.880 141.560 284.260 ;
        RECT 134.910 282.810 135.290 283.190 ;
        RECT 134.910 280.965 135.290 281.345 ;
        RECT 137.355 280.880 137.735 281.260 ;
        RECT 139.395 280.880 139.775 281.260 ;
        RECT 141.180 280.880 141.560 281.260 ;
        RECT 134.910 278.325 135.290 278.705 ;
        RECT 137.355 277.880 137.735 278.260 ;
        RECT 139.395 277.880 139.775 278.260 ;
        RECT 141.180 277.880 141.560 278.260 ;
        RECT 0.240 276.380 0.620 276.760 ;
        RECT 4.160 276.380 4.540 276.760 ;
        RECT 37.560 276.485 37.940 276.865 ;
        RECT 70.010 276.485 70.390 276.865 ;
        RECT 102.460 276.485 102.840 276.865 ;
        RECT 134.910 276.485 135.290 276.865 ;
        RECT 6.700 275.925 9.560 276.305 ;
        RECT 39.150 275.925 42.010 276.305 ;
        RECT 71.600 275.925 74.460 276.305 ;
        RECT 104.050 275.925 106.910 276.305 ;
        RECT 6.700 275.205 9.560 275.585 ;
        RECT 39.150 275.205 42.010 275.585 ;
        RECT 71.600 275.205 74.460 275.585 ;
        RECT 104.050 275.205 106.910 275.585 ;
        RECT 37.560 274.645 37.940 275.025 ;
        RECT 70.010 274.645 70.390 275.025 ;
        RECT 102.460 274.645 102.840 275.025 ;
        RECT 134.910 274.645 135.290 275.025 ;
        RECT 0.240 272.995 0.620 273.375 ;
        RECT 4.160 272.995 4.540 273.375 ;
        RECT 6.700 273.365 9.560 273.745 ;
        RECT 6.700 271.480 9.560 271.860 ;
        RECT 6.700 270.720 9.560 271.100 ;
        RECT 0.240 269.995 0.620 270.375 ;
        RECT 4.160 269.995 4.540 270.375 ;
        RECT 6.700 268.880 9.560 269.260 ;
        RECT 0.240 266.995 0.620 267.375 ;
        RECT 4.160 266.995 4.540 267.375 ;
        RECT 6.700 267.040 9.560 267.420 ;
        RECT 6.700 265.155 9.560 265.535 ;
        RECT 6.700 264.395 9.560 264.775 ;
        RECT 0.240 263.995 0.620 264.375 ;
        RECT 4.160 263.995 4.540 264.375 ;
        RECT 6.700 262.555 9.560 262.935 ;
        RECT 0.240 260.995 0.620 261.375 ;
        RECT 4.160 260.995 4.540 261.375 ;
        RECT 6.700 260.715 9.560 261.095 ;
        RECT 0.240 257.995 0.620 258.375 ;
        RECT 4.160 257.995 4.540 258.375 ;
        RECT 10.335 258.005 12.085 261.815 ;
        RECT 14.175 258.005 15.925 263.655 ;
        RECT 18.015 258.005 19.765 266.300 ;
        RECT 21.855 258.005 23.605 268.140 ;
        RECT 25.695 258.005 27.445 269.980 ;
        RECT 29.535 258.005 31.285 272.625 ;
        RECT 33.375 258.005 35.125 274.465 ;
        RECT 39.150 273.365 42.010 273.745 ;
        RECT 37.560 272.805 37.940 273.185 ;
        RECT 39.150 271.480 42.010 271.860 ;
        RECT 39.150 270.720 42.010 271.100 ;
        RECT 37.560 270.160 37.940 270.540 ;
        RECT 39.150 268.880 42.010 269.260 ;
        RECT 37.560 268.320 37.940 268.700 ;
        RECT 39.150 267.040 42.010 267.420 ;
        RECT 37.560 266.480 37.940 266.860 ;
        RECT 39.150 265.155 42.010 265.535 ;
        RECT 39.150 264.395 42.010 264.775 ;
        RECT 37.560 263.835 37.940 264.215 ;
        RECT 39.150 262.555 42.010 262.935 ;
        RECT 37.560 261.995 37.940 262.375 ;
        RECT 39.150 260.715 42.010 261.095 ;
        RECT 37.560 260.155 37.940 260.535 ;
        RECT 42.785 258.005 44.535 261.815 ;
        RECT 46.625 258.005 48.375 263.655 ;
        RECT 50.465 258.005 52.215 266.300 ;
        RECT 54.305 258.005 56.055 268.140 ;
        RECT 58.145 258.005 59.895 269.980 ;
        RECT 61.985 258.005 63.735 272.625 ;
        RECT 65.825 258.005 67.575 274.465 ;
        RECT 71.600 273.365 74.460 273.745 ;
        RECT 70.010 272.805 70.390 273.185 ;
        RECT 71.600 271.480 74.460 271.860 ;
        RECT 71.600 270.720 74.460 271.100 ;
        RECT 70.010 270.160 70.390 270.540 ;
        RECT 71.600 268.880 74.460 269.260 ;
        RECT 70.010 268.320 70.390 268.700 ;
        RECT 71.600 267.040 74.460 267.420 ;
        RECT 70.010 266.480 70.390 266.860 ;
        RECT 71.600 265.155 74.460 265.535 ;
        RECT 71.600 264.395 74.460 264.775 ;
        RECT 70.010 263.835 70.390 264.215 ;
        RECT 71.600 262.555 74.460 262.935 ;
        RECT 70.010 261.995 70.390 262.375 ;
        RECT 71.600 260.715 74.460 261.095 ;
        RECT 70.010 260.155 70.390 260.535 ;
        RECT 75.235 258.005 76.985 261.815 ;
        RECT 79.075 258.005 80.825 263.655 ;
        RECT 82.915 258.005 84.665 266.300 ;
        RECT 86.755 258.005 88.505 268.140 ;
        RECT 90.595 258.005 92.345 269.980 ;
        RECT 94.435 258.005 96.185 272.625 ;
        RECT 98.275 258.005 100.025 274.465 ;
        RECT 104.050 273.365 106.910 273.745 ;
        RECT 102.460 272.805 102.840 273.185 ;
        RECT 104.050 271.480 106.910 271.860 ;
        RECT 104.050 270.720 106.910 271.100 ;
        RECT 102.460 270.160 102.840 270.540 ;
        RECT 104.050 268.880 106.910 269.260 ;
        RECT 102.460 268.320 102.840 268.700 ;
        RECT 104.050 267.040 106.910 267.420 ;
        RECT 102.460 266.480 102.840 266.860 ;
        RECT 104.050 265.155 106.910 265.535 ;
        RECT 104.050 264.395 106.910 264.775 ;
        RECT 102.460 263.835 102.840 264.215 ;
        RECT 104.050 262.555 106.910 262.935 ;
        RECT 102.460 261.995 102.840 262.375 ;
        RECT 104.050 260.715 106.910 261.095 ;
        RECT 102.460 260.155 102.840 260.535 ;
        RECT 107.685 258.005 109.435 261.815 ;
        RECT 111.525 258.005 113.275 263.655 ;
        RECT 115.365 258.005 117.115 266.300 ;
        RECT 119.205 258.005 120.955 268.140 ;
        RECT 123.045 258.005 124.795 269.980 ;
        RECT 126.885 258.005 128.635 272.625 ;
        RECT 130.725 258.005 132.475 274.465 ;
        RECT 134.910 272.805 135.290 273.185 ;
        RECT 137.355 271.495 137.735 271.875 ;
        RECT 139.395 271.495 139.775 271.875 ;
        RECT 141.180 271.495 141.560 271.875 ;
        RECT 134.910 270.160 135.290 270.540 ;
        RECT 134.910 268.320 135.290 268.700 ;
        RECT 137.355 268.495 137.735 268.875 ;
        RECT 139.395 268.495 139.775 268.875 ;
        RECT 141.180 268.495 141.560 268.875 ;
        RECT 134.910 266.480 135.290 266.860 ;
        RECT 137.355 265.495 137.735 265.875 ;
        RECT 139.395 265.495 139.775 265.875 ;
        RECT 141.180 265.495 141.560 265.875 ;
        RECT 134.910 263.835 135.290 264.215 ;
        RECT 137.355 262.495 137.735 262.875 ;
        RECT 139.395 262.495 139.775 262.875 ;
        RECT 141.180 262.495 141.560 262.875 ;
        RECT 134.910 261.995 135.290 262.375 ;
        RECT 134.910 260.155 135.290 260.535 ;
        RECT 137.355 259.495 137.735 259.875 ;
        RECT 139.395 259.495 139.775 259.875 ;
        RECT 141.180 259.495 141.560 259.875 ;
        RECT 9.100 257.620 9.480 257.810 ;
        RECT 12.940 257.620 13.320 257.810 ;
        RECT 16.780 257.620 17.160 257.810 ;
        RECT 20.620 257.620 21.000 257.810 ;
        RECT 24.460 257.620 24.840 257.810 ;
        RECT 28.300 257.620 28.680 257.810 ;
        RECT 32.140 257.620 32.520 257.810 ;
        RECT 35.980 257.620 36.360 257.810 ;
        RECT 41.550 257.620 41.930 257.810 ;
        RECT 45.390 257.620 45.770 257.810 ;
        RECT 49.230 257.620 49.610 257.810 ;
        RECT 53.070 257.620 53.450 257.810 ;
        RECT 56.910 257.620 57.290 257.810 ;
        RECT 60.750 257.620 61.130 257.810 ;
        RECT 64.590 257.620 64.970 257.810 ;
        RECT 68.430 257.620 68.810 257.810 ;
        RECT 74.000 257.620 74.380 257.810 ;
        RECT 77.840 257.620 78.220 257.810 ;
        RECT 81.680 257.620 82.060 257.810 ;
        RECT 85.520 257.620 85.900 257.810 ;
        RECT 89.360 257.620 89.740 257.810 ;
        RECT 93.200 257.620 93.580 257.810 ;
        RECT 97.040 257.620 97.420 257.810 ;
        RECT 100.880 257.620 101.260 257.810 ;
        RECT 106.450 257.620 106.830 257.810 ;
        RECT 110.290 257.620 110.670 257.810 ;
        RECT 114.130 257.620 114.510 257.810 ;
        RECT 117.970 257.620 118.350 257.810 ;
        RECT 121.810 257.620 122.190 257.810 ;
        RECT 125.650 257.620 126.030 257.810 ;
        RECT 129.490 257.620 129.870 257.810 ;
        RECT 133.330 257.620 133.710 257.810 ;
        RECT 3.430 256.810 141.830 257.620 ;
        RECT 0.240 254.995 0.620 255.375 ;
        RECT 3.430 255.360 4.240 256.810 ;
        RECT 136.340 256.620 136.720 256.810 ;
        RECT 138.380 256.620 138.760 256.810 ;
        RECT 140.420 256.620 140.800 256.810 ;
        RECT 136.340 255.360 136.720 255.550 ;
        RECT 138.380 255.360 138.760 255.550 ;
        RECT 140.420 255.360 140.800 255.550 ;
        RECT 3.430 254.550 141.830 255.360 ;
        RECT 7.180 254.360 7.560 254.550 ;
        RECT 11.020 254.360 11.400 254.550 ;
        RECT 14.860 254.360 15.240 254.550 ;
        RECT 18.700 254.360 19.080 254.550 ;
        RECT 22.540 254.360 22.920 254.550 ;
        RECT 26.380 254.360 26.760 254.550 ;
        RECT 30.220 254.360 30.600 254.550 ;
        RECT 34.060 254.360 34.440 254.550 ;
        RECT 39.630 254.360 40.010 254.550 ;
        RECT 43.470 254.360 43.850 254.550 ;
        RECT 47.310 254.360 47.690 254.550 ;
        RECT 51.150 254.360 51.530 254.550 ;
        RECT 54.990 254.360 55.370 254.550 ;
        RECT 58.830 254.360 59.210 254.550 ;
        RECT 62.670 254.360 63.050 254.550 ;
        RECT 66.510 254.360 66.890 254.550 ;
        RECT 72.080 254.360 72.460 254.550 ;
        RECT 75.920 254.360 76.300 254.550 ;
        RECT 79.760 254.360 80.140 254.550 ;
        RECT 83.600 254.360 83.980 254.550 ;
        RECT 87.440 254.360 87.820 254.550 ;
        RECT 91.280 254.360 91.660 254.550 ;
        RECT 95.120 254.360 95.500 254.550 ;
        RECT 98.960 254.360 99.340 254.550 ;
        RECT 104.530 254.360 104.910 254.550 ;
        RECT 108.370 254.360 108.750 254.550 ;
        RECT 112.210 254.360 112.590 254.550 ;
        RECT 116.050 254.360 116.430 254.550 ;
        RECT 119.890 254.360 120.270 254.550 ;
        RECT 123.730 254.360 124.110 254.550 ;
        RECT 127.570 254.360 127.950 254.550 ;
        RECT 131.410 254.360 131.790 254.550 ;
        RECT 0.240 251.995 0.620 252.375 ;
        RECT 2.520 249.705 2.870 253.895 ;
        RECT 0.240 248.995 0.620 249.375 ;
        RECT 3.150 248.350 3.500 252.265 ;
        RECT 4.160 251.995 4.540 252.375 ;
        RECT 6.700 251.030 9.560 251.410 ;
        RECT 12.255 250.310 14.005 254.165 ;
        RECT 4.160 248.995 4.540 249.375 ;
        RECT 6.700 249.190 9.560 249.570 ;
        RECT 16.095 248.465 17.845 254.165 ;
        RECT 2.745 248.025 3.500 248.350 ;
        RECT 2.300 247.340 2.680 247.720 ;
        RECT 6.700 247.345 9.560 247.725 ;
        RECT 6.700 246.585 9.560 246.965 ;
        RECT 0.240 245.995 0.620 246.375 ;
        RECT 4.160 245.995 4.540 246.375 ;
        RECT 19.935 245.825 21.685 254.165 ;
        RECT 6.700 244.705 9.560 245.085 ;
        RECT 23.775 243.985 25.525 254.165 ;
        RECT 0.240 242.995 0.620 243.375 ;
        RECT 4.160 242.995 4.540 243.375 ;
        RECT 6.700 242.865 9.560 243.245 ;
        RECT 27.615 242.140 29.365 254.165 ;
        RECT 6.700 241.020 9.560 241.400 ;
        RECT 0.240 239.995 0.620 240.375 ;
        RECT 4.160 239.995 4.540 240.375 ;
        RECT 6.700 240.260 9.560 240.640 ;
        RECT 31.455 239.500 33.205 254.165 ;
        RECT 6.700 238.380 9.560 238.760 ;
        RECT 35.295 237.660 37.045 254.165 ;
        RECT 37.560 251.590 37.940 251.970 ;
        RECT 39.150 251.030 42.010 251.410 ;
        RECT 44.705 250.310 46.455 254.165 ;
        RECT 37.560 249.750 37.940 250.130 ;
        RECT 39.150 249.190 42.010 249.570 ;
        RECT 48.545 248.465 50.295 254.165 ;
        RECT 37.560 247.905 37.940 248.285 ;
        RECT 39.150 247.345 42.010 247.725 ;
        RECT 39.150 246.585 42.010 246.965 ;
        RECT 52.385 245.825 54.135 254.165 ;
        RECT 37.560 245.265 37.940 245.645 ;
        RECT 39.150 244.705 42.010 245.085 ;
        RECT 56.225 243.985 57.975 254.165 ;
        RECT 37.560 243.425 37.940 243.805 ;
        RECT 39.150 242.865 42.010 243.245 ;
        RECT 60.065 242.140 61.815 254.165 ;
        RECT 37.560 241.580 37.940 241.960 ;
        RECT 39.150 241.020 42.010 241.400 ;
        RECT 39.150 240.260 42.010 240.640 ;
        RECT 63.905 239.500 65.655 254.165 ;
        RECT 37.560 238.940 37.940 239.320 ;
        RECT 39.150 238.380 42.010 238.760 ;
        RECT 67.745 237.660 69.495 254.165 ;
        RECT 70.010 251.590 70.390 251.970 ;
        RECT 71.600 251.030 74.460 251.410 ;
        RECT 77.155 250.310 78.905 254.165 ;
        RECT 70.010 249.750 70.390 250.130 ;
        RECT 71.600 249.190 74.460 249.570 ;
        RECT 80.995 248.465 82.745 254.165 ;
        RECT 70.010 247.905 70.390 248.285 ;
        RECT 71.600 247.345 74.460 247.725 ;
        RECT 71.600 246.585 74.460 246.965 ;
        RECT 84.835 245.825 86.585 254.165 ;
        RECT 70.010 245.265 70.390 245.645 ;
        RECT 71.600 244.705 74.460 245.085 ;
        RECT 88.675 243.985 90.425 254.165 ;
        RECT 70.010 243.425 70.390 243.805 ;
        RECT 71.600 242.865 74.460 243.245 ;
        RECT 92.515 242.140 94.265 254.165 ;
        RECT 70.010 241.580 70.390 241.960 ;
        RECT 71.600 241.020 74.460 241.400 ;
        RECT 71.600 240.260 74.460 240.640 ;
        RECT 96.355 239.500 98.105 254.165 ;
        RECT 70.010 238.940 70.390 239.320 ;
        RECT 71.600 238.380 74.460 238.760 ;
        RECT 100.195 237.660 101.945 254.165 ;
        RECT 102.460 251.590 102.840 251.970 ;
        RECT 104.050 251.030 106.910 251.410 ;
        RECT 109.605 250.310 111.355 254.165 ;
        RECT 102.460 249.750 102.840 250.130 ;
        RECT 104.050 249.190 106.910 249.570 ;
        RECT 113.445 248.465 115.195 254.165 ;
        RECT 102.460 247.905 102.840 248.285 ;
        RECT 104.050 247.345 106.910 247.725 ;
        RECT 104.050 246.585 106.910 246.965 ;
        RECT 117.285 245.825 119.035 254.165 ;
        RECT 102.460 245.265 102.840 245.645 ;
        RECT 104.050 244.705 106.910 245.085 ;
        RECT 121.125 243.985 122.875 254.165 ;
        RECT 102.460 243.425 102.840 243.805 ;
        RECT 104.050 242.865 106.910 243.245 ;
        RECT 124.965 242.140 126.715 254.165 ;
        RECT 102.460 241.580 102.840 241.960 ;
        RECT 104.050 241.020 106.910 241.400 ;
        RECT 104.050 240.260 106.910 240.640 ;
        RECT 128.805 239.500 130.555 254.165 ;
        RECT 102.460 238.940 102.840 239.320 ;
        RECT 104.050 238.380 106.910 238.760 ;
        RECT 132.645 237.660 134.395 254.165 ;
        RECT 137.355 253.495 137.735 253.875 ;
        RECT 139.395 253.495 139.775 253.875 ;
        RECT 141.180 253.495 141.560 253.875 ;
        RECT 134.910 251.590 135.290 251.970 ;
        RECT 137.355 250.495 137.735 250.875 ;
        RECT 139.395 250.495 139.775 250.875 ;
        RECT 141.180 250.495 141.560 250.875 ;
        RECT 134.910 249.750 135.290 250.130 ;
        RECT 134.910 247.905 135.290 248.285 ;
        RECT 137.355 247.495 137.735 247.875 ;
        RECT 139.395 247.495 139.775 247.875 ;
        RECT 141.180 247.495 141.560 247.875 ;
        RECT 134.910 245.265 135.290 245.645 ;
        RECT 137.355 244.495 137.735 244.875 ;
        RECT 139.395 244.495 139.775 244.875 ;
        RECT 141.180 244.495 141.560 244.875 ;
        RECT 134.910 243.425 135.290 243.805 ;
        RECT 134.910 241.580 135.290 241.960 ;
        RECT 137.355 241.495 137.735 241.875 ;
        RECT 139.395 241.495 139.775 241.875 ;
        RECT 141.180 241.495 141.560 241.875 ;
        RECT 134.910 238.940 135.290 239.320 ;
        RECT 137.355 238.495 137.735 238.875 ;
        RECT 139.395 238.495 139.775 238.875 ;
        RECT 141.180 238.495 141.560 238.875 ;
        RECT 0.240 236.995 0.620 237.375 ;
        RECT 4.160 236.995 4.540 237.375 ;
        RECT 37.560 237.100 37.940 237.480 ;
        RECT 70.010 237.100 70.390 237.480 ;
        RECT 102.460 237.100 102.840 237.480 ;
        RECT 134.910 237.100 135.290 237.480 ;
        RECT 6.700 236.540 9.560 236.920 ;
        RECT 39.150 236.540 42.010 236.920 ;
        RECT 71.600 236.540 74.460 236.920 ;
        RECT 104.050 236.540 106.910 236.920 ;
        RECT 6.700 235.820 9.560 236.200 ;
        RECT 39.150 235.820 42.010 236.200 ;
        RECT 71.600 235.820 74.460 236.200 ;
        RECT 104.050 235.820 106.910 236.200 ;
        RECT 37.560 235.260 37.940 235.640 ;
        RECT 70.010 235.260 70.390 235.640 ;
        RECT 102.460 235.260 102.840 235.640 ;
        RECT 134.910 235.260 135.290 235.640 ;
        RECT 0.240 233.610 0.620 233.990 ;
        RECT 4.160 233.610 4.540 233.990 ;
        RECT 6.700 233.980 9.560 234.360 ;
        RECT 6.700 232.095 9.560 232.475 ;
        RECT 6.700 231.335 9.560 231.715 ;
        RECT 0.240 230.610 0.620 230.990 ;
        RECT 4.160 230.610 4.540 230.990 ;
        RECT 6.700 229.495 9.560 229.875 ;
        RECT 0.240 227.610 0.620 227.990 ;
        RECT 4.160 227.610 4.540 227.990 ;
        RECT 6.700 227.655 9.560 228.035 ;
        RECT 6.700 225.770 9.560 226.150 ;
        RECT 6.700 225.010 9.560 225.390 ;
        RECT 0.240 224.610 0.620 224.990 ;
        RECT 4.160 224.610 4.540 224.990 ;
        RECT 6.700 223.170 9.560 223.550 ;
        RECT 0.240 221.610 0.620 221.990 ;
        RECT 4.160 221.610 4.540 221.990 ;
        RECT 6.700 221.330 9.560 221.710 ;
        RECT 0.240 218.610 0.620 218.990 ;
        RECT 4.160 218.610 4.540 218.990 ;
        RECT 10.335 218.620 12.085 222.430 ;
        RECT 14.175 218.620 15.925 224.270 ;
        RECT 18.015 218.620 19.765 226.915 ;
        RECT 21.855 218.620 23.605 228.755 ;
        RECT 25.695 218.620 27.445 230.595 ;
        RECT 29.535 218.620 31.285 233.240 ;
        RECT 33.375 218.620 35.125 235.080 ;
        RECT 39.150 233.980 42.010 234.360 ;
        RECT 37.560 233.420 37.940 233.800 ;
        RECT 39.150 232.095 42.010 232.475 ;
        RECT 39.150 231.335 42.010 231.715 ;
        RECT 37.560 230.775 37.940 231.155 ;
        RECT 39.150 229.495 42.010 229.875 ;
        RECT 37.560 228.935 37.940 229.315 ;
        RECT 39.150 227.655 42.010 228.035 ;
        RECT 37.560 227.095 37.940 227.475 ;
        RECT 39.150 225.770 42.010 226.150 ;
        RECT 39.150 225.010 42.010 225.390 ;
        RECT 37.560 224.450 37.940 224.830 ;
        RECT 39.150 223.170 42.010 223.550 ;
        RECT 37.560 222.610 37.940 222.990 ;
        RECT 39.150 221.330 42.010 221.710 ;
        RECT 37.560 220.770 37.940 221.150 ;
        RECT 42.785 218.620 44.535 222.430 ;
        RECT 46.625 218.620 48.375 224.270 ;
        RECT 50.465 218.620 52.215 226.915 ;
        RECT 54.305 218.620 56.055 228.755 ;
        RECT 58.145 218.620 59.895 230.595 ;
        RECT 61.985 218.620 63.735 233.240 ;
        RECT 65.825 218.620 67.575 235.080 ;
        RECT 71.600 233.980 74.460 234.360 ;
        RECT 70.010 233.420 70.390 233.800 ;
        RECT 71.600 232.095 74.460 232.475 ;
        RECT 71.600 231.335 74.460 231.715 ;
        RECT 70.010 230.775 70.390 231.155 ;
        RECT 71.600 229.495 74.460 229.875 ;
        RECT 70.010 228.935 70.390 229.315 ;
        RECT 71.600 227.655 74.460 228.035 ;
        RECT 70.010 227.095 70.390 227.475 ;
        RECT 71.600 225.770 74.460 226.150 ;
        RECT 71.600 225.010 74.460 225.390 ;
        RECT 70.010 224.450 70.390 224.830 ;
        RECT 71.600 223.170 74.460 223.550 ;
        RECT 70.010 222.610 70.390 222.990 ;
        RECT 71.600 221.330 74.460 221.710 ;
        RECT 70.010 220.770 70.390 221.150 ;
        RECT 75.235 218.620 76.985 222.430 ;
        RECT 79.075 218.620 80.825 224.270 ;
        RECT 82.915 218.620 84.665 226.915 ;
        RECT 86.755 218.620 88.505 228.755 ;
        RECT 90.595 218.620 92.345 230.595 ;
        RECT 94.435 218.620 96.185 233.240 ;
        RECT 98.275 218.620 100.025 235.080 ;
        RECT 104.050 233.980 106.910 234.360 ;
        RECT 102.460 233.420 102.840 233.800 ;
        RECT 104.050 232.095 106.910 232.475 ;
        RECT 104.050 231.335 106.910 231.715 ;
        RECT 102.460 230.775 102.840 231.155 ;
        RECT 104.050 229.495 106.910 229.875 ;
        RECT 102.460 228.935 102.840 229.315 ;
        RECT 104.050 227.655 106.910 228.035 ;
        RECT 102.460 227.095 102.840 227.475 ;
        RECT 104.050 225.770 106.910 226.150 ;
        RECT 104.050 225.010 106.910 225.390 ;
        RECT 102.460 224.450 102.840 224.830 ;
        RECT 104.050 223.170 106.910 223.550 ;
        RECT 102.460 222.610 102.840 222.990 ;
        RECT 104.050 221.330 106.910 221.710 ;
        RECT 102.460 220.770 102.840 221.150 ;
        RECT 107.685 218.620 109.435 222.430 ;
        RECT 111.525 218.620 113.275 224.270 ;
        RECT 115.365 218.620 117.115 226.915 ;
        RECT 119.205 218.620 120.955 228.755 ;
        RECT 123.045 218.620 124.795 230.595 ;
        RECT 126.885 218.620 128.635 233.240 ;
        RECT 130.725 218.620 132.475 235.080 ;
        RECT 134.910 233.420 135.290 233.800 ;
        RECT 137.355 232.110 137.735 232.490 ;
        RECT 139.395 232.110 139.775 232.490 ;
        RECT 141.180 232.110 141.560 232.490 ;
        RECT 134.910 230.775 135.290 231.155 ;
        RECT 134.910 228.935 135.290 229.315 ;
        RECT 137.355 229.110 137.735 229.490 ;
        RECT 139.395 229.110 139.775 229.490 ;
        RECT 141.180 229.110 141.560 229.490 ;
        RECT 134.910 227.095 135.290 227.475 ;
        RECT 137.355 226.110 137.735 226.490 ;
        RECT 139.395 226.110 139.775 226.490 ;
        RECT 141.180 226.110 141.560 226.490 ;
        RECT 134.910 224.450 135.290 224.830 ;
        RECT 137.355 223.110 137.735 223.490 ;
        RECT 139.395 223.110 139.775 223.490 ;
        RECT 141.180 223.110 141.560 223.490 ;
        RECT 134.910 222.610 135.290 222.990 ;
        RECT 134.910 220.770 135.290 221.150 ;
        RECT 137.355 220.110 137.735 220.490 ;
        RECT 139.395 220.110 139.775 220.490 ;
        RECT 141.180 220.110 141.560 220.490 ;
        RECT 9.100 218.235 9.480 218.425 ;
        RECT 12.940 218.235 13.320 218.425 ;
        RECT 16.780 218.235 17.160 218.425 ;
        RECT 20.620 218.235 21.000 218.425 ;
        RECT 24.460 218.235 24.840 218.425 ;
        RECT 28.300 218.235 28.680 218.425 ;
        RECT 32.140 218.235 32.520 218.425 ;
        RECT 35.980 218.235 36.360 218.425 ;
        RECT 41.550 218.235 41.930 218.425 ;
        RECT 45.390 218.235 45.770 218.425 ;
        RECT 49.230 218.235 49.610 218.425 ;
        RECT 53.070 218.235 53.450 218.425 ;
        RECT 56.910 218.235 57.290 218.425 ;
        RECT 60.750 218.235 61.130 218.425 ;
        RECT 64.590 218.235 64.970 218.425 ;
        RECT 68.430 218.235 68.810 218.425 ;
        RECT 74.000 218.235 74.380 218.425 ;
        RECT 77.840 218.235 78.220 218.425 ;
        RECT 81.680 218.235 82.060 218.425 ;
        RECT 85.520 218.235 85.900 218.425 ;
        RECT 89.360 218.235 89.740 218.425 ;
        RECT 93.200 218.235 93.580 218.425 ;
        RECT 97.040 218.235 97.420 218.425 ;
        RECT 100.880 218.235 101.260 218.425 ;
        RECT 106.450 218.235 106.830 218.425 ;
        RECT 110.290 218.235 110.670 218.425 ;
        RECT 114.130 218.235 114.510 218.425 ;
        RECT 117.970 218.235 118.350 218.425 ;
        RECT 121.810 218.235 122.190 218.425 ;
        RECT 125.650 218.235 126.030 218.425 ;
        RECT 129.490 218.235 129.870 218.425 ;
        RECT 133.330 218.235 133.710 218.425 ;
        RECT 3.430 217.425 141.830 218.235 ;
        RECT 0.240 215.610 0.620 215.990 ;
        RECT 3.430 215.975 4.240 217.425 ;
        RECT 136.340 217.235 136.720 217.425 ;
        RECT 138.380 217.235 138.760 217.425 ;
        RECT 140.420 217.235 140.800 217.425 ;
        RECT 136.340 215.975 136.720 216.165 ;
        RECT 138.380 215.975 138.760 216.165 ;
        RECT 140.420 215.975 140.800 216.165 ;
        RECT 3.430 215.165 141.830 215.975 ;
        RECT 7.180 214.975 7.560 215.165 ;
        RECT 11.020 214.975 11.400 215.165 ;
        RECT 14.860 214.975 15.240 215.165 ;
        RECT 18.700 214.975 19.080 215.165 ;
        RECT 22.540 214.975 22.920 215.165 ;
        RECT 26.380 214.975 26.760 215.165 ;
        RECT 30.220 214.975 30.600 215.165 ;
        RECT 34.060 214.975 34.440 215.165 ;
        RECT 39.630 214.975 40.010 215.165 ;
        RECT 43.470 214.975 43.850 215.165 ;
        RECT 47.310 214.975 47.690 215.165 ;
        RECT 51.150 214.975 51.530 215.165 ;
        RECT 54.990 214.975 55.370 215.165 ;
        RECT 58.830 214.975 59.210 215.165 ;
        RECT 62.670 214.975 63.050 215.165 ;
        RECT 66.510 214.975 66.890 215.165 ;
        RECT 72.080 214.975 72.460 215.165 ;
        RECT 75.920 214.975 76.300 215.165 ;
        RECT 79.760 214.975 80.140 215.165 ;
        RECT 83.600 214.975 83.980 215.165 ;
        RECT 87.440 214.975 87.820 215.165 ;
        RECT 91.280 214.975 91.660 215.165 ;
        RECT 95.120 214.975 95.500 215.165 ;
        RECT 98.960 214.975 99.340 215.165 ;
        RECT 104.530 214.975 104.910 215.165 ;
        RECT 108.370 214.975 108.750 215.165 ;
        RECT 112.210 214.975 112.590 215.165 ;
        RECT 116.050 214.975 116.430 215.165 ;
        RECT 119.890 214.975 120.270 215.165 ;
        RECT 123.730 214.975 124.110 215.165 ;
        RECT 127.570 214.975 127.950 215.165 ;
        RECT 131.410 214.975 131.790 215.165 ;
        RECT 0.240 212.610 0.620 212.990 ;
        RECT 2.520 210.320 2.870 214.510 ;
        RECT 0.240 209.610 0.620 209.990 ;
        RECT 3.150 208.965 3.500 212.880 ;
        RECT 4.160 212.610 4.540 212.990 ;
        RECT 6.700 211.645 9.560 212.025 ;
        RECT 12.255 210.925 14.005 214.780 ;
        RECT 4.160 209.610 4.540 209.990 ;
        RECT 6.700 209.805 9.560 210.185 ;
        RECT 16.095 209.080 17.845 214.780 ;
        RECT 2.745 208.640 3.500 208.965 ;
        RECT 2.300 207.955 2.680 208.335 ;
        RECT 6.700 207.960 9.560 208.340 ;
        RECT 6.700 207.200 9.560 207.580 ;
        RECT 0.240 206.610 0.620 206.990 ;
        RECT 4.160 206.610 4.540 206.990 ;
        RECT 19.935 206.440 21.685 214.780 ;
        RECT 6.700 205.320 9.560 205.700 ;
        RECT 23.775 204.600 25.525 214.780 ;
        RECT 0.240 203.610 0.620 203.990 ;
        RECT 4.160 203.610 4.540 203.990 ;
        RECT 6.700 203.480 9.560 203.860 ;
        RECT 27.615 202.755 29.365 214.780 ;
        RECT 6.700 201.635 9.560 202.015 ;
        RECT 0.240 200.610 0.620 200.990 ;
        RECT 4.160 200.610 4.540 200.990 ;
        RECT 6.700 200.875 9.560 201.255 ;
        RECT 31.455 200.115 33.205 214.780 ;
        RECT 6.700 198.995 9.560 199.375 ;
        RECT 35.295 198.275 37.045 214.780 ;
        RECT 37.560 212.205 37.940 212.585 ;
        RECT 39.150 211.645 42.010 212.025 ;
        RECT 44.705 210.925 46.455 214.780 ;
        RECT 37.560 210.365 37.940 210.745 ;
        RECT 39.150 209.805 42.010 210.185 ;
        RECT 48.545 209.080 50.295 214.780 ;
        RECT 37.560 208.520 37.940 208.900 ;
        RECT 39.150 207.960 42.010 208.340 ;
        RECT 39.150 207.200 42.010 207.580 ;
        RECT 52.385 206.440 54.135 214.780 ;
        RECT 37.560 205.880 37.940 206.260 ;
        RECT 39.150 205.320 42.010 205.700 ;
        RECT 56.225 204.600 57.975 214.780 ;
        RECT 37.560 204.040 37.940 204.420 ;
        RECT 39.150 203.480 42.010 203.860 ;
        RECT 60.065 202.755 61.815 214.780 ;
        RECT 37.560 202.195 37.940 202.575 ;
        RECT 39.150 201.635 42.010 202.015 ;
        RECT 39.150 200.875 42.010 201.255 ;
        RECT 63.905 200.115 65.655 214.780 ;
        RECT 37.560 199.555 37.940 199.935 ;
        RECT 39.150 198.995 42.010 199.375 ;
        RECT 67.745 198.275 69.495 214.780 ;
        RECT 70.010 212.205 70.390 212.585 ;
        RECT 71.600 211.645 74.460 212.025 ;
        RECT 77.155 210.925 78.905 214.780 ;
        RECT 70.010 210.365 70.390 210.745 ;
        RECT 71.600 209.805 74.460 210.185 ;
        RECT 80.995 209.080 82.745 214.780 ;
        RECT 70.010 208.520 70.390 208.900 ;
        RECT 71.600 207.960 74.460 208.340 ;
        RECT 71.600 207.200 74.460 207.580 ;
        RECT 84.835 206.440 86.585 214.780 ;
        RECT 70.010 205.880 70.390 206.260 ;
        RECT 71.600 205.320 74.460 205.700 ;
        RECT 88.675 204.600 90.425 214.780 ;
        RECT 70.010 204.040 70.390 204.420 ;
        RECT 71.600 203.480 74.460 203.860 ;
        RECT 92.515 202.755 94.265 214.780 ;
        RECT 70.010 202.195 70.390 202.575 ;
        RECT 71.600 201.635 74.460 202.015 ;
        RECT 71.600 200.875 74.460 201.255 ;
        RECT 96.355 200.115 98.105 214.780 ;
        RECT 70.010 199.555 70.390 199.935 ;
        RECT 71.600 198.995 74.460 199.375 ;
        RECT 100.195 198.275 101.945 214.780 ;
        RECT 102.460 212.205 102.840 212.585 ;
        RECT 104.050 211.645 106.910 212.025 ;
        RECT 109.605 210.925 111.355 214.780 ;
        RECT 102.460 210.365 102.840 210.745 ;
        RECT 104.050 209.805 106.910 210.185 ;
        RECT 113.445 209.080 115.195 214.780 ;
        RECT 102.460 208.520 102.840 208.900 ;
        RECT 104.050 207.960 106.910 208.340 ;
        RECT 104.050 207.200 106.910 207.580 ;
        RECT 117.285 206.440 119.035 214.780 ;
        RECT 102.460 205.880 102.840 206.260 ;
        RECT 104.050 205.320 106.910 205.700 ;
        RECT 121.125 204.600 122.875 214.780 ;
        RECT 102.460 204.040 102.840 204.420 ;
        RECT 104.050 203.480 106.910 203.860 ;
        RECT 124.965 202.755 126.715 214.780 ;
        RECT 102.460 202.195 102.840 202.575 ;
        RECT 104.050 201.635 106.910 202.015 ;
        RECT 104.050 200.875 106.910 201.255 ;
        RECT 128.805 200.115 130.555 214.780 ;
        RECT 102.460 199.555 102.840 199.935 ;
        RECT 104.050 198.995 106.910 199.375 ;
        RECT 132.645 198.275 134.395 214.780 ;
        RECT 137.355 214.110 137.735 214.490 ;
        RECT 139.395 214.110 139.775 214.490 ;
        RECT 141.180 214.110 141.560 214.490 ;
        RECT 134.910 212.205 135.290 212.585 ;
        RECT 137.355 211.110 137.735 211.490 ;
        RECT 139.395 211.110 139.775 211.490 ;
        RECT 141.180 211.110 141.560 211.490 ;
        RECT 134.910 210.365 135.290 210.745 ;
        RECT 134.910 208.520 135.290 208.900 ;
        RECT 137.355 208.110 137.735 208.490 ;
        RECT 139.395 208.110 139.775 208.490 ;
        RECT 141.180 208.110 141.560 208.490 ;
        RECT 134.910 205.880 135.290 206.260 ;
        RECT 137.355 205.110 137.735 205.490 ;
        RECT 139.395 205.110 139.775 205.490 ;
        RECT 141.180 205.110 141.560 205.490 ;
        RECT 134.910 204.040 135.290 204.420 ;
        RECT 134.910 202.195 135.290 202.575 ;
        RECT 137.355 202.110 137.735 202.490 ;
        RECT 139.395 202.110 139.775 202.490 ;
        RECT 141.180 202.110 141.560 202.490 ;
        RECT 134.910 199.555 135.290 199.935 ;
        RECT 137.355 199.110 137.735 199.490 ;
        RECT 139.395 199.110 139.775 199.490 ;
        RECT 141.180 199.110 141.560 199.490 ;
        RECT 0.240 197.610 0.620 197.990 ;
        RECT 4.160 197.610 4.540 197.990 ;
        RECT 37.560 197.715 37.940 198.095 ;
        RECT 70.010 197.715 70.390 198.095 ;
        RECT 102.460 197.715 102.840 198.095 ;
        RECT 134.910 197.715 135.290 198.095 ;
        RECT 6.700 197.155 9.560 197.535 ;
        RECT 39.150 197.155 42.010 197.535 ;
        RECT 71.600 197.155 74.460 197.535 ;
        RECT 104.050 197.155 106.910 197.535 ;
        RECT 6.700 196.435 9.560 196.815 ;
        RECT 39.150 196.435 42.010 196.815 ;
        RECT 71.600 196.435 74.460 196.815 ;
        RECT 104.050 196.435 106.910 196.815 ;
        RECT 37.560 195.875 37.940 196.255 ;
        RECT 70.010 195.875 70.390 196.255 ;
        RECT 102.460 195.875 102.840 196.255 ;
        RECT 134.910 195.875 135.290 196.255 ;
        RECT 0.240 194.225 0.620 194.605 ;
        RECT 4.160 194.225 4.540 194.605 ;
        RECT 6.700 194.595 9.560 194.975 ;
        RECT 6.700 192.710 9.560 193.090 ;
        RECT 6.700 191.950 9.560 192.330 ;
        RECT 0.240 191.225 0.620 191.605 ;
        RECT 4.160 191.225 4.540 191.605 ;
        RECT 6.700 190.110 9.560 190.490 ;
        RECT 0.240 188.225 0.620 188.605 ;
        RECT 4.160 188.225 4.540 188.605 ;
        RECT 6.700 188.270 9.560 188.650 ;
        RECT 6.700 186.385 9.560 186.765 ;
        RECT 6.700 185.625 9.560 186.005 ;
        RECT 0.240 185.225 0.620 185.605 ;
        RECT 4.160 185.225 4.540 185.605 ;
        RECT 6.700 183.785 9.560 184.165 ;
        RECT 0.240 182.225 0.620 182.605 ;
        RECT 4.160 182.225 4.540 182.605 ;
        RECT 6.700 181.945 9.560 182.325 ;
        RECT 0.240 179.225 0.620 179.605 ;
        RECT 4.160 179.225 4.540 179.605 ;
        RECT 10.335 179.235 12.085 183.045 ;
        RECT 14.175 179.235 15.925 184.885 ;
        RECT 18.015 179.235 19.765 187.530 ;
        RECT 21.855 179.235 23.605 189.370 ;
        RECT 25.695 179.235 27.445 191.210 ;
        RECT 29.535 179.235 31.285 193.855 ;
        RECT 33.375 179.235 35.125 195.695 ;
        RECT 39.150 194.595 42.010 194.975 ;
        RECT 37.560 194.035 37.940 194.415 ;
        RECT 39.150 192.710 42.010 193.090 ;
        RECT 39.150 191.950 42.010 192.330 ;
        RECT 37.560 191.390 37.940 191.770 ;
        RECT 39.150 190.110 42.010 190.490 ;
        RECT 37.560 189.550 37.940 189.930 ;
        RECT 39.150 188.270 42.010 188.650 ;
        RECT 37.560 187.710 37.940 188.090 ;
        RECT 39.150 186.385 42.010 186.765 ;
        RECT 39.150 185.625 42.010 186.005 ;
        RECT 37.560 185.065 37.940 185.445 ;
        RECT 39.150 183.785 42.010 184.165 ;
        RECT 37.560 183.225 37.940 183.605 ;
        RECT 39.150 181.945 42.010 182.325 ;
        RECT 37.560 181.385 37.940 181.765 ;
        RECT 42.785 179.235 44.535 183.045 ;
        RECT 46.625 179.235 48.375 184.885 ;
        RECT 50.465 179.235 52.215 187.530 ;
        RECT 54.305 179.235 56.055 189.370 ;
        RECT 58.145 179.235 59.895 191.210 ;
        RECT 61.985 179.235 63.735 193.855 ;
        RECT 65.825 179.235 67.575 195.695 ;
        RECT 71.600 194.595 74.460 194.975 ;
        RECT 70.010 194.035 70.390 194.415 ;
        RECT 71.600 192.710 74.460 193.090 ;
        RECT 71.600 191.950 74.460 192.330 ;
        RECT 70.010 191.390 70.390 191.770 ;
        RECT 71.600 190.110 74.460 190.490 ;
        RECT 70.010 189.550 70.390 189.930 ;
        RECT 71.600 188.270 74.460 188.650 ;
        RECT 70.010 187.710 70.390 188.090 ;
        RECT 71.600 186.385 74.460 186.765 ;
        RECT 71.600 185.625 74.460 186.005 ;
        RECT 70.010 185.065 70.390 185.445 ;
        RECT 71.600 183.785 74.460 184.165 ;
        RECT 70.010 183.225 70.390 183.605 ;
        RECT 71.600 181.945 74.460 182.325 ;
        RECT 70.010 181.385 70.390 181.765 ;
        RECT 75.235 179.235 76.985 183.045 ;
        RECT 79.075 179.235 80.825 184.885 ;
        RECT 82.915 179.235 84.665 187.530 ;
        RECT 86.755 179.235 88.505 189.370 ;
        RECT 90.595 179.235 92.345 191.210 ;
        RECT 94.435 179.235 96.185 193.855 ;
        RECT 98.275 179.235 100.025 195.695 ;
        RECT 104.050 194.595 106.910 194.975 ;
        RECT 102.460 194.035 102.840 194.415 ;
        RECT 104.050 192.710 106.910 193.090 ;
        RECT 104.050 191.950 106.910 192.330 ;
        RECT 102.460 191.390 102.840 191.770 ;
        RECT 104.050 190.110 106.910 190.490 ;
        RECT 102.460 189.550 102.840 189.930 ;
        RECT 104.050 188.270 106.910 188.650 ;
        RECT 102.460 187.710 102.840 188.090 ;
        RECT 104.050 186.385 106.910 186.765 ;
        RECT 104.050 185.625 106.910 186.005 ;
        RECT 102.460 185.065 102.840 185.445 ;
        RECT 104.050 183.785 106.910 184.165 ;
        RECT 102.460 183.225 102.840 183.605 ;
        RECT 104.050 181.945 106.910 182.325 ;
        RECT 102.460 181.385 102.840 181.765 ;
        RECT 107.685 179.235 109.435 183.045 ;
        RECT 111.525 179.235 113.275 184.885 ;
        RECT 115.365 179.235 117.115 187.530 ;
        RECT 119.205 179.235 120.955 189.370 ;
        RECT 123.045 179.235 124.795 191.210 ;
        RECT 126.885 179.235 128.635 193.855 ;
        RECT 130.725 179.235 132.475 195.695 ;
        RECT 134.910 194.035 135.290 194.415 ;
        RECT 137.355 192.725 137.735 193.105 ;
        RECT 139.395 192.725 139.775 193.105 ;
        RECT 141.180 192.725 141.560 193.105 ;
        RECT 134.910 191.390 135.290 191.770 ;
        RECT 134.910 189.550 135.290 189.930 ;
        RECT 137.355 189.725 137.735 190.105 ;
        RECT 139.395 189.725 139.775 190.105 ;
        RECT 141.180 189.725 141.560 190.105 ;
        RECT 134.910 187.710 135.290 188.090 ;
        RECT 137.355 186.725 137.735 187.105 ;
        RECT 139.395 186.725 139.775 187.105 ;
        RECT 141.180 186.725 141.560 187.105 ;
        RECT 134.910 185.065 135.290 185.445 ;
        RECT 137.355 183.725 137.735 184.105 ;
        RECT 139.395 183.725 139.775 184.105 ;
        RECT 141.180 183.725 141.560 184.105 ;
        RECT 134.910 183.225 135.290 183.605 ;
        RECT 134.910 181.385 135.290 181.765 ;
        RECT 137.355 180.725 137.735 181.105 ;
        RECT 139.395 180.725 139.775 181.105 ;
        RECT 141.180 180.725 141.560 181.105 ;
        RECT 9.100 178.850 9.480 179.040 ;
        RECT 12.940 178.850 13.320 179.040 ;
        RECT 16.780 178.850 17.160 179.040 ;
        RECT 20.620 178.850 21.000 179.040 ;
        RECT 24.460 178.850 24.840 179.040 ;
        RECT 28.300 178.850 28.680 179.040 ;
        RECT 32.140 178.850 32.520 179.040 ;
        RECT 35.980 178.850 36.360 179.040 ;
        RECT 41.550 178.850 41.930 179.040 ;
        RECT 45.390 178.850 45.770 179.040 ;
        RECT 49.230 178.850 49.610 179.040 ;
        RECT 53.070 178.850 53.450 179.040 ;
        RECT 56.910 178.850 57.290 179.040 ;
        RECT 60.750 178.850 61.130 179.040 ;
        RECT 64.590 178.850 64.970 179.040 ;
        RECT 68.430 178.850 68.810 179.040 ;
        RECT 74.000 178.850 74.380 179.040 ;
        RECT 77.840 178.850 78.220 179.040 ;
        RECT 81.680 178.850 82.060 179.040 ;
        RECT 85.520 178.850 85.900 179.040 ;
        RECT 89.360 178.850 89.740 179.040 ;
        RECT 93.200 178.850 93.580 179.040 ;
        RECT 97.040 178.850 97.420 179.040 ;
        RECT 100.880 178.850 101.260 179.040 ;
        RECT 106.450 178.850 106.830 179.040 ;
        RECT 110.290 178.850 110.670 179.040 ;
        RECT 114.130 178.850 114.510 179.040 ;
        RECT 117.970 178.850 118.350 179.040 ;
        RECT 121.810 178.850 122.190 179.040 ;
        RECT 125.650 178.850 126.030 179.040 ;
        RECT 129.490 178.850 129.870 179.040 ;
        RECT 133.330 178.850 133.710 179.040 ;
        RECT 3.430 178.040 141.830 178.850 ;
        RECT 0.240 176.225 0.620 176.605 ;
        RECT 3.430 176.590 4.240 178.040 ;
        RECT 136.340 177.850 136.720 178.040 ;
        RECT 138.380 177.850 138.760 178.040 ;
        RECT 140.420 177.850 140.800 178.040 ;
        RECT 136.340 176.590 136.720 176.780 ;
        RECT 138.380 176.590 138.760 176.780 ;
        RECT 140.420 176.590 140.800 176.780 ;
        RECT 3.430 175.780 141.830 176.590 ;
        RECT 7.180 175.590 7.560 175.780 ;
        RECT 11.020 175.590 11.400 175.780 ;
        RECT 14.860 175.590 15.240 175.780 ;
        RECT 18.700 175.590 19.080 175.780 ;
        RECT 22.540 175.590 22.920 175.780 ;
        RECT 26.380 175.590 26.760 175.780 ;
        RECT 30.220 175.590 30.600 175.780 ;
        RECT 34.060 175.590 34.440 175.780 ;
        RECT 39.630 175.590 40.010 175.780 ;
        RECT 43.470 175.590 43.850 175.780 ;
        RECT 47.310 175.590 47.690 175.780 ;
        RECT 51.150 175.590 51.530 175.780 ;
        RECT 54.990 175.590 55.370 175.780 ;
        RECT 58.830 175.590 59.210 175.780 ;
        RECT 62.670 175.590 63.050 175.780 ;
        RECT 66.510 175.590 66.890 175.780 ;
        RECT 72.080 175.590 72.460 175.780 ;
        RECT 75.920 175.590 76.300 175.780 ;
        RECT 79.760 175.590 80.140 175.780 ;
        RECT 83.600 175.590 83.980 175.780 ;
        RECT 87.440 175.590 87.820 175.780 ;
        RECT 91.280 175.590 91.660 175.780 ;
        RECT 95.120 175.590 95.500 175.780 ;
        RECT 98.960 175.590 99.340 175.780 ;
        RECT 104.530 175.590 104.910 175.780 ;
        RECT 108.370 175.590 108.750 175.780 ;
        RECT 112.210 175.590 112.590 175.780 ;
        RECT 116.050 175.590 116.430 175.780 ;
        RECT 119.890 175.590 120.270 175.780 ;
        RECT 123.730 175.590 124.110 175.780 ;
        RECT 127.570 175.590 127.950 175.780 ;
        RECT 131.410 175.590 131.790 175.780 ;
        RECT 0.240 173.225 0.620 173.605 ;
        RECT 2.520 170.935 2.870 175.125 ;
        RECT 0.240 170.225 0.620 170.605 ;
        RECT 3.150 169.580 3.500 173.495 ;
        RECT 4.160 173.225 4.540 173.605 ;
        RECT 6.700 172.260 9.560 172.640 ;
        RECT 12.255 171.540 14.005 175.395 ;
        RECT 4.160 170.225 4.540 170.605 ;
        RECT 6.700 170.420 9.560 170.800 ;
        RECT 16.095 169.695 17.845 175.395 ;
        RECT 2.745 169.255 3.500 169.580 ;
        RECT 2.300 168.570 2.680 168.950 ;
        RECT 6.700 168.575 9.560 168.955 ;
        RECT 6.700 167.815 9.560 168.195 ;
        RECT 0.240 167.225 0.620 167.605 ;
        RECT 4.160 167.225 4.540 167.605 ;
        RECT 19.935 167.055 21.685 175.395 ;
        RECT 6.700 165.935 9.560 166.315 ;
        RECT 23.775 165.215 25.525 175.395 ;
        RECT 0.240 164.225 0.620 164.605 ;
        RECT 4.160 164.225 4.540 164.605 ;
        RECT 6.700 164.095 9.560 164.475 ;
        RECT 27.615 163.370 29.365 175.395 ;
        RECT 6.700 162.250 9.560 162.630 ;
        RECT 0.240 161.225 0.620 161.605 ;
        RECT 4.160 161.225 4.540 161.605 ;
        RECT 6.700 161.490 9.560 161.870 ;
        RECT 31.455 160.730 33.205 175.395 ;
        RECT 6.700 159.610 9.560 159.990 ;
        RECT 35.295 158.890 37.045 175.395 ;
        RECT 37.560 172.820 37.940 173.200 ;
        RECT 39.150 172.260 42.010 172.640 ;
        RECT 44.705 171.540 46.455 175.395 ;
        RECT 37.560 170.980 37.940 171.360 ;
        RECT 39.150 170.420 42.010 170.800 ;
        RECT 48.545 169.695 50.295 175.395 ;
        RECT 37.560 169.135 37.940 169.515 ;
        RECT 39.150 168.575 42.010 168.955 ;
        RECT 39.150 167.815 42.010 168.195 ;
        RECT 52.385 167.055 54.135 175.395 ;
        RECT 37.560 166.495 37.940 166.875 ;
        RECT 39.150 165.935 42.010 166.315 ;
        RECT 56.225 165.215 57.975 175.395 ;
        RECT 37.560 164.655 37.940 165.035 ;
        RECT 39.150 164.095 42.010 164.475 ;
        RECT 60.065 163.370 61.815 175.395 ;
        RECT 37.560 162.810 37.940 163.190 ;
        RECT 39.150 162.250 42.010 162.630 ;
        RECT 39.150 161.490 42.010 161.870 ;
        RECT 63.905 160.730 65.655 175.395 ;
        RECT 37.560 160.170 37.940 160.550 ;
        RECT 39.150 159.610 42.010 159.990 ;
        RECT 67.745 158.890 69.495 175.395 ;
        RECT 70.010 172.820 70.390 173.200 ;
        RECT 71.600 172.260 74.460 172.640 ;
        RECT 77.155 171.540 78.905 175.395 ;
        RECT 70.010 170.980 70.390 171.360 ;
        RECT 71.600 170.420 74.460 170.800 ;
        RECT 80.995 169.695 82.745 175.395 ;
        RECT 70.010 169.135 70.390 169.515 ;
        RECT 71.600 168.575 74.460 168.955 ;
        RECT 71.600 167.815 74.460 168.195 ;
        RECT 84.835 167.055 86.585 175.395 ;
        RECT 70.010 166.495 70.390 166.875 ;
        RECT 71.600 165.935 74.460 166.315 ;
        RECT 88.675 165.215 90.425 175.395 ;
        RECT 70.010 164.655 70.390 165.035 ;
        RECT 71.600 164.095 74.460 164.475 ;
        RECT 92.515 163.370 94.265 175.395 ;
        RECT 70.010 162.810 70.390 163.190 ;
        RECT 71.600 162.250 74.460 162.630 ;
        RECT 71.600 161.490 74.460 161.870 ;
        RECT 96.355 160.730 98.105 175.395 ;
        RECT 70.010 160.170 70.390 160.550 ;
        RECT 71.600 159.610 74.460 159.990 ;
        RECT 100.195 158.890 101.945 175.395 ;
        RECT 102.460 172.820 102.840 173.200 ;
        RECT 104.050 172.260 106.910 172.640 ;
        RECT 109.605 171.540 111.355 175.395 ;
        RECT 102.460 170.980 102.840 171.360 ;
        RECT 104.050 170.420 106.910 170.800 ;
        RECT 113.445 169.695 115.195 175.395 ;
        RECT 102.460 169.135 102.840 169.515 ;
        RECT 104.050 168.575 106.910 168.955 ;
        RECT 104.050 167.815 106.910 168.195 ;
        RECT 117.285 167.055 119.035 175.395 ;
        RECT 102.460 166.495 102.840 166.875 ;
        RECT 104.050 165.935 106.910 166.315 ;
        RECT 121.125 165.215 122.875 175.395 ;
        RECT 102.460 164.655 102.840 165.035 ;
        RECT 104.050 164.095 106.910 164.475 ;
        RECT 124.965 163.370 126.715 175.395 ;
        RECT 102.460 162.810 102.840 163.190 ;
        RECT 104.050 162.250 106.910 162.630 ;
        RECT 104.050 161.490 106.910 161.870 ;
        RECT 128.805 160.730 130.555 175.395 ;
        RECT 102.460 160.170 102.840 160.550 ;
        RECT 104.050 159.610 106.910 159.990 ;
        RECT 132.645 158.890 134.395 175.395 ;
        RECT 137.355 174.725 137.735 175.105 ;
        RECT 139.395 174.725 139.775 175.105 ;
        RECT 141.180 174.725 141.560 175.105 ;
        RECT 134.910 172.820 135.290 173.200 ;
        RECT 137.355 171.725 137.735 172.105 ;
        RECT 139.395 171.725 139.775 172.105 ;
        RECT 141.180 171.725 141.560 172.105 ;
        RECT 134.910 170.980 135.290 171.360 ;
        RECT 134.910 169.135 135.290 169.515 ;
        RECT 137.355 168.725 137.735 169.105 ;
        RECT 139.395 168.725 139.775 169.105 ;
        RECT 141.180 168.725 141.560 169.105 ;
        RECT 134.910 166.495 135.290 166.875 ;
        RECT 137.355 165.725 137.735 166.105 ;
        RECT 139.395 165.725 139.775 166.105 ;
        RECT 141.180 165.725 141.560 166.105 ;
        RECT 134.910 164.655 135.290 165.035 ;
        RECT 134.910 162.810 135.290 163.190 ;
        RECT 137.355 162.725 137.735 163.105 ;
        RECT 139.395 162.725 139.775 163.105 ;
        RECT 141.180 162.725 141.560 163.105 ;
        RECT 134.910 160.170 135.290 160.550 ;
        RECT 137.355 159.725 137.735 160.105 ;
        RECT 139.395 159.725 139.775 160.105 ;
        RECT 141.180 159.725 141.560 160.105 ;
        RECT 0.240 158.225 0.620 158.605 ;
        RECT 4.160 158.225 4.540 158.605 ;
        RECT 37.560 158.330 37.940 158.710 ;
        RECT 70.010 158.330 70.390 158.710 ;
        RECT 102.460 158.330 102.840 158.710 ;
        RECT 134.910 158.330 135.290 158.710 ;
        RECT 6.700 157.770 9.560 158.150 ;
        RECT 39.150 157.770 42.010 158.150 ;
        RECT 71.600 157.770 74.460 158.150 ;
        RECT 104.050 157.770 106.910 158.150 ;
        RECT 6.700 157.050 9.560 157.430 ;
        RECT 39.150 157.050 42.010 157.430 ;
        RECT 71.600 157.050 74.460 157.430 ;
        RECT 104.050 157.050 106.910 157.430 ;
        RECT 37.560 156.490 37.940 156.870 ;
        RECT 70.010 156.490 70.390 156.870 ;
        RECT 102.460 156.490 102.840 156.870 ;
        RECT 134.910 156.490 135.290 156.870 ;
        RECT 0.240 154.840 0.620 155.220 ;
        RECT 4.160 154.840 4.540 155.220 ;
        RECT 6.700 155.210 9.560 155.590 ;
        RECT 6.700 153.325 9.560 153.705 ;
        RECT 6.700 152.565 9.560 152.945 ;
        RECT 0.240 151.840 0.620 152.220 ;
        RECT 4.160 151.840 4.540 152.220 ;
        RECT 6.700 150.725 9.560 151.105 ;
        RECT 0.240 148.840 0.620 149.220 ;
        RECT 4.160 148.840 4.540 149.220 ;
        RECT 6.700 148.885 9.560 149.265 ;
        RECT 6.700 147.000 9.560 147.380 ;
        RECT 6.700 146.240 9.560 146.620 ;
        RECT 0.240 145.840 0.620 146.220 ;
        RECT 4.160 145.840 4.540 146.220 ;
        RECT 6.700 144.400 9.560 144.780 ;
        RECT 0.240 142.840 0.620 143.220 ;
        RECT 4.160 142.840 4.540 143.220 ;
        RECT 6.700 142.560 9.560 142.940 ;
        RECT 0.240 139.840 0.620 140.220 ;
        RECT 4.160 139.840 4.540 140.220 ;
        RECT 10.335 139.850 12.085 143.660 ;
        RECT 14.175 139.850 15.925 145.500 ;
        RECT 18.015 139.850 19.765 148.145 ;
        RECT 21.855 139.850 23.605 149.985 ;
        RECT 25.695 139.850 27.445 151.825 ;
        RECT 29.535 139.850 31.285 154.470 ;
        RECT 33.375 139.850 35.125 156.310 ;
        RECT 39.150 155.210 42.010 155.590 ;
        RECT 37.560 154.650 37.940 155.030 ;
        RECT 39.150 153.325 42.010 153.705 ;
        RECT 39.150 152.565 42.010 152.945 ;
        RECT 37.560 152.005 37.940 152.385 ;
        RECT 39.150 150.725 42.010 151.105 ;
        RECT 37.560 150.165 37.940 150.545 ;
        RECT 39.150 148.885 42.010 149.265 ;
        RECT 37.560 148.325 37.940 148.705 ;
        RECT 39.150 147.000 42.010 147.380 ;
        RECT 39.150 146.240 42.010 146.620 ;
        RECT 37.560 145.680 37.940 146.060 ;
        RECT 39.150 144.400 42.010 144.780 ;
        RECT 37.560 143.840 37.940 144.220 ;
        RECT 39.150 142.560 42.010 142.940 ;
        RECT 37.560 142.000 37.940 142.380 ;
        RECT 42.785 139.850 44.535 143.660 ;
        RECT 46.625 139.850 48.375 145.500 ;
        RECT 50.465 139.850 52.215 148.145 ;
        RECT 54.305 139.850 56.055 149.985 ;
        RECT 58.145 139.850 59.895 151.825 ;
        RECT 61.985 139.850 63.735 154.470 ;
        RECT 65.825 139.850 67.575 156.310 ;
        RECT 71.600 155.210 74.460 155.590 ;
        RECT 70.010 154.650 70.390 155.030 ;
        RECT 71.600 153.325 74.460 153.705 ;
        RECT 71.600 152.565 74.460 152.945 ;
        RECT 70.010 152.005 70.390 152.385 ;
        RECT 71.600 150.725 74.460 151.105 ;
        RECT 70.010 150.165 70.390 150.545 ;
        RECT 71.600 148.885 74.460 149.265 ;
        RECT 70.010 148.325 70.390 148.705 ;
        RECT 71.600 147.000 74.460 147.380 ;
        RECT 71.600 146.240 74.460 146.620 ;
        RECT 70.010 145.680 70.390 146.060 ;
        RECT 71.600 144.400 74.460 144.780 ;
        RECT 70.010 143.840 70.390 144.220 ;
        RECT 71.600 142.560 74.460 142.940 ;
        RECT 70.010 142.000 70.390 142.380 ;
        RECT 75.235 139.850 76.985 143.660 ;
        RECT 79.075 139.850 80.825 145.500 ;
        RECT 82.915 139.850 84.665 148.145 ;
        RECT 86.755 139.850 88.505 149.985 ;
        RECT 90.595 139.850 92.345 151.825 ;
        RECT 94.435 139.850 96.185 154.470 ;
        RECT 98.275 139.850 100.025 156.310 ;
        RECT 104.050 155.210 106.910 155.590 ;
        RECT 102.460 154.650 102.840 155.030 ;
        RECT 104.050 153.325 106.910 153.705 ;
        RECT 104.050 152.565 106.910 152.945 ;
        RECT 102.460 152.005 102.840 152.385 ;
        RECT 104.050 150.725 106.910 151.105 ;
        RECT 102.460 150.165 102.840 150.545 ;
        RECT 104.050 148.885 106.910 149.265 ;
        RECT 102.460 148.325 102.840 148.705 ;
        RECT 104.050 147.000 106.910 147.380 ;
        RECT 104.050 146.240 106.910 146.620 ;
        RECT 102.460 145.680 102.840 146.060 ;
        RECT 104.050 144.400 106.910 144.780 ;
        RECT 102.460 143.840 102.840 144.220 ;
        RECT 104.050 142.560 106.910 142.940 ;
        RECT 102.460 142.000 102.840 142.380 ;
        RECT 107.685 139.850 109.435 143.660 ;
        RECT 111.525 139.850 113.275 145.500 ;
        RECT 115.365 139.850 117.115 148.145 ;
        RECT 119.205 139.850 120.955 149.985 ;
        RECT 123.045 139.850 124.795 151.825 ;
        RECT 126.885 139.850 128.635 154.470 ;
        RECT 130.725 139.850 132.475 156.310 ;
        RECT 134.910 154.650 135.290 155.030 ;
        RECT 137.355 153.340 137.735 153.720 ;
        RECT 139.395 153.340 139.775 153.720 ;
        RECT 141.180 153.340 141.560 153.720 ;
        RECT 134.910 152.005 135.290 152.385 ;
        RECT 134.910 150.165 135.290 150.545 ;
        RECT 137.355 150.340 137.735 150.720 ;
        RECT 139.395 150.340 139.775 150.720 ;
        RECT 141.180 150.340 141.560 150.720 ;
        RECT 134.910 148.325 135.290 148.705 ;
        RECT 137.355 147.340 137.735 147.720 ;
        RECT 139.395 147.340 139.775 147.720 ;
        RECT 141.180 147.340 141.560 147.720 ;
        RECT 134.910 145.680 135.290 146.060 ;
        RECT 137.355 144.340 137.735 144.720 ;
        RECT 139.395 144.340 139.775 144.720 ;
        RECT 141.180 144.340 141.560 144.720 ;
        RECT 134.910 143.840 135.290 144.220 ;
        RECT 134.910 142.000 135.290 142.380 ;
        RECT 137.355 141.340 137.735 141.720 ;
        RECT 139.395 141.340 139.775 141.720 ;
        RECT 141.180 141.340 141.560 141.720 ;
        RECT 9.100 139.465 9.480 139.655 ;
        RECT 12.940 139.465 13.320 139.655 ;
        RECT 16.780 139.465 17.160 139.655 ;
        RECT 20.620 139.465 21.000 139.655 ;
        RECT 24.460 139.465 24.840 139.655 ;
        RECT 28.300 139.465 28.680 139.655 ;
        RECT 32.140 139.465 32.520 139.655 ;
        RECT 35.980 139.465 36.360 139.655 ;
        RECT 41.550 139.465 41.930 139.655 ;
        RECT 45.390 139.465 45.770 139.655 ;
        RECT 49.230 139.465 49.610 139.655 ;
        RECT 53.070 139.465 53.450 139.655 ;
        RECT 56.910 139.465 57.290 139.655 ;
        RECT 60.750 139.465 61.130 139.655 ;
        RECT 64.590 139.465 64.970 139.655 ;
        RECT 68.430 139.465 68.810 139.655 ;
        RECT 74.000 139.465 74.380 139.655 ;
        RECT 77.840 139.465 78.220 139.655 ;
        RECT 81.680 139.465 82.060 139.655 ;
        RECT 85.520 139.465 85.900 139.655 ;
        RECT 89.360 139.465 89.740 139.655 ;
        RECT 93.200 139.465 93.580 139.655 ;
        RECT 97.040 139.465 97.420 139.655 ;
        RECT 100.880 139.465 101.260 139.655 ;
        RECT 106.450 139.465 106.830 139.655 ;
        RECT 110.290 139.465 110.670 139.655 ;
        RECT 114.130 139.465 114.510 139.655 ;
        RECT 117.970 139.465 118.350 139.655 ;
        RECT 121.810 139.465 122.190 139.655 ;
        RECT 125.650 139.465 126.030 139.655 ;
        RECT 129.490 139.465 129.870 139.655 ;
        RECT 133.330 139.465 133.710 139.655 ;
        RECT 3.430 138.655 141.830 139.465 ;
        RECT 0.240 136.840 0.620 137.220 ;
        RECT 3.430 137.205 4.240 138.655 ;
        RECT 136.340 138.465 136.720 138.655 ;
        RECT 138.380 138.465 138.760 138.655 ;
        RECT 140.420 138.465 140.800 138.655 ;
        RECT 136.340 137.205 136.720 137.395 ;
        RECT 138.380 137.205 138.760 137.395 ;
        RECT 140.420 137.205 140.800 137.395 ;
        RECT 3.430 136.395 141.830 137.205 ;
        RECT 7.180 136.205 7.560 136.395 ;
        RECT 11.020 136.205 11.400 136.395 ;
        RECT 14.860 136.205 15.240 136.395 ;
        RECT 18.700 136.205 19.080 136.395 ;
        RECT 22.540 136.205 22.920 136.395 ;
        RECT 26.380 136.205 26.760 136.395 ;
        RECT 30.220 136.205 30.600 136.395 ;
        RECT 34.060 136.205 34.440 136.395 ;
        RECT 39.630 136.205 40.010 136.395 ;
        RECT 43.470 136.205 43.850 136.395 ;
        RECT 47.310 136.205 47.690 136.395 ;
        RECT 51.150 136.205 51.530 136.395 ;
        RECT 54.990 136.205 55.370 136.395 ;
        RECT 58.830 136.205 59.210 136.395 ;
        RECT 62.670 136.205 63.050 136.395 ;
        RECT 66.510 136.205 66.890 136.395 ;
        RECT 72.080 136.205 72.460 136.395 ;
        RECT 75.920 136.205 76.300 136.395 ;
        RECT 79.760 136.205 80.140 136.395 ;
        RECT 83.600 136.205 83.980 136.395 ;
        RECT 87.440 136.205 87.820 136.395 ;
        RECT 91.280 136.205 91.660 136.395 ;
        RECT 95.120 136.205 95.500 136.395 ;
        RECT 98.960 136.205 99.340 136.395 ;
        RECT 104.530 136.205 104.910 136.395 ;
        RECT 108.370 136.205 108.750 136.395 ;
        RECT 112.210 136.205 112.590 136.395 ;
        RECT 116.050 136.205 116.430 136.395 ;
        RECT 119.890 136.205 120.270 136.395 ;
        RECT 123.730 136.205 124.110 136.395 ;
        RECT 127.570 136.205 127.950 136.395 ;
        RECT 131.410 136.205 131.790 136.395 ;
        RECT 0.240 133.840 0.620 134.220 ;
        RECT 2.520 131.550 2.870 135.740 ;
        RECT 0.240 130.840 0.620 131.220 ;
        RECT 3.150 130.195 3.500 134.110 ;
        RECT 4.160 133.840 4.540 134.220 ;
        RECT 6.700 132.875 9.560 133.255 ;
        RECT 12.255 132.155 14.005 136.010 ;
        RECT 4.160 130.840 4.540 131.220 ;
        RECT 6.700 131.035 9.560 131.415 ;
        RECT 16.095 130.310 17.845 136.010 ;
        RECT 2.745 129.870 3.500 130.195 ;
        RECT 2.300 129.185 2.680 129.565 ;
        RECT 6.700 129.190 9.560 129.570 ;
        RECT 6.700 128.430 9.560 128.810 ;
        RECT 0.240 127.840 0.620 128.220 ;
        RECT 4.160 127.840 4.540 128.220 ;
        RECT 19.935 127.670 21.685 136.010 ;
        RECT 6.700 126.550 9.560 126.930 ;
        RECT 23.775 125.830 25.525 136.010 ;
        RECT 0.240 124.840 0.620 125.220 ;
        RECT 4.160 124.840 4.540 125.220 ;
        RECT 6.700 124.710 9.560 125.090 ;
        RECT 27.615 123.985 29.365 136.010 ;
        RECT 6.700 122.865 9.560 123.245 ;
        RECT 0.240 121.840 0.620 122.220 ;
        RECT 4.160 121.840 4.540 122.220 ;
        RECT 6.700 122.105 9.560 122.485 ;
        RECT 31.455 121.345 33.205 136.010 ;
        RECT 6.700 120.225 9.560 120.605 ;
        RECT 35.295 119.505 37.045 136.010 ;
        RECT 37.560 133.435 37.940 133.815 ;
        RECT 39.150 132.875 42.010 133.255 ;
        RECT 44.705 132.155 46.455 136.010 ;
        RECT 37.560 131.595 37.940 131.975 ;
        RECT 39.150 131.035 42.010 131.415 ;
        RECT 48.545 130.310 50.295 136.010 ;
        RECT 37.560 129.750 37.940 130.130 ;
        RECT 39.150 129.190 42.010 129.570 ;
        RECT 39.150 128.430 42.010 128.810 ;
        RECT 52.385 127.670 54.135 136.010 ;
        RECT 37.560 127.110 37.940 127.490 ;
        RECT 39.150 126.550 42.010 126.930 ;
        RECT 56.225 125.830 57.975 136.010 ;
        RECT 37.560 125.270 37.940 125.650 ;
        RECT 39.150 124.710 42.010 125.090 ;
        RECT 60.065 123.985 61.815 136.010 ;
        RECT 37.560 123.425 37.940 123.805 ;
        RECT 39.150 122.865 42.010 123.245 ;
        RECT 39.150 122.105 42.010 122.485 ;
        RECT 63.905 121.345 65.655 136.010 ;
        RECT 37.560 120.785 37.940 121.165 ;
        RECT 39.150 120.225 42.010 120.605 ;
        RECT 67.745 119.505 69.495 136.010 ;
        RECT 70.010 133.435 70.390 133.815 ;
        RECT 71.600 132.875 74.460 133.255 ;
        RECT 77.155 132.155 78.905 136.010 ;
        RECT 70.010 131.595 70.390 131.975 ;
        RECT 71.600 131.035 74.460 131.415 ;
        RECT 80.995 130.310 82.745 136.010 ;
        RECT 70.010 129.750 70.390 130.130 ;
        RECT 71.600 129.190 74.460 129.570 ;
        RECT 71.600 128.430 74.460 128.810 ;
        RECT 84.835 127.670 86.585 136.010 ;
        RECT 70.010 127.110 70.390 127.490 ;
        RECT 71.600 126.550 74.460 126.930 ;
        RECT 88.675 125.830 90.425 136.010 ;
        RECT 70.010 125.270 70.390 125.650 ;
        RECT 71.600 124.710 74.460 125.090 ;
        RECT 92.515 123.985 94.265 136.010 ;
        RECT 70.010 123.425 70.390 123.805 ;
        RECT 71.600 122.865 74.460 123.245 ;
        RECT 71.600 122.105 74.460 122.485 ;
        RECT 96.355 121.345 98.105 136.010 ;
        RECT 70.010 120.785 70.390 121.165 ;
        RECT 71.600 120.225 74.460 120.605 ;
        RECT 100.195 119.505 101.945 136.010 ;
        RECT 102.460 133.435 102.840 133.815 ;
        RECT 104.050 132.875 106.910 133.255 ;
        RECT 109.605 132.155 111.355 136.010 ;
        RECT 102.460 131.595 102.840 131.975 ;
        RECT 104.050 131.035 106.910 131.415 ;
        RECT 113.445 130.310 115.195 136.010 ;
        RECT 102.460 129.750 102.840 130.130 ;
        RECT 104.050 129.190 106.910 129.570 ;
        RECT 104.050 128.430 106.910 128.810 ;
        RECT 117.285 127.670 119.035 136.010 ;
        RECT 102.460 127.110 102.840 127.490 ;
        RECT 104.050 126.550 106.910 126.930 ;
        RECT 121.125 125.830 122.875 136.010 ;
        RECT 102.460 125.270 102.840 125.650 ;
        RECT 104.050 124.710 106.910 125.090 ;
        RECT 124.965 123.985 126.715 136.010 ;
        RECT 102.460 123.425 102.840 123.805 ;
        RECT 104.050 122.865 106.910 123.245 ;
        RECT 104.050 122.105 106.910 122.485 ;
        RECT 128.805 121.345 130.555 136.010 ;
        RECT 102.460 120.785 102.840 121.165 ;
        RECT 104.050 120.225 106.910 120.605 ;
        RECT 132.645 119.505 134.395 136.010 ;
        RECT 137.355 135.340 137.735 135.720 ;
        RECT 139.395 135.340 139.775 135.720 ;
        RECT 141.180 135.340 141.560 135.720 ;
        RECT 134.910 133.435 135.290 133.815 ;
        RECT 137.355 132.340 137.735 132.720 ;
        RECT 139.395 132.340 139.775 132.720 ;
        RECT 141.180 132.340 141.560 132.720 ;
        RECT 134.910 131.595 135.290 131.975 ;
        RECT 134.910 129.750 135.290 130.130 ;
        RECT 137.355 129.340 137.735 129.720 ;
        RECT 139.395 129.340 139.775 129.720 ;
        RECT 141.180 129.340 141.560 129.720 ;
        RECT 134.910 127.110 135.290 127.490 ;
        RECT 137.355 126.340 137.735 126.720 ;
        RECT 139.395 126.340 139.775 126.720 ;
        RECT 141.180 126.340 141.560 126.720 ;
        RECT 134.910 125.270 135.290 125.650 ;
        RECT 134.910 123.425 135.290 123.805 ;
        RECT 137.355 123.340 137.735 123.720 ;
        RECT 139.395 123.340 139.775 123.720 ;
        RECT 141.180 123.340 141.560 123.720 ;
        RECT 134.910 120.785 135.290 121.165 ;
        RECT 137.355 120.340 137.735 120.720 ;
        RECT 139.395 120.340 139.775 120.720 ;
        RECT 141.180 120.340 141.560 120.720 ;
        RECT 0.240 118.840 0.620 119.220 ;
        RECT 4.160 118.840 4.540 119.220 ;
        RECT 37.560 118.945 37.940 119.325 ;
        RECT 70.010 118.945 70.390 119.325 ;
        RECT 102.460 118.945 102.840 119.325 ;
        RECT 134.910 118.945 135.290 119.325 ;
        RECT 6.700 118.385 9.560 118.765 ;
        RECT 39.150 118.385 42.010 118.765 ;
        RECT 71.600 118.385 74.460 118.765 ;
        RECT 104.050 118.385 106.910 118.765 ;
        RECT 6.700 117.665 9.560 118.045 ;
        RECT 39.150 117.665 42.010 118.045 ;
        RECT 71.600 117.665 74.460 118.045 ;
        RECT 104.050 117.665 106.910 118.045 ;
        RECT 37.560 117.105 37.940 117.485 ;
        RECT 70.010 117.105 70.390 117.485 ;
        RECT 102.460 117.105 102.840 117.485 ;
        RECT 134.910 117.105 135.290 117.485 ;
        RECT 0.240 115.455 0.620 115.835 ;
        RECT 4.160 115.455 4.540 115.835 ;
        RECT 6.700 115.825 9.560 116.205 ;
        RECT 6.700 113.940 9.560 114.320 ;
        RECT 6.700 113.180 9.560 113.560 ;
        RECT 0.240 112.455 0.620 112.835 ;
        RECT 4.160 112.455 4.540 112.835 ;
        RECT 6.700 111.340 9.560 111.720 ;
        RECT 0.240 109.455 0.620 109.835 ;
        RECT 4.160 109.455 4.540 109.835 ;
        RECT 6.700 109.500 9.560 109.880 ;
        RECT 6.700 107.615 9.560 107.995 ;
        RECT 6.700 106.855 9.560 107.235 ;
        RECT 0.240 106.455 0.620 106.835 ;
        RECT 4.160 106.455 4.540 106.835 ;
        RECT 6.700 105.015 9.560 105.395 ;
        RECT 0.240 103.455 0.620 103.835 ;
        RECT 4.160 103.455 4.540 103.835 ;
        RECT 6.700 103.175 9.560 103.555 ;
        RECT 0.240 100.455 0.620 100.835 ;
        RECT 4.160 100.455 4.540 100.835 ;
        RECT 10.335 100.465 12.085 104.275 ;
        RECT 14.175 100.465 15.925 106.115 ;
        RECT 18.015 100.465 19.765 108.760 ;
        RECT 21.855 100.465 23.605 110.600 ;
        RECT 25.695 100.465 27.445 112.440 ;
        RECT 29.535 100.465 31.285 115.085 ;
        RECT 33.375 100.465 35.125 116.925 ;
        RECT 39.150 115.825 42.010 116.205 ;
        RECT 37.560 115.265 37.940 115.645 ;
        RECT 39.150 113.940 42.010 114.320 ;
        RECT 39.150 113.180 42.010 113.560 ;
        RECT 37.560 112.620 37.940 113.000 ;
        RECT 39.150 111.340 42.010 111.720 ;
        RECT 37.560 110.780 37.940 111.160 ;
        RECT 39.150 109.500 42.010 109.880 ;
        RECT 37.560 108.940 37.940 109.320 ;
        RECT 39.150 107.615 42.010 107.995 ;
        RECT 39.150 106.855 42.010 107.235 ;
        RECT 37.560 106.295 37.940 106.675 ;
        RECT 39.150 105.015 42.010 105.395 ;
        RECT 37.560 104.455 37.940 104.835 ;
        RECT 39.150 103.175 42.010 103.555 ;
        RECT 37.560 102.615 37.940 102.995 ;
        RECT 42.785 100.465 44.535 104.275 ;
        RECT 46.625 100.465 48.375 106.115 ;
        RECT 50.465 100.465 52.215 108.760 ;
        RECT 54.305 100.465 56.055 110.600 ;
        RECT 58.145 100.465 59.895 112.440 ;
        RECT 61.985 100.465 63.735 115.085 ;
        RECT 65.825 100.465 67.575 116.925 ;
        RECT 71.600 115.825 74.460 116.205 ;
        RECT 70.010 115.265 70.390 115.645 ;
        RECT 71.600 113.940 74.460 114.320 ;
        RECT 71.600 113.180 74.460 113.560 ;
        RECT 70.010 112.620 70.390 113.000 ;
        RECT 71.600 111.340 74.460 111.720 ;
        RECT 70.010 110.780 70.390 111.160 ;
        RECT 71.600 109.500 74.460 109.880 ;
        RECT 70.010 108.940 70.390 109.320 ;
        RECT 71.600 107.615 74.460 107.995 ;
        RECT 71.600 106.855 74.460 107.235 ;
        RECT 70.010 106.295 70.390 106.675 ;
        RECT 71.600 105.015 74.460 105.395 ;
        RECT 70.010 104.455 70.390 104.835 ;
        RECT 71.600 103.175 74.460 103.555 ;
        RECT 70.010 102.615 70.390 102.995 ;
        RECT 75.235 100.465 76.985 104.275 ;
        RECT 79.075 100.465 80.825 106.115 ;
        RECT 82.915 100.465 84.665 108.760 ;
        RECT 86.755 100.465 88.505 110.600 ;
        RECT 90.595 100.465 92.345 112.440 ;
        RECT 94.435 100.465 96.185 115.085 ;
        RECT 98.275 100.465 100.025 116.925 ;
        RECT 104.050 115.825 106.910 116.205 ;
        RECT 102.460 115.265 102.840 115.645 ;
        RECT 104.050 113.940 106.910 114.320 ;
        RECT 104.050 113.180 106.910 113.560 ;
        RECT 102.460 112.620 102.840 113.000 ;
        RECT 104.050 111.340 106.910 111.720 ;
        RECT 102.460 110.780 102.840 111.160 ;
        RECT 104.050 109.500 106.910 109.880 ;
        RECT 102.460 108.940 102.840 109.320 ;
        RECT 104.050 107.615 106.910 107.995 ;
        RECT 104.050 106.855 106.910 107.235 ;
        RECT 102.460 106.295 102.840 106.675 ;
        RECT 104.050 105.015 106.910 105.395 ;
        RECT 102.460 104.455 102.840 104.835 ;
        RECT 104.050 103.175 106.910 103.555 ;
        RECT 102.460 102.615 102.840 102.995 ;
        RECT 107.685 100.465 109.435 104.275 ;
        RECT 111.525 100.465 113.275 106.115 ;
        RECT 115.365 100.465 117.115 108.760 ;
        RECT 119.205 100.465 120.955 110.600 ;
        RECT 123.045 100.465 124.795 112.440 ;
        RECT 126.885 100.465 128.635 115.085 ;
        RECT 130.725 100.465 132.475 116.925 ;
        RECT 134.910 115.265 135.290 115.645 ;
        RECT 137.355 113.955 137.735 114.335 ;
        RECT 139.395 113.955 139.775 114.335 ;
        RECT 141.180 113.955 141.560 114.335 ;
        RECT 134.910 112.620 135.290 113.000 ;
        RECT 134.910 110.780 135.290 111.160 ;
        RECT 137.355 110.955 137.735 111.335 ;
        RECT 139.395 110.955 139.775 111.335 ;
        RECT 141.180 110.955 141.560 111.335 ;
        RECT 134.910 108.940 135.290 109.320 ;
        RECT 137.355 107.955 137.735 108.335 ;
        RECT 139.395 107.955 139.775 108.335 ;
        RECT 141.180 107.955 141.560 108.335 ;
        RECT 134.910 106.295 135.290 106.675 ;
        RECT 137.355 104.955 137.735 105.335 ;
        RECT 139.395 104.955 139.775 105.335 ;
        RECT 141.180 104.955 141.560 105.335 ;
        RECT 134.910 104.455 135.290 104.835 ;
        RECT 134.910 102.615 135.290 102.995 ;
        RECT 137.355 101.955 137.735 102.335 ;
        RECT 139.395 101.955 139.775 102.335 ;
        RECT 141.180 101.955 141.560 102.335 ;
        RECT 9.100 100.080 9.480 100.270 ;
        RECT 12.940 100.080 13.320 100.270 ;
        RECT 16.780 100.080 17.160 100.270 ;
        RECT 20.620 100.080 21.000 100.270 ;
        RECT 24.460 100.080 24.840 100.270 ;
        RECT 28.300 100.080 28.680 100.270 ;
        RECT 32.140 100.080 32.520 100.270 ;
        RECT 35.980 100.080 36.360 100.270 ;
        RECT 41.550 100.080 41.930 100.270 ;
        RECT 45.390 100.080 45.770 100.270 ;
        RECT 49.230 100.080 49.610 100.270 ;
        RECT 53.070 100.080 53.450 100.270 ;
        RECT 56.910 100.080 57.290 100.270 ;
        RECT 60.750 100.080 61.130 100.270 ;
        RECT 64.590 100.080 64.970 100.270 ;
        RECT 68.430 100.080 68.810 100.270 ;
        RECT 74.000 100.080 74.380 100.270 ;
        RECT 77.840 100.080 78.220 100.270 ;
        RECT 81.680 100.080 82.060 100.270 ;
        RECT 85.520 100.080 85.900 100.270 ;
        RECT 89.360 100.080 89.740 100.270 ;
        RECT 93.200 100.080 93.580 100.270 ;
        RECT 97.040 100.080 97.420 100.270 ;
        RECT 100.880 100.080 101.260 100.270 ;
        RECT 106.450 100.080 106.830 100.270 ;
        RECT 110.290 100.080 110.670 100.270 ;
        RECT 114.130 100.080 114.510 100.270 ;
        RECT 117.970 100.080 118.350 100.270 ;
        RECT 121.810 100.080 122.190 100.270 ;
        RECT 125.650 100.080 126.030 100.270 ;
        RECT 129.490 100.080 129.870 100.270 ;
        RECT 133.330 100.080 133.710 100.270 ;
        RECT 3.430 99.270 141.830 100.080 ;
        RECT 0.240 97.455 0.620 97.835 ;
        RECT 3.430 97.820 4.240 99.270 ;
        RECT 136.340 99.080 136.720 99.270 ;
        RECT 138.380 99.080 138.760 99.270 ;
        RECT 140.420 99.080 140.800 99.270 ;
        RECT 136.340 97.820 136.720 98.010 ;
        RECT 138.380 97.820 138.760 98.010 ;
        RECT 140.420 97.820 140.800 98.010 ;
        RECT 3.430 97.010 141.830 97.820 ;
        RECT 7.180 96.820 7.560 97.010 ;
        RECT 11.020 96.820 11.400 97.010 ;
        RECT 14.860 96.820 15.240 97.010 ;
        RECT 18.700 96.820 19.080 97.010 ;
        RECT 22.540 96.820 22.920 97.010 ;
        RECT 26.380 96.820 26.760 97.010 ;
        RECT 30.220 96.820 30.600 97.010 ;
        RECT 34.060 96.820 34.440 97.010 ;
        RECT 39.630 96.820 40.010 97.010 ;
        RECT 43.470 96.820 43.850 97.010 ;
        RECT 47.310 96.820 47.690 97.010 ;
        RECT 51.150 96.820 51.530 97.010 ;
        RECT 54.990 96.820 55.370 97.010 ;
        RECT 58.830 96.820 59.210 97.010 ;
        RECT 62.670 96.820 63.050 97.010 ;
        RECT 66.510 96.820 66.890 97.010 ;
        RECT 72.080 96.820 72.460 97.010 ;
        RECT 75.920 96.820 76.300 97.010 ;
        RECT 79.760 96.820 80.140 97.010 ;
        RECT 83.600 96.820 83.980 97.010 ;
        RECT 87.440 96.820 87.820 97.010 ;
        RECT 91.280 96.820 91.660 97.010 ;
        RECT 95.120 96.820 95.500 97.010 ;
        RECT 98.960 96.820 99.340 97.010 ;
        RECT 104.530 96.820 104.910 97.010 ;
        RECT 108.370 96.820 108.750 97.010 ;
        RECT 112.210 96.820 112.590 97.010 ;
        RECT 116.050 96.820 116.430 97.010 ;
        RECT 119.890 96.820 120.270 97.010 ;
        RECT 123.730 96.820 124.110 97.010 ;
        RECT 127.570 96.820 127.950 97.010 ;
        RECT 131.410 96.820 131.790 97.010 ;
        RECT 0.240 94.455 0.620 94.835 ;
        RECT 2.520 92.165 2.870 96.355 ;
        RECT 0.240 91.455 0.620 91.835 ;
        RECT 3.150 90.810 3.500 94.725 ;
        RECT 4.160 94.455 4.540 94.835 ;
        RECT 6.700 93.490 9.560 93.870 ;
        RECT 12.255 92.770 14.005 96.625 ;
        RECT 4.160 91.455 4.540 91.835 ;
        RECT 6.700 91.650 9.560 92.030 ;
        RECT 16.095 90.925 17.845 96.625 ;
        RECT 2.745 90.485 3.500 90.810 ;
        RECT 2.300 89.800 2.680 90.180 ;
        RECT 6.700 89.805 9.560 90.185 ;
        RECT 6.700 89.045 9.560 89.425 ;
        RECT 0.240 88.455 0.620 88.835 ;
        RECT 4.160 88.455 4.540 88.835 ;
        RECT 19.935 88.285 21.685 96.625 ;
        RECT 6.700 87.165 9.560 87.545 ;
        RECT 23.775 86.445 25.525 96.625 ;
        RECT 0.240 85.455 0.620 85.835 ;
        RECT 4.160 85.455 4.540 85.835 ;
        RECT 6.700 85.325 9.560 85.705 ;
        RECT 27.615 84.600 29.365 96.625 ;
        RECT 6.700 83.480 9.560 83.860 ;
        RECT 0.240 82.455 0.620 82.835 ;
        RECT 4.160 82.455 4.540 82.835 ;
        RECT 6.700 82.720 9.560 83.100 ;
        RECT 31.455 81.960 33.205 96.625 ;
        RECT 6.700 80.840 9.560 81.220 ;
        RECT 35.295 80.120 37.045 96.625 ;
        RECT 37.560 94.050 37.940 94.430 ;
        RECT 39.150 93.490 42.010 93.870 ;
        RECT 44.705 92.770 46.455 96.625 ;
        RECT 37.560 92.210 37.940 92.590 ;
        RECT 39.150 91.650 42.010 92.030 ;
        RECT 48.545 90.925 50.295 96.625 ;
        RECT 37.560 90.365 37.940 90.745 ;
        RECT 39.150 89.805 42.010 90.185 ;
        RECT 39.150 89.045 42.010 89.425 ;
        RECT 52.385 88.285 54.135 96.625 ;
        RECT 37.560 87.725 37.940 88.105 ;
        RECT 39.150 87.165 42.010 87.545 ;
        RECT 56.225 86.445 57.975 96.625 ;
        RECT 37.560 85.885 37.940 86.265 ;
        RECT 39.150 85.325 42.010 85.705 ;
        RECT 60.065 84.600 61.815 96.625 ;
        RECT 37.560 84.040 37.940 84.420 ;
        RECT 39.150 83.480 42.010 83.860 ;
        RECT 39.150 82.720 42.010 83.100 ;
        RECT 63.905 81.960 65.655 96.625 ;
        RECT 37.560 81.400 37.940 81.780 ;
        RECT 39.150 80.840 42.010 81.220 ;
        RECT 67.745 80.120 69.495 96.625 ;
        RECT 70.010 94.050 70.390 94.430 ;
        RECT 71.600 93.490 74.460 93.870 ;
        RECT 77.155 92.770 78.905 96.625 ;
        RECT 70.010 92.210 70.390 92.590 ;
        RECT 71.600 91.650 74.460 92.030 ;
        RECT 80.995 90.925 82.745 96.625 ;
        RECT 70.010 90.365 70.390 90.745 ;
        RECT 71.600 89.805 74.460 90.185 ;
        RECT 71.600 89.045 74.460 89.425 ;
        RECT 84.835 88.285 86.585 96.625 ;
        RECT 70.010 87.725 70.390 88.105 ;
        RECT 71.600 87.165 74.460 87.545 ;
        RECT 88.675 86.445 90.425 96.625 ;
        RECT 70.010 85.885 70.390 86.265 ;
        RECT 71.600 85.325 74.460 85.705 ;
        RECT 92.515 84.600 94.265 96.625 ;
        RECT 70.010 84.040 70.390 84.420 ;
        RECT 71.600 83.480 74.460 83.860 ;
        RECT 71.600 82.720 74.460 83.100 ;
        RECT 96.355 81.960 98.105 96.625 ;
        RECT 70.010 81.400 70.390 81.780 ;
        RECT 71.600 80.840 74.460 81.220 ;
        RECT 100.195 80.120 101.945 96.625 ;
        RECT 102.460 94.050 102.840 94.430 ;
        RECT 104.050 93.490 106.910 93.870 ;
        RECT 109.605 92.770 111.355 96.625 ;
        RECT 102.460 92.210 102.840 92.590 ;
        RECT 104.050 91.650 106.910 92.030 ;
        RECT 113.445 90.925 115.195 96.625 ;
        RECT 102.460 90.365 102.840 90.745 ;
        RECT 104.050 89.805 106.910 90.185 ;
        RECT 104.050 89.045 106.910 89.425 ;
        RECT 117.285 88.285 119.035 96.625 ;
        RECT 102.460 87.725 102.840 88.105 ;
        RECT 104.050 87.165 106.910 87.545 ;
        RECT 121.125 86.445 122.875 96.625 ;
        RECT 102.460 85.885 102.840 86.265 ;
        RECT 104.050 85.325 106.910 85.705 ;
        RECT 124.965 84.600 126.715 96.625 ;
        RECT 102.460 84.040 102.840 84.420 ;
        RECT 104.050 83.480 106.910 83.860 ;
        RECT 104.050 82.720 106.910 83.100 ;
        RECT 128.805 81.960 130.555 96.625 ;
        RECT 102.460 81.400 102.840 81.780 ;
        RECT 104.050 80.840 106.910 81.220 ;
        RECT 132.645 80.120 134.395 96.625 ;
        RECT 137.355 95.955 137.735 96.335 ;
        RECT 139.395 95.955 139.775 96.335 ;
        RECT 141.180 95.955 141.560 96.335 ;
        RECT 134.910 94.050 135.290 94.430 ;
        RECT 137.355 92.955 137.735 93.335 ;
        RECT 139.395 92.955 139.775 93.335 ;
        RECT 141.180 92.955 141.560 93.335 ;
        RECT 134.910 92.210 135.290 92.590 ;
        RECT 134.910 90.365 135.290 90.745 ;
        RECT 137.355 89.955 137.735 90.335 ;
        RECT 139.395 89.955 139.775 90.335 ;
        RECT 141.180 89.955 141.560 90.335 ;
        RECT 134.910 87.725 135.290 88.105 ;
        RECT 137.355 86.955 137.735 87.335 ;
        RECT 139.395 86.955 139.775 87.335 ;
        RECT 141.180 86.955 141.560 87.335 ;
        RECT 134.910 85.885 135.290 86.265 ;
        RECT 134.910 84.040 135.290 84.420 ;
        RECT 137.355 83.955 137.735 84.335 ;
        RECT 139.395 83.955 139.775 84.335 ;
        RECT 141.180 83.955 141.560 84.335 ;
        RECT 134.910 81.400 135.290 81.780 ;
        RECT 137.355 80.955 137.735 81.335 ;
        RECT 139.395 80.955 139.775 81.335 ;
        RECT 141.180 80.955 141.560 81.335 ;
        RECT 0.240 79.455 0.620 79.835 ;
        RECT 4.160 79.455 4.540 79.835 ;
        RECT 37.560 79.560 37.940 79.940 ;
        RECT 70.010 79.560 70.390 79.940 ;
        RECT 102.460 79.560 102.840 79.940 ;
        RECT 134.910 79.560 135.290 79.940 ;
        RECT 6.700 79.000 9.560 79.380 ;
        RECT 39.150 79.000 42.010 79.380 ;
        RECT 71.600 79.000 74.460 79.380 ;
        RECT 104.050 79.000 106.910 79.380 ;
        RECT 6.700 78.280 9.560 78.660 ;
        RECT 39.150 78.280 42.010 78.660 ;
        RECT 71.600 78.280 74.460 78.660 ;
        RECT 104.050 78.280 106.910 78.660 ;
        RECT 37.560 77.720 37.940 78.100 ;
        RECT 70.010 77.720 70.390 78.100 ;
        RECT 102.460 77.720 102.840 78.100 ;
        RECT 134.910 77.720 135.290 78.100 ;
        RECT 0.240 76.070 0.620 76.450 ;
        RECT 4.160 76.070 4.540 76.450 ;
        RECT 6.700 76.440 9.560 76.820 ;
        RECT 6.700 74.555 9.560 74.935 ;
        RECT 6.700 73.795 9.560 74.175 ;
        RECT 0.240 73.070 0.620 73.450 ;
        RECT 4.160 73.070 4.540 73.450 ;
        RECT 6.700 71.955 9.560 72.335 ;
        RECT 0.240 70.070 0.620 70.450 ;
        RECT 4.160 70.070 4.540 70.450 ;
        RECT 6.700 70.115 9.560 70.495 ;
        RECT 6.700 68.230 9.560 68.610 ;
        RECT 6.700 67.470 9.560 67.850 ;
        RECT 0.240 67.070 0.620 67.450 ;
        RECT 4.160 67.070 4.540 67.450 ;
        RECT 6.700 65.630 9.560 66.010 ;
        RECT 0.240 64.070 0.620 64.450 ;
        RECT 4.160 64.070 4.540 64.450 ;
        RECT 6.700 63.790 9.560 64.170 ;
        RECT 0.240 61.070 0.620 61.450 ;
        RECT 4.160 61.070 4.540 61.450 ;
        RECT 10.335 61.080 12.085 64.890 ;
        RECT 14.175 61.080 15.925 66.730 ;
        RECT 18.015 61.080 19.765 69.375 ;
        RECT 21.855 61.080 23.605 71.215 ;
        RECT 25.695 61.080 27.445 73.055 ;
        RECT 29.535 61.080 31.285 75.700 ;
        RECT 33.375 61.080 35.125 77.540 ;
        RECT 39.150 76.440 42.010 76.820 ;
        RECT 37.560 75.880 37.940 76.260 ;
        RECT 39.150 74.555 42.010 74.935 ;
        RECT 39.150 73.795 42.010 74.175 ;
        RECT 37.560 73.235 37.940 73.615 ;
        RECT 39.150 71.955 42.010 72.335 ;
        RECT 37.560 71.395 37.940 71.775 ;
        RECT 39.150 70.115 42.010 70.495 ;
        RECT 37.560 69.555 37.940 69.935 ;
        RECT 39.150 68.230 42.010 68.610 ;
        RECT 39.150 67.470 42.010 67.850 ;
        RECT 37.560 66.910 37.940 67.290 ;
        RECT 39.150 65.630 42.010 66.010 ;
        RECT 37.560 65.070 37.940 65.450 ;
        RECT 39.150 63.790 42.010 64.170 ;
        RECT 37.560 63.230 37.940 63.610 ;
        RECT 42.785 61.080 44.535 64.890 ;
        RECT 46.625 61.080 48.375 66.730 ;
        RECT 50.465 61.080 52.215 69.375 ;
        RECT 54.305 61.080 56.055 71.215 ;
        RECT 58.145 61.080 59.895 73.055 ;
        RECT 61.985 61.080 63.735 75.700 ;
        RECT 65.825 61.080 67.575 77.540 ;
        RECT 71.600 76.440 74.460 76.820 ;
        RECT 70.010 75.880 70.390 76.260 ;
        RECT 71.600 74.555 74.460 74.935 ;
        RECT 71.600 73.795 74.460 74.175 ;
        RECT 70.010 73.235 70.390 73.615 ;
        RECT 71.600 71.955 74.460 72.335 ;
        RECT 70.010 71.395 70.390 71.775 ;
        RECT 71.600 70.115 74.460 70.495 ;
        RECT 70.010 69.555 70.390 69.935 ;
        RECT 71.600 68.230 74.460 68.610 ;
        RECT 71.600 67.470 74.460 67.850 ;
        RECT 70.010 66.910 70.390 67.290 ;
        RECT 71.600 65.630 74.460 66.010 ;
        RECT 70.010 65.070 70.390 65.450 ;
        RECT 71.600 63.790 74.460 64.170 ;
        RECT 70.010 63.230 70.390 63.610 ;
        RECT 75.235 61.080 76.985 64.890 ;
        RECT 79.075 61.080 80.825 66.730 ;
        RECT 82.915 61.080 84.665 69.375 ;
        RECT 86.755 61.080 88.505 71.215 ;
        RECT 90.595 61.080 92.345 73.055 ;
        RECT 94.435 61.080 96.185 75.700 ;
        RECT 98.275 61.080 100.025 77.540 ;
        RECT 104.050 76.440 106.910 76.820 ;
        RECT 102.460 75.880 102.840 76.260 ;
        RECT 104.050 74.555 106.910 74.935 ;
        RECT 104.050 73.795 106.910 74.175 ;
        RECT 102.460 73.235 102.840 73.615 ;
        RECT 104.050 71.955 106.910 72.335 ;
        RECT 102.460 71.395 102.840 71.775 ;
        RECT 104.050 70.115 106.910 70.495 ;
        RECT 102.460 69.555 102.840 69.935 ;
        RECT 104.050 68.230 106.910 68.610 ;
        RECT 104.050 67.470 106.910 67.850 ;
        RECT 102.460 66.910 102.840 67.290 ;
        RECT 104.050 65.630 106.910 66.010 ;
        RECT 102.460 65.070 102.840 65.450 ;
        RECT 104.050 63.790 106.910 64.170 ;
        RECT 102.460 63.230 102.840 63.610 ;
        RECT 107.685 61.080 109.435 64.890 ;
        RECT 111.525 61.080 113.275 66.730 ;
        RECT 115.365 61.080 117.115 69.375 ;
        RECT 119.205 61.080 120.955 71.215 ;
        RECT 123.045 61.080 124.795 73.055 ;
        RECT 126.885 61.080 128.635 75.700 ;
        RECT 130.725 61.080 132.475 77.540 ;
        RECT 134.910 75.880 135.290 76.260 ;
        RECT 137.355 74.570 137.735 74.950 ;
        RECT 139.395 74.570 139.775 74.950 ;
        RECT 141.180 74.570 141.560 74.950 ;
        RECT 134.910 73.235 135.290 73.615 ;
        RECT 134.910 71.395 135.290 71.775 ;
        RECT 137.355 71.570 137.735 71.950 ;
        RECT 139.395 71.570 139.775 71.950 ;
        RECT 141.180 71.570 141.560 71.950 ;
        RECT 134.910 69.555 135.290 69.935 ;
        RECT 137.355 68.570 137.735 68.950 ;
        RECT 139.395 68.570 139.775 68.950 ;
        RECT 141.180 68.570 141.560 68.950 ;
        RECT 134.910 66.910 135.290 67.290 ;
        RECT 137.355 65.570 137.735 65.950 ;
        RECT 139.395 65.570 139.775 65.950 ;
        RECT 141.180 65.570 141.560 65.950 ;
        RECT 134.910 65.070 135.290 65.450 ;
        RECT 134.910 63.230 135.290 63.610 ;
        RECT 137.355 62.570 137.735 62.950 ;
        RECT 139.395 62.570 139.775 62.950 ;
        RECT 141.180 62.570 141.560 62.950 ;
        RECT 9.100 60.695 9.480 60.885 ;
        RECT 12.940 60.695 13.320 60.885 ;
        RECT 16.780 60.695 17.160 60.885 ;
        RECT 20.620 60.695 21.000 60.885 ;
        RECT 24.460 60.695 24.840 60.885 ;
        RECT 28.300 60.695 28.680 60.885 ;
        RECT 32.140 60.695 32.520 60.885 ;
        RECT 35.980 60.695 36.360 60.885 ;
        RECT 41.550 60.695 41.930 60.885 ;
        RECT 45.390 60.695 45.770 60.885 ;
        RECT 49.230 60.695 49.610 60.885 ;
        RECT 53.070 60.695 53.450 60.885 ;
        RECT 56.910 60.695 57.290 60.885 ;
        RECT 60.750 60.695 61.130 60.885 ;
        RECT 64.590 60.695 64.970 60.885 ;
        RECT 68.430 60.695 68.810 60.885 ;
        RECT 74.000 60.695 74.380 60.885 ;
        RECT 77.840 60.695 78.220 60.885 ;
        RECT 81.680 60.695 82.060 60.885 ;
        RECT 85.520 60.695 85.900 60.885 ;
        RECT 89.360 60.695 89.740 60.885 ;
        RECT 93.200 60.695 93.580 60.885 ;
        RECT 97.040 60.695 97.420 60.885 ;
        RECT 100.880 60.695 101.260 60.885 ;
        RECT 106.450 60.695 106.830 60.885 ;
        RECT 110.290 60.695 110.670 60.885 ;
        RECT 114.130 60.695 114.510 60.885 ;
        RECT 117.970 60.695 118.350 60.885 ;
        RECT 121.810 60.695 122.190 60.885 ;
        RECT 125.650 60.695 126.030 60.885 ;
        RECT 129.490 60.695 129.870 60.885 ;
        RECT 133.330 60.695 133.710 60.885 ;
        RECT 3.430 59.885 141.830 60.695 ;
        RECT 0.240 58.070 0.620 58.450 ;
        RECT 3.430 58.435 4.240 59.885 ;
        RECT 136.340 59.695 136.720 59.885 ;
        RECT 138.380 59.695 138.760 59.885 ;
        RECT 140.420 59.695 140.800 59.885 ;
        RECT 136.340 58.435 136.720 58.625 ;
        RECT 138.380 58.435 138.760 58.625 ;
        RECT 140.420 58.435 140.800 58.625 ;
        RECT 3.430 57.625 141.830 58.435 ;
        RECT 7.180 57.435 7.560 57.625 ;
        RECT 11.020 57.435 11.400 57.625 ;
        RECT 14.860 57.435 15.240 57.625 ;
        RECT 18.700 57.435 19.080 57.625 ;
        RECT 22.540 57.435 22.920 57.625 ;
        RECT 26.380 57.435 26.760 57.625 ;
        RECT 30.220 57.435 30.600 57.625 ;
        RECT 34.060 57.435 34.440 57.625 ;
        RECT 39.630 57.435 40.010 57.625 ;
        RECT 43.470 57.435 43.850 57.625 ;
        RECT 47.310 57.435 47.690 57.625 ;
        RECT 51.150 57.435 51.530 57.625 ;
        RECT 54.990 57.435 55.370 57.625 ;
        RECT 58.830 57.435 59.210 57.625 ;
        RECT 62.670 57.435 63.050 57.625 ;
        RECT 66.510 57.435 66.890 57.625 ;
        RECT 72.080 57.435 72.460 57.625 ;
        RECT 75.920 57.435 76.300 57.625 ;
        RECT 79.760 57.435 80.140 57.625 ;
        RECT 83.600 57.435 83.980 57.625 ;
        RECT 87.440 57.435 87.820 57.625 ;
        RECT 91.280 57.435 91.660 57.625 ;
        RECT 95.120 57.435 95.500 57.625 ;
        RECT 98.960 57.435 99.340 57.625 ;
        RECT 104.530 57.435 104.910 57.625 ;
        RECT 108.370 57.435 108.750 57.625 ;
        RECT 112.210 57.435 112.590 57.625 ;
        RECT 116.050 57.435 116.430 57.625 ;
        RECT 119.890 57.435 120.270 57.625 ;
        RECT 123.730 57.435 124.110 57.625 ;
        RECT 127.570 57.435 127.950 57.625 ;
        RECT 131.410 57.435 131.790 57.625 ;
        RECT 0.240 55.070 0.620 55.450 ;
        RECT 2.520 52.780 2.870 56.970 ;
        RECT 0.240 52.070 0.620 52.450 ;
        RECT 3.150 51.425 3.500 55.340 ;
        RECT 4.160 55.070 4.540 55.450 ;
        RECT 6.700 54.105 9.560 54.485 ;
        RECT 12.255 53.385 14.005 57.240 ;
        RECT 4.160 52.070 4.540 52.450 ;
        RECT 6.700 52.265 9.560 52.645 ;
        RECT 16.095 51.540 17.845 57.240 ;
        RECT 2.745 51.100 3.500 51.425 ;
        RECT 2.300 50.415 2.680 50.795 ;
        RECT 6.700 50.420 9.560 50.800 ;
        RECT 6.700 49.660 9.560 50.040 ;
        RECT 0.240 49.070 0.620 49.450 ;
        RECT 4.160 49.070 4.540 49.450 ;
        RECT 19.935 48.900 21.685 57.240 ;
        RECT 6.700 47.780 9.560 48.160 ;
        RECT 23.775 47.060 25.525 57.240 ;
        RECT 0.240 46.070 0.620 46.450 ;
        RECT 4.160 46.070 4.540 46.450 ;
        RECT 6.700 45.940 9.560 46.320 ;
        RECT 27.615 45.215 29.365 57.240 ;
        RECT 6.700 44.095 9.560 44.475 ;
        RECT 0.240 43.070 0.620 43.450 ;
        RECT 4.160 43.070 4.540 43.450 ;
        RECT 6.700 43.335 9.560 43.715 ;
        RECT 31.455 42.575 33.205 57.240 ;
        RECT 6.700 41.455 9.560 41.835 ;
        RECT 35.295 40.735 37.045 57.240 ;
        RECT 37.560 54.665 37.940 55.045 ;
        RECT 39.150 54.105 42.010 54.485 ;
        RECT 44.705 53.385 46.455 57.240 ;
        RECT 37.560 52.825 37.940 53.205 ;
        RECT 39.150 52.265 42.010 52.645 ;
        RECT 48.545 51.540 50.295 57.240 ;
        RECT 37.560 50.980 37.940 51.360 ;
        RECT 39.150 50.420 42.010 50.800 ;
        RECT 39.150 49.660 42.010 50.040 ;
        RECT 52.385 48.900 54.135 57.240 ;
        RECT 37.560 48.340 37.940 48.720 ;
        RECT 39.150 47.780 42.010 48.160 ;
        RECT 56.225 47.060 57.975 57.240 ;
        RECT 37.560 46.500 37.940 46.880 ;
        RECT 39.150 45.940 42.010 46.320 ;
        RECT 60.065 45.215 61.815 57.240 ;
        RECT 37.560 44.655 37.940 45.035 ;
        RECT 39.150 44.095 42.010 44.475 ;
        RECT 39.150 43.335 42.010 43.715 ;
        RECT 63.905 42.575 65.655 57.240 ;
        RECT 37.560 42.015 37.940 42.395 ;
        RECT 39.150 41.455 42.010 41.835 ;
        RECT 67.745 40.735 69.495 57.240 ;
        RECT 70.010 54.665 70.390 55.045 ;
        RECT 71.600 54.105 74.460 54.485 ;
        RECT 77.155 53.385 78.905 57.240 ;
        RECT 70.010 52.825 70.390 53.205 ;
        RECT 71.600 52.265 74.460 52.645 ;
        RECT 80.995 51.540 82.745 57.240 ;
        RECT 70.010 50.980 70.390 51.360 ;
        RECT 71.600 50.420 74.460 50.800 ;
        RECT 71.600 49.660 74.460 50.040 ;
        RECT 84.835 48.900 86.585 57.240 ;
        RECT 70.010 48.340 70.390 48.720 ;
        RECT 71.600 47.780 74.460 48.160 ;
        RECT 88.675 47.060 90.425 57.240 ;
        RECT 70.010 46.500 70.390 46.880 ;
        RECT 71.600 45.940 74.460 46.320 ;
        RECT 92.515 45.215 94.265 57.240 ;
        RECT 70.010 44.655 70.390 45.035 ;
        RECT 71.600 44.095 74.460 44.475 ;
        RECT 71.600 43.335 74.460 43.715 ;
        RECT 96.355 42.575 98.105 57.240 ;
        RECT 70.010 42.015 70.390 42.395 ;
        RECT 71.600 41.455 74.460 41.835 ;
        RECT 100.195 40.735 101.945 57.240 ;
        RECT 102.460 54.665 102.840 55.045 ;
        RECT 104.050 54.105 106.910 54.485 ;
        RECT 109.605 53.385 111.355 57.240 ;
        RECT 102.460 52.825 102.840 53.205 ;
        RECT 104.050 52.265 106.910 52.645 ;
        RECT 113.445 51.540 115.195 57.240 ;
        RECT 102.460 50.980 102.840 51.360 ;
        RECT 104.050 50.420 106.910 50.800 ;
        RECT 104.050 49.660 106.910 50.040 ;
        RECT 117.285 48.900 119.035 57.240 ;
        RECT 102.460 48.340 102.840 48.720 ;
        RECT 104.050 47.780 106.910 48.160 ;
        RECT 121.125 47.060 122.875 57.240 ;
        RECT 102.460 46.500 102.840 46.880 ;
        RECT 104.050 45.940 106.910 46.320 ;
        RECT 124.965 45.215 126.715 57.240 ;
        RECT 102.460 44.655 102.840 45.035 ;
        RECT 104.050 44.095 106.910 44.475 ;
        RECT 104.050 43.335 106.910 43.715 ;
        RECT 128.805 42.575 130.555 57.240 ;
        RECT 102.460 42.015 102.840 42.395 ;
        RECT 104.050 41.455 106.910 41.835 ;
        RECT 132.645 40.735 134.395 57.240 ;
        RECT 137.355 56.570 137.735 56.950 ;
        RECT 139.395 56.570 139.775 56.950 ;
        RECT 141.180 56.570 141.560 56.950 ;
        RECT 134.910 54.665 135.290 55.045 ;
        RECT 137.355 53.570 137.735 53.950 ;
        RECT 139.395 53.570 139.775 53.950 ;
        RECT 141.180 53.570 141.560 53.950 ;
        RECT 134.910 52.825 135.290 53.205 ;
        RECT 134.910 50.980 135.290 51.360 ;
        RECT 137.355 50.570 137.735 50.950 ;
        RECT 139.395 50.570 139.775 50.950 ;
        RECT 141.180 50.570 141.560 50.950 ;
        RECT 134.910 48.340 135.290 48.720 ;
        RECT 137.355 47.570 137.735 47.950 ;
        RECT 139.395 47.570 139.775 47.950 ;
        RECT 141.180 47.570 141.560 47.950 ;
        RECT 134.910 46.500 135.290 46.880 ;
        RECT 134.910 44.655 135.290 45.035 ;
        RECT 137.355 44.570 137.735 44.950 ;
        RECT 139.395 44.570 139.775 44.950 ;
        RECT 141.180 44.570 141.560 44.950 ;
        RECT 134.910 42.015 135.290 42.395 ;
        RECT 137.355 41.570 137.735 41.950 ;
        RECT 139.395 41.570 139.775 41.950 ;
        RECT 141.180 41.570 141.560 41.950 ;
        RECT 0.240 40.070 0.620 40.450 ;
        RECT 4.160 40.070 4.540 40.450 ;
        RECT 37.560 40.175 37.940 40.555 ;
        RECT 70.010 40.175 70.390 40.555 ;
        RECT 102.460 40.175 102.840 40.555 ;
        RECT 134.910 40.175 135.290 40.555 ;
        RECT 6.700 39.615 9.560 39.995 ;
        RECT 39.150 39.615 42.010 39.995 ;
        RECT 71.600 39.615 74.460 39.995 ;
        RECT 104.050 39.615 106.910 39.995 ;
        RECT 6.700 38.895 9.560 39.275 ;
        RECT 39.150 38.895 42.010 39.275 ;
        RECT 71.600 38.895 74.460 39.275 ;
        RECT 104.050 38.895 106.910 39.275 ;
        RECT 37.560 38.335 37.940 38.715 ;
        RECT 70.010 38.335 70.390 38.715 ;
        RECT 102.460 38.335 102.840 38.715 ;
        RECT 134.910 38.335 135.290 38.715 ;
        RECT 0.240 36.685 0.620 37.065 ;
        RECT 4.160 36.685 4.540 37.065 ;
        RECT 6.700 37.055 9.560 37.435 ;
        RECT 6.700 35.170 9.560 35.550 ;
        RECT 6.700 34.410 9.560 34.790 ;
        RECT 0.240 33.685 0.620 34.065 ;
        RECT 4.160 33.685 4.540 34.065 ;
        RECT 6.700 32.570 9.560 32.950 ;
        RECT 0.240 30.685 0.620 31.065 ;
        RECT 4.160 30.685 4.540 31.065 ;
        RECT 6.700 30.730 9.560 31.110 ;
        RECT 6.700 28.845 9.560 29.225 ;
        RECT 6.700 28.085 9.560 28.465 ;
        RECT 0.240 27.685 0.620 28.065 ;
        RECT 4.160 27.685 4.540 28.065 ;
        RECT 6.700 26.245 9.560 26.625 ;
        RECT 0.240 24.685 0.620 25.065 ;
        RECT 4.160 24.685 4.540 25.065 ;
        RECT 6.700 24.405 9.560 24.785 ;
        RECT 0.240 21.685 0.620 22.065 ;
        RECT 4.160 21.685 4.540 22.065 ;
        RECT 10.335 21.695 12.085 25.505 ;
        RECT 14.175 21.695 15.925 27.345 ;
        RECT 18.015 21.695 19.765 29.990 ;
        RECT 21.855 21.695 23.605 31.830 ;
        RECT 25.695 21.695 27.445 33.670 ;
        RECT 29.535 21.695 31.285 36.315 ;
        RECT 33.375 21.695 35.125 38.155 ;
        RECT 39.150 37.055 42.010 37.435 ;
        RECT 37.560 36.495 37.940 36.875 ;
        RECT 39.150 35.170 42.010 35.550 ;
        RECT 39.150 34.410 42.010 34.790 ;
        RECT 37.560 33.850 37.940 34.230 ;
        RECT 39.150 32.570 42.010 32.950 ;
        RECT 37.560 32.010 37.940 32.390 ;
        RECT 39.150 30.730 42.010 31.110 ;
        RECT 37.560 30.170 37.940 30.550 ;
        RECT 39.150 28.845 42.010 29.225 ;
        RECT 39.150 28.085 42.010 28.465 ;
        RECT 37.560 27.525 37.940 27.905 ;
        RECT 39.150 26.245 42.010 26.625 ;
        RECT 37.560 25.685 37.940 26.065 ;
        RECT 39.150 24.405 42.010 24.785 ;
        RECT 37.560 23.845 37.940 24.225 ;
        RECT 42.785 21.695 44.535 25.505 ;
        RECT 46.625 21.695 48.375 27.345 ;
        RECT 50.465 21.695 52.215 29.990 ;
        RECT 54.305 21.695 56.055 31.830 ;
        RECT 58.145 21.695 59.895 33.670 ;
        RECT 61.985 21.695 63.735 36.315 ;
        RECT 65.825 21.695 67.575 38.155 ;
        RECT 71.600 37.055 74.460 37.435 ;
        RECT 70.010 36.495 70.390 36.875 ;
        RECT 71.600 35.170 74.460 35.550 ;
        RECT 71.600 34.410 74.460 34.790 ;
        RECT 70.010 33.850 70.390 34.230 ;
        RECT 71.600 32.570 74.460 32.950 ;
        RECT 70.010 32.010 70.390 32.390 ;
        RECT 71.600 30.730 74.460 31.110 ;
        RECT 70.010 30.170 70.390 30.550 ;
        RECT 71.600 28.845 74.460 29.225 ;
        RECT 71.600 28.085 74.460 28.465 ;
        RECT 70.010 27.525 70.390 27.905 ;
        RECT 71.600 26.245 74.460 26.625 ;
        RECT 70.010 25.685 70.390 26.065 ;
        RECT 71.600 24.405 74.460 24.785 ;
        RECT 70.010 23.845 70.390 24.225 ;
        RECT 75.235 21.695 76.985 25.505 ;
        RECT 79.075 21.695 80.825 27.345 ;
        RECT 82.915 21.695 84.665 29.990 ;
        RECT 86.755 21.695 88.505 31.830 ;
        RECT 90.595 21.695 92.345 33.670 ;
        RECT 94.435 21.695 96.185 36.315 ;
        RECT 98.275 21.695 100.025 38.155 ;
        RECT 104.050 37.055 106.910 37.435 ;
        RECT 102.460 36.495 102.840 36.875 ;
        RECT 104.050 35.170 106.910 35.550 ;
        RECT 104.050 34.410 106.910 34.790 ;
        RECT 102.460 33.850 102.840 34.230 ;
        RECT 104.050 32.570 106.910 32.950 ;
        RECT 102.460 32.010 102.840 32.390 ;
        RECT 104.050 30.730 106.910 31.110 ;
        RECT 102.460 30.170 102.840 30.550 ;
        RECT 104.050 28.845 106.910 29.225 ;
        RECT 104.050 28.085 106.910 28.465 ;
        RECT 102.460 27.525 102.840 27.905 ;
        RECT 104.050 26.245 106.910 26.625 ;
        RECT 102.460 25.685 102.840 26.065 ;
        RECT 104.050 24.405 106.910 24.785 ;
        RECT 102.460 23.845 102.840 24.225 ;
        RECT 107.685 21.695 109.435 25.505 ;
        RECT 111.525 21.695 113.275 27.345 ;
        RECT 115.365 21.695 117.115 29.990 ;
        RECT 119.205 21.695 120.955 31.830 ;
        RECT 123.045 21.695 124.795 33.670 ;
        RECT 126.885 21.695 128.635 36.315 ;
        RECT 130.725 21.695 132.475 38.155 ;
        RECT 134.910 36.495 135.290 36.875 ;
        RECT 137.355 35.185 137.735 35.565 ;
        RECT 139.395 35.185 139.775 35.565 ;
        RECT 141.180 35.185 141.560 35.565 ;
        RECT 134.910 33.850 135.290 34.230 ;
        RECT 134.910 32.010 135.290 32.390 ;
        RECT 137.355 32.185 137.735 32.565 ;
        RECT 139.395 32.185 139.775 32.565 ;
        RECT 141.180 32.185 141.560 32.565 ;
        RECT 134.910 30.170 135.290 30.550 ;
        RECT 137.355 29.185 137.735 29.565 ;
        RECT 139.395 29.185 139.775 29.565 ;
        RECT 141.180 29.185 141.560 29.565 ;
        RECT 134.910 27.525 135.290 27.905 ;
        RECT 137.355 26.185 137.735 26.565 ;
        RECT 139.395 26.185 139.775 26.565 ;
        RECT 141.180 26.185 141.560 26.565 ;
        RECT 134.910 25.685 135.290 26.065 ;
        RECT 134.910 23.845 135.290 24.225 ;
        RECT 137.355 23.185 137.735 23.565 ;
        RECT 139.395 23.185 139.775 23.565 ;
        RECT 141.180 23.185 141.560 23.565 ;
        RECT 9.100 21.310 9.480 21.500 ;
        RECT 12.940 21.310 13.320 21.500 ;
        RECT 16.780 21.310 17.160 21.500 ;
        RECT 20.620 21.310 21.000 21.500 ;
        RECT 24.460 21.310 24.840 21.500 ;
        RECT 28.300 21.310 28.680 21.500 ;
        RECT 32.140 21.310 32.520 21.500 ;
        RECT 35.980 21.310 36.360 21.500 ;
        RECT 41.550 21.310 41.930 21.500 ;
        RECT 45.390 21.310 45.770 21.500 ;
        RECT 49.230 21.310 49.610 21.500 ;
        RECT 53.070 21.310 53.450 21.500 ;
        RECT 56.910 21.310 57.290 21.500 ;
        RECT 60.750 21.310 61.130 21.500 ;
        RECT 64.590 21.310 64.970 21.500 ;
        RECT 68.430 21.310 68.810 21.500 ;
        RECT 74.000 21.310 74.380 21.500 ;
        RECT 77.840 21.310 78.220 21.500 ;
        RECT 81.680 21.310 82.060 21.500 ;
        RECT 85.520 21.310 85.900 21.500 ;
        RECT 89.360 21.310 89.740 21.500 ;
        RECT 93.200 21.310 93.580 21.500 ;
        RECT 97.040 21.310 97.420 21.500 ;
        RECT 100.880 21.310 101.260 21.500 ;
        RECT 106.450 21.310 106.830 21.500 ;
        RECT 110.290 21.310 110.670 21.500 ;
        RECT 114.130 21.310 114.510 21.500 ;
        RECT 117.970 21.310 118.350 21.500 ;
        RECT 121.810 21.310 122.190 21.500 ;
        RECT 125.650 21.310 126.030 21.500 ;
        RECT 129.490 21.310 129.870 21.500 ;
        RECT 133.330 21.310 133.710 21.500 ;
        RECT 3.430 20.500 141.830 21.310 ;
        RECT 0.240 18.685 0.620 19.065 ;
        RECT 3.430 19.050 4.240 20.500 ;
        RECT 136.340 20.310 136.720 20.500 ;
        RECT 138.380 20.310 138.760 20.500 ;
        RECT 140.420 20.310 140.800 20.500 ;
        RECT 136.340 19.050 136.720 19.240 ;
        RECT 138.380 19.050 138.760 19.240 ;
        RECT 140.420 19.050 140.800 19.240 ;
        RECT 3.430 18.240 141.830 19.050 ;
        RECT 7.180 18.050 7.560 18.240 ;
        RECT 11.020 18.050 11.400 18.240 ;
        RECT 14.860 18.050 15.240 18.240 ;
        RECT 18.700 18.050 19.080 18.240 ;
        RECT 22.540 18.050 22.920 18.240 ;
        RECT 26.380 18.050 26.760 18.240 ;
        RECT 30.220 18.050 30.600 18.240 ;
        RECT 34.060 18.050 34.440 18.240 ;
        RECT 39.630 18.050 40.010 18.240 ;
        RECT 43.470 18.050 43.850 18.240 ;
        RECT 47.310 18.050 47.690 18.240 ;
        RECT 51.150 18.050 51.530 18.240 ;
        RECT 54.990 18.050 55.370 18.240 ;
        RECT 58.830 18.050 59.210 18.240 ;
        RECT 62.670 18.050 63.050 18.240 ;
        RECT 66.510 18.050 66.890 18.240 ;
        RECT 72.080 18.050 72.460 18.240 ;
        RECT 75.920 18.050 76.300 18.240 ;
        RECT 79.760 18.050 80.140 18.240 ;
        RECT 83.600 18.050 83.980 18.240 ;
        RECT 87.440 18.050 87.820 18.240 ;
        RECT 91.280 18.050 91.660 18.240 ;
        RECT 95.120 18.050 95.500 18.240 ;
        RECT 98.960 18.050 99.340 18.240 ;
        RECT 104.530 18.050 104.910 18.240 ;
        RECT 108.370 18.050 108.750 18.240 ;
        RECT 112.210 18.050 112.590 18.240 ;
        RECT 116.050 18.050 116.430 18.240 ;
        RECT 119.890 18.050 120.270 18.240 ;
        RECT 123.730 18.050 124.110 18.240 ;
        RECT 127.570 18.050 127.950 18.240 ;
        RECT 131.410 18.050 131.790 18.240 ;
        RECT 0.240 15.685 0.620 16.065 ;
        RECT 2.520 13.395 2.870 17.585 ;
        RECT 0.240 12.685 0.620 13.065 ;
        RECT 3.150 12.040 3.500 15.955 ;
        RECT 4.160 15.685 4.540 16.065 ;
        RECT 6.700 14.720 9.560 15.100 ;
        RECT 12.255 14.000 14.005 17.855 ;
        RECT 4.160 12.685 4.540 13.065 ;
        RECT 6.700 12.880 9.560 13.260 ;
        RECT 16.095 12.155 17.845 17.855 ;
        RECT 2.745 11.715 3.500 12.040 ;
        RECT 2.300 11.030 2.680 11.410 ;
        RECT 6.700 11.035 9.560 11.415 ;
        RECT 6.700 10.275 9.560 10.655 ;
        RECT 0.240 9.685 0.620 10.065 ;
        RECT 4.160 9.685 4.540 10.065 ;
        RECT 19.935 9.515 21.685 17.855 ;
        RECT 6.700 8.395 9.560 8.775 ;
        RECT 23.775 7.675 25.525 17.855 ;
        RECT 0.240 6.685 0.620 7.065 ;
        RECT 4.160 6.685 4.540 7.065 ;
        RECT 6.700 6.555 9.560 6.935 ;
        RECT 27.615 5.830 29.365 17.855 ;
        RECT 6.700 4.710 9.560 5.090 ;
        RECT 0.240 3.685 0.620 4.065 ;
        RECT 4.160 3.685 4.540 4.065 ;
        RECT 6.700 3.950 9.560 4.330 ;
        RECT 31.455 3.190 33.205 17.855 ;
        RECT 6.700 2.070 9.560 2.450 ;
        RECT 35.295 1.350 37.045 17.855 ;
        RECT 37.560 15.280 37.940 15.660 ;
        RECT 39.150 14.720 42.010 15.100 ;
        RECT 44.705 14.000 46.455 17.855 ;
        RECT 37.560 13.440 37.940 13.820 ;
        RECT 39.150 12.880 42.010 13.260 ;
        RECT 48.545 12.155 50.295 17.855 ;
        RECT 37.560 11.595 37.940 11.975 ;
        RECT 39.150 11.035 42.010 11.415 ;
        RECT 39.150 10.275 42.010 10.655 ;
        RECT 52.385 9.515 54.135 17.855 ;
        RECT 37.560 8.955 37.940 9.335 ;
        RECT 39.150 8.395 42.010 8.775 ;
        RECT 56.225 7.675 57.975 17.855 ;
        RECT 37.560 7.115 37.940 7.495 ;
        RECT 39.150 6.555 42.010 6.935 ;
        RECT 60.065 5.830 61.815 17.855 ;
        RECT 37.560 5.270 37.940 5.650 ;
        RECT 39.150 4.710 42.010 5.090 ;
        RECT 39.150 3.950 42.010 4.330 ;
        RECT 63.905 3.190 65.655 17.855 ;
        RECT 37.560 2.630 37.940 3.010 ;
        RECT 39.150 2.070 42.010 2.450 ;
        RECT 67.745 1.350 69.495 17.855 ;
        RECT 70.010 15.280 70.390 15.660 ;
        RECT 71.600 14.720 74.460 15.100 ;
        RECT 77.155 14.000 78.905 17.855 ;
        RECT 70.010 13.440 70.390 13.820 ;
        RECT 71.600 12.880 74.460 13.260 ;
        RECT 80.995 12.155 82.745 17.855 ;
        RECT 70.010 11.595 70.390 11.975 ;
        RECT 71.600 11.035 74.460 11.415 ;
        RECT 71.600 10.275 74.460 10.655 ;
        RECT 84.835 9.515 86.585 17.855 ;
        RECT 70.010 8.955 70.390 9.335 ;
        RECT 71.600 8.395 74.460 8.775 ;
        RECT 88.675 7.675 90.425 17.855 ;
        RECT 70.010 7.115 70.390 7.495 ;
        RECT 71.600 6.555 74.460 6.935 ;
        RECT 92.515 5.830 94.265 17.855 ;
        RECT 70.010 5.270 70.390 5.650 ;
        RECT 71.600 4.710 74.460 5.090 ;
        RECT 71.600 3.950 74.460 4.330 ;
        RECT 96.355 3.190 98.105 17.855 ;
        RECT 70.010 2.630 70.390 3.010 ;
        RECT 71.600 2.070 74.460 2.450 ;
        RECT 100.195 1.350 101.945 17.855 ;
        RECT 102.460 15.280 102.840 15.660 ;
        RECT 104.050 14.720 106.910 15.100 ;
        RECT 109.605 14.000 111.355 17.855 ;
        RECT 102.460 13.440 102.840 13.820 ;
        RECT 104.050 12.880 106.910 13.260 ;
        RECT 113.445 12.155 115.195 17.855 ;
        RECT 102.460 11.595 102.840 11.975 ;
        RECT 104.050 11.035 106.910 11.415 ;
        RECT 104.050 10.275 106.910 10.655 ;
        RECT 117.285 9.515 119.035 17.855 ;
        RECT 102.460 8.955 102.840 9.335 ;
        RECT 104.050 8.395 106.910 8.775 ;
        RECT 121.125 7.675 122.875 17.855 ;
        RECT 102.460 7.115 102.840 7.495 ;
        RECT 104.050 6.555 106.910 6.935 ;
        RECT 124.965 5.830 126.715 17.855 ;
        RECT 102.460 5.270 102.840 5.650 ;
        RECT 104.050 4.710 106.910 5.090 ;
        RECT 104.050 3.950 106.910 4.330 ;
        RECT 128.805 3.190 130.555 17.855 ;
        RECT 102.460 2.630 102.840 3.010 ;
        RECT 104.050 2.070 106.910 2.450 ;
        RECT 132.645 1.350 134.395 17.855 ;
        RECT 137.355 17.185 137.735 17.565 ;
        RECT 139.395 17.185 139.775 17.565 ;
        RECT 141.180 17.185 141.560 17.565 ;
        RECT 134.910 15.280 135.290 15.660 ;
        RECT 137.355 14.185 137.735 14.565 ;
        RECT 139.395 14.185 139.775 14.565 ;
        RECT 141.180 14.185 141.560 14.565 ;
        RECT 134.910 13.440 135.290 13.820 ;
        RECT 134.910 11.595 135.290 11.975 ;
        RECT 137.355 11.185 137.735 11.565 ;
        RECT 139.395 11.185 139.775 11.565 ;
        RECT 141.180 11.185 141.560 11.565 ;
        RECT 134.910 8.955 135.290 9.335 ;
        RECT 137.355 8.185 137.735 8.565 ;
        RECT 139.395 8.185 139.775 8.565 ;
        RECT 141.180 8.185 141.560 8.565 ;
        RECT 134.910 7.115 135.290 7.495 ;
        RECT 134.910 5.270 135.290 5.650 ;
        RECT 137.355 5.185 137.735 5.565 ;
        RECT 139.395 5.185 139.775 5.565 ;
        RECT 141.180 5.185 141.560 5.565 ;
        RECT 134.910 2.630 135.290 3.010 ;
        RECT 137.355 2.185 137.735 2.565 ;
        RECT 139.395 2.185 139.775 2.565 ;
        RECT 141.180 2.185 141.560 2.565 ;
        RECT 0.240 0.685 0.620 1.065 ;
        RECT 4.160 0.685 4.540 1.065 ;
        RECT 37.560 0.790 37.940 1.170 ;
        RECT 70.010 0.790 70.390 1.170 ;
        RECT 102.460 0.790 102.840 1.170 ;
        RECT 134.910 0.790 135.290 1.170 ;
        RECT 6.700 0.230 9.560 0.610 ;
        RECT 39.150 0.230 42.010 0.610 ;
        RECT 71.600 0.230 74.460 0.610 ;
        RECT 104.050 0.230 106.910 0.610 ;
      LAYER Metal3 ;
        RECT 6.700 314.590 9.560 314.970 ;
        RECT 39.150 314.590 42.010 314.970 ;
        RECT 71.600 314.590 74.460 314.970 ;
        RECT 104.050 314.590 106.910 314.970 ;
        RECT 28.740 314.360 29.120 314.410 ;
        RECT 37.560 314.360 37.940 314.410 ;
        RECT 28.740 314.080 37.940 314.360 ;
        RECT 28.740 314.030 29.120 314.080 ;
        RECT 37.560 314.030 37.940 314.080 ;
        RECT 61.190 314.360 61.570 314.410 ;
        RECT 70.010 314.360 70.390 314.410 ;
        RECT 61.190 314.080 70.390 314.360 ;
        RECT 61.190 314.030 61.570 314.080 ;
        RECT 70.010 314.030 70.390 314.080 ;
        RECT 93.640 314.360 94.020 314.410 ;
        RECT 102.460 314.360 102.840 314.410 ;
        RECT 93.640 314.080 102.840 314.360 ;
        RECT 93.640 314.030 94.020 314.080 ;
        RECT 102.460 314.030 102.840 314.080 ;
        RECT 126.090 314.360 126.470 314.410 ;
        RECT 134.910 314.360 135.290 314.410 ;
        RECT 126.090 314.080 135.290 314.360 ;
        RECT 126.090 314.030 126.470 314.080 ;
        RECT 134.910 314.030 135.290 314.080 ;
        RECT 0.240 312.380 0.620 312.760 ;
        RECT 4.160 312.380 4.540 312.760 ;
        RECT 6.700 312.750 9.560 313.130 ;
        RECT 39.150 312.750 42.010 313.130 ;
        RECT 71.600 312.750 74.460 313.130 ;
        RECT 104.050 312.750 106.910 313.130 ;
        RECT 30.020 312.520 30.400 312.570 ;
        RECT 37.560 312.520 37.940 312.570 ;
        RECT 30.020 312.240 37.940 312.520 ;
        RECT 30.020 312.190 30.400 312.240 ;
        RECT 37.560 312.190 37.940 312.240 ;
        RECT 62.470 312.520 62.850 312.570 ;
        RECT 70.010 312.520 70.390 312.570 ;
        RECT 62.470 312.240 70.390 312.520 ;
        RECT 62.470 312.190 62.850 312.240 ;
        RECT 70.010 312.190 70.390 312.240 ;
        RECT 94.920 312.520 95.300 312.570 ;
        RECT 102.460 312.520 102.840 312.570 ;
        RECT 94.920 312.240 102.840 312.520 ;
        RECT 94.920 312.190 95.300 312.240 ;
        RECT 102.460 312.190 102.840 312.240 ;
        RECT 127.370 312.520 127.750 312.570 ;
        RECT 134.910 312.520 135.290 312.570 ;
        RECT 127.370 312.240 135.290 312.520 ;
        RECT 127.370 312.190 127.750 312.240 ;
        RECT 134.910 312.190 135.290 312.240 ;
        RECT 6.700 310.865 9.560 311.245 ;
        RECT 39.150 310.865 42.010 311.245 ;
        RECT 71.600 310.865 74.460 311.245 ;
        RECT 104.050 310.865 106.910 311.245 ;
        RECT 137.355 310.880 137.735 311.260 ;
        RECT 139.395 310.880 139.775 311.260 ;
        RECT 141.180 310.880 141.560 311.260 ;
        RECT 6.700 310.105 9.560 310.485 ;
        RECT 39.150 310.105 42.010 310.485 ;
        RECT 71.600 310.105 74.460 310.485 ;
        RECT 104.050 310.105 106.910 310.485 ;
        RECT 31.300 309.875 31.680 309.925 ;
        RECT 37.560 309.875 37.940 309.925 ;
        RECT 0.240 309.380 0.620 309.760 ;
        RECT 4.160 309.380 4.540 309.760 ;
        RECT 31.300 309.595 37.940 309.875 ;
        RECT 31.300 309.545 31.680 309.595 ;
        RECT 37.560 309.545 37.940 309.595 ;
        RECT 63.750 309.875 64.130 309.925 ;
        RECT 70.010 309.875 70.390 309.925 ;
        RECT 63.750 309.595 70.390 309.875 ;
        RECT 63.750 309.545 64.130 309.595 ;
        RECT 70.010 309.545 70.390 309.595 ;
        RECT 96.200 309.875 96.580 309.925 ;
        RECT 102.460 309.875 102.840 309.925 ;
        RECT 96.200 309.595 102.840 309.875 ;
        RECT 96.200 309.545 96.580 309.595 ;
        RECT 102.460 309.545 102.840 309.595 ;
        RECT 128.650 309.875 129.030 309.925 ;
        RECT 134.910 309.875 135.290 309.925 ;
        RECT 128.650 309.595 135.290 309.875 ;
        RECT 128.650 309.545 129.030 309.595 ;
        RECT 134.910 309.545 135.290 309.595 ;
        RECT 6.700 308.265 9.560 308.645 ;
        RECT 39.150 308.265 42.010 308.645 ;
        RECT 71.600 308.265 74.460 308.645 ;
        RECT 104.050 308.265 106.910 308.645 ;
        RECT 32.580 308.035 32.960 308.085 ;
        RECT 37.560 308.035 37.940 308.085 ;
        RECT 32.580 307.755 37.940 308.035 ;
        RECT 32.580 307.705 32.960 307.755 ;
        RECT 37.560 307.705 37.940 307.755 ;
        RECT 65.030 308.035 65.410 308.085 ;
        RECT 70.010 308.035 70.390 308.085 ;
        RECT 65.030 307.755 70.390 308.035 ;
        RECT 65.030 307.705 65.410 307.755 ;
        RECT 70.010 307.705 70.390 307.755 ;
        RECT 97.480 308.035 97.860 308.085 ;
        RECT 102.460 308.035 102.840 308.085 ;
        RECT 97.480 307.755 102.840 308.035 ;
        RECT 97.480 307.705 97.860 307.755 ;
        RECT 102.460 307.705 102.840 307.755 ;
        RECT 129.930 308.035 130.310 308.085 ;
        RECT 134.910 308.035 135.290 308.085 ;
        RECT 129.930 307.755 135.290 308.035 ;
        RECT 137.355 307.880 137.735 308.260 ;
        RECT 139.395 307.880 139.775 308.260 ;
        RECT 141.180 307.880 141.560 308.260 ;
        RECT 129.930 307.705 130.310 307.755 ;
        RECT 134.910 307.705 135.290 307.755 ;
        RECT 0.240 306.380 0.620 306.760 ;
        RECT 4.160 306.380 4.540 306.760 ;
        RECT 6.700 306.425 9.560 306.805 ;
        RECT 39.150 306.425 42.010 306.805 ;
        RECT 71.600 306.425 74.460 306.805 ;
        RECT 104.050 306.425 106.910 306.805 ;
        RECT 33.860 306.195 34.240 306.245 ;
        RECT 37.560 306.195 37.940 306.245 ;
        RECT 33.860 305.915 37.940 306.195 ;
        RECT 33.860 305.865 34.240 305.915 ;
        RECT 37.560 305.865 37.940 305.915 ;
        RECT 66.310 306.195 66.690 306.245 ;
        RECT 70.010 306.195 70.390 306.245 ;
        RECT 66.310 305.915 70.390 306.195 ;
        RECT 66.310 305.865 66.690 305.915 ;
        RECT 70.010 305.865 70.390 305.915 ;
        RECT 98.760 306.195 99.140 306.245 ;
        RECT 102.460 306.195 102.840 306.245 ;
        RECT 98.760 305.915 102.840 306.195 ;
        RECT 98.760 305.865 99.140 305.915 ;
        RECT 102.460 305.865 102.840 305.915 ;
        RECT 131.210 306.195 131.590 306.245 ;
        RECT 134.910 306.195 135.290 306.245 ;
        RECT 131.210 305.915 135.290 306.195 ;
        RECT 131.210 305.865 131.590 305.915 ;
        RECT 134.910 305.865 135.290 305.915 ;
        RECT 6.700 304.540 9.560 304.920 ;
        RECT 39.150 304.540 42.010 304.920 ;
        RECT 71.600 304.540 74.460 304.920 ;
        RECT 104.050 304.540 106.910 304.920 ;
        RECT 137.355 304.880 137.735 305.260 ;
        RECT 139.395 304.880 139.775 305.260 ;
        RECT 141.180 304.880 141.560 305.260 ;
        RECT 6.700 303.780 9.560 304.160 ;
        RECT 39.150 303.780 42.010 304.160 ;
        RECT 71.600 303.780 74.460 304.160 ;
        RECT 104.050 303.780 106.910 304.160 ;
        RECT 0.240 303.380 0.620 303.760 ;
        RECT 4.160 303.380 4.540 303.760 ;
        RECT 35.140 303.550 35.520 303.600 ;
        RECT 37.560 303.550 37.940 303.600 ;
        RECT 35.140 303.270 37.940 303.550 ;
        RECT 35.140 303.220 35.520 303.270 ;
        RECT 37.560 303.220 37.940 303.270 ;
        RECT 67.590 303.550 67.970 303.600 ;
        RECT 70.010 303.550 70.390 303.600 ;
        RECT 67.590 303.270 70.390 303.550 ;
        RECT 67.590 303.220 67.970 303.270 ;
        RECT 70.010 303.220 70.390 303.270 ;
        RECT 100.040 303.550 100.420 303.600 ;
        RECT 102.460 303.550 102.840 303.600 ;
        RECT 100.040 303.270 102.840 303.550 ;
        RECT 100.040 303.220 100.420 303.270 ;
        RECT 102.460 303.220 102.840 303.270 ;
        RECT 132.490 303.550 132.870 303.600 ;
        RECT 134.910 303.550 135.290 303.600 ;
        RECT 132.490 303.270 135.290 303.550 ;
        RECT 132.490 303.220 132.870 303.270 ;
        RECT 134.910 303.220 135.290 303.270 ;
        RECT 6.700 301.940 9.560 302.320 ;
        RECT 39.150 301.940 42.010 302.320 ;
        RECT 71.600 301.940 74.460 302.320 ;
        RECT 104.050 301.940 106.910 302.320 ;
        RECT 137.355 301.880 137.735 302.260 ;
        RECT 139.395 301.880 139.775 302.260 ;
        RECT 141.180 301.880 141.560 302.260 ;
        RECT 36.420 301.710 36.800 301.760 ;
        RECT 37.560 301.710 37.940 301.760 ;
        RECT 36.420 301.430 37.940 301.710 ;
        RECT 36.420 301.380 36.800 301.430 ;
        RECT 37.560 301.380 37.940 301.430 ;
        RECT 68.870 301.710 69.250 301.760 ;
        RECT 70.010 301.710 70.390 301.760 ;
        RECT 68.870 301.430 70.390 301.710 ;
        RECT 68.870 301.380 69.250 301.430 ;
        RECT 70.010 301.380 70.390 301.430 ;
        RECT 101.320 301.710 101.700 301.760 ;
        RECT 102.460 301.710 102.840 301.760 ;
        RECT 101.320 301.430 102.840 301.710 ;
        RECT 101.320 301.380 101.700 301.430 ;
        RECT 102.460 301.380 102.840 301.430 ;
        RECT 133.770 301.710 134.150 301.760 ;
        RECT 134.910 301.710 135.290 301.760 ;
        RECT 133.770 301.430 135.290 301.710 ;
        RECT 133.770 301.380 134.150 301.430 ;
        RECT 134.910 301.380 135.290 301.430 ;
        RECT 0.240 300.380 0.620 300.760 ;
        RECT 4.160 300.380 4.540 300.760 ;
        RECT 6.700 300.100 9.560 300.480 ;
        RECT 39.150 300.100 42.010 300.480 ;
        RECT 71.600 300.100 74.460 300.480 ;
        RECT 104.050 300.100 106.910 300.480 ;
        RECT 37.560 299.540 38.080 299.920 ;
        RECT 70.010 299.540 70.530 299.920 ;
        RECT 102.460 299.540 102.980 299.920 ;
        RECT 134.910 299.540 135.430 299.920 ;
        RECT 137.355 298.880 137.735 299.260 ;
        RECT 139.395 298.880 139.775 299.260 ;
        RECT 141.180 298.880 141.560 299.260 ;
        RECT 0.240 297.380 0.620 297.760 ;
        RECT 4.160 297.380 4.540 297.760 ;
        RECT 0.240 294.380 0.620 294.760 ;
        RECT 137.355 292.880 137.735 293.260 ;
        RECT 139.395 292.880 139.775 293.260 ;
        RECT 141.180 292.880 141.560 293.260 ;
        RECT 0.240 291.380 0.620 291.760 ;
        RECT 4.160 291.380 4.540 291.760 ;
        RECT 37.060 290.975 37.940 291.355 ;
        RECT 69.510 290.975 70.390 291.355 ;
        RECT 101.960 290.975 102.840 291.355 ;
        RECT 134.410 290.975 135.290 291.355 ;
        RECT 6.700 290.415 9.560 290.795 ;
        RECT 39.150 290.415 42.010 290.795 ;
        RECT 71.600 290.415 74.460 290.795 ;
        RECT 104.050 290.415 106.910 290.795 ;
        RECT 137.355 289.880 137.735 290.260 ;
        RECT 139.395 289.880 139.775 290.260 ;
        RECT 141.180 289.880 141.560 290.260 ;
        RECT 35.780 289.465 36.160 289.515 ;
        RECT 37.560 289.465 37.940 289.515 ;
        RECT 35.780 289.185 37.940 289.465 ;
        RECT 35.780 289.135 36.160 289.185 ;
        RECT 37.560 289.135 37.940 289.185 ;
        RECT 68.230 289.465 68.610 289.515 ;
        RECT 70.010 289.465 70.390 289.515 ;
        RECT 68.230 289.185 70.390 289.465 ;
        RECT 68.230 289.135 68.610 289.185 ;
        RECT 70.010 289.135 70.390 289.185 ;
        RECT 100.680 289.465 101.060 289.515 ;
        RECT 102.460 289.465 102.840 289.515 ;
        RECT 100.680 289.185 102.840 289.465 ;
        RECT 100.680 289.135 101.060 289.185 ;
        RECT 102.460 289.135 102.840 289.185 ;
        RECT 133.130 289.465 133.510 289.515 ;
        RECT 134.910 289.465 135.290 289.515 ;
        RECT 133.130 289.185 135.290 289.465 ;
        RECT 133.130 289.135 133.510 289.185 ;
        RECT 134.910 289.135 135.290 289.185 ;
        RECT 0.240 288.380 0.620 288.760 ;
        RECT 4.160 288.380 4.540 288.760 ;
        RECT 6.700 288.575 9.560 288.955 ;
        RECT 39.150 288.575 42.010 288.955 ;
        RECT 71.600 288.575 74.460 288.955 ;
        RECT 104.050 288.575 106.910 288.955 ;
        RECT 34.500 287.620 34.880 287.670 ;
        RECT 37.560 287.620 37.940 287.670 ;
        RECT 34.500 287.340 37.940 287.620 ;
        RECT 34.500 287.290 34.880 287.340 ;
        RECT 37.560 287.290 37.940 287.340 ;
        RECT 66.950 287.620 67.330 287.670 ;
        RECT 70.010 287.620 70.390 287.670 ;
        RECT 66.950 287.340 70.390 287.620 ;
        RECT 66.950 287.290 67.330 287.340 ;
        RECT 70.010 287.290 70.390 287.340 ;
        RECT 99.400 287.620 99.780 287.670 ;
        RECT 102.460 287.620 102.840 287.670 ;
        RECT 99.400 287.340 102.840 287.620 ;
        RECT 99.400 287.290 99.780 287.340 ;
        RECT 102.460 287.290 102.840 287.340 ;
        RECT 131.850 287.620 132.230 287.670 ;
        RECT 134.910 287.620 135.290 287.670 ;
        RECT 131.850 287.340 135.290 287.620 ;
        RECT 131.850 287.290 132.230 287.340 ;
        RECT 134.910 287.290 135.290 287.340 ;
        RECT 6.700 286.730 9.560 287.110 ;
        RECT 39.150 286.730 42.010 287.110 ;
        RECT 71.600 286.730 74.460 287.110 ;
        RECT 104.050 286.730 106.910 287.110 ;
        RECT 137.355 286.880 137.735 287.260 ;
        RECT 139.395 286.880 139.775 287.260 ;
        RECT 141.180 286.880 141.560 287.260 ;
        RECT 6.700 285.970 9.560 286.350 ;
        RECT 39.150 285.970 42.010 286.350 ;
        RECT 71.600 285.970 74.460 286.350 ;
        RECT 104.050 285.970 106.910 286.350 ;
        RECT 0.240 285.380 0.620 285.760 ;
        RECT 4.160 285.380 4.540 285.760 ;
        RECT 33.220 284.980 33.600 285.030 ;
        RECT 37.560 284.980 37.940 285.030 ;
        RECT 33.220 284.700 37.940 284.980 ;
        RECT 33.220 284.650 33.600 284.700 ;
        RECT 37.560 284.650 37.940 284.700 ;
        RECT 65.670 284.980 66.050 285.030 ;
        RECT 70.010 284.980 70.390 285.030 ;
        RECT 65.670 284.700 70.390 284.980 ;
        RECT 65.670 284.650 66.050 284.700 ;
        RECT 70.010 284.650 70.390 284.700 ;
        RECT 98.120 284.980 98.500 285.030 ;
        RECT 102.460 284.980 102.840 285.030 ;
        RECT 98.120 284.700 102.840 284.980 ;
        RECT 98.120 284.650 98.500 284.700 ;
        RECT 102.460 284.650 102.840 284.700 ;
        RECT 130.570 284.980 130.950 285.030 ;
        RECT 134.910 284.980 135.290 285.030 ;
        RECT 130.570 284.700 135.290 284.980 ;
        RECT 130.570 284.650 130.950 284.700 ;
        RECT 134.910 284.650 135.290 284.700 ;
        RECT 6.700 284.090 9.560 284.470 ;
        RECT 39.150 284.090 42.010 284.470 ;
        RECT 71.600 284.090 74.460 284.470 ;
        RECT 104.050 284.090 106.910 284.470 ;
        RECT 137.355 283.880 137.735 284.260 ;
        RECT 139.395 283.880 139.775 284.260 ;
        RECT 141.180 283.880 141.560 284.260 ;
        RECT 31.940 283.140 32.320 283.190 ;
        RECT 37.560 283.140 37.940 283.190 ;
        RECT 31.940 282.860 37.940 283.140 ;
        RECT 31.940 282.810 32.320 282.860 ;
        RECT 37.560 282.810 37.940 282.860 ;
        RECT 64.390 283.140 64.770 283.190 ;
        RECT 70.010 283.140 70.390 283.190 ;
        RECT 64.390 282.860 70.390 283.140 ;
        RECT 64.390 282.810 64.770 282.860 ;
        RECT 70.010 282.810 70.390 282.860 ;
        RECT 96.840 283.140 97.220 283.190 ;
        RECT 102.460 283.140 102.840 283.190 ;
        RECT 96.840 282.860 102.840 283.140 ;
        RECT 96.840 282.810 97.220 282.860 ;
        RECT 102.460 282.810 102.840 282.860 ;
        RECT 129.290 283.140 129.670 283.190 ;
        RECT 134.910 283.140 135.290 283.190 ;
        RECT 129.290 282.860 135.290 283.140 ;
        RECT 129.290 282.810 129.670 282.860 ;
        RECT 134.910 282.810 135.290 282.860 ;
        RECT 0.240 282.380 0.620 282.760 ;
        RECT 4.160 282.380 4.540 282.760 ;
        RECT 6.700 282.250 9.560 282.630 ;
        RECT 39.150 282.250 42.010 282.630 ;
        RECT 71.600 282.250 74.460 282.630 ;
        RECT 104.050 282.250 106.910 282.630 ;
        RECT 30.660 281.295 31.040 281.345 ;
        RECT 37.560 281.295 37.940 281.345 ;
        RECT 30.660 281.015 37.940 281.295 ;
        RECT 30.660 280.965 31.040 281.015 ;
        RECT 37.560 280.965 37.940 281.015 ;
        RECT 63.110 281.295 63.490 281.345 ;
        RECT 70.010 281.295 70.390 281.345 ;
        RECT 63.110 281.015 70.390 281.295 ;
        RECT 63.110 280.965 63.490 281.015 ;
        RECT 70.010 280.965 70.390 281.015 ;
        RECT 95.560 281.295 95.940 281.345 ;
        RECT 102.460 281.295 102.840 281.345 ;
        RECT 95.560 281.015 102.840 281.295 ;
        RECT 95.560 280.965 95.940 281.015 ;
        RECT 102.460 280.965 102.840 281.015 ;
        RECT 128.010 281.295 128.390 281.345 ;
        RECT 134.910 281.295 135.290 281.345 ;
        RECT 128.010 281.015 135.290 281.295 ;
        RECT 128.010 280.965 128.390 281.015 ;
        RECT 134.910 280.965 135.290 281.015 ;
        RECT 137.355 280.880 137.735 281.260 ;
        RECT 139.395 280.880 139.775 281.260 ;
        RECT 141.180 280.880 141.560 281.260 ;
        RECT 6.700 280.405 9.560 280.785 ;
        RECT 39.150 280.405 42.010 280.785 ;
        RECT 71.600 280.405 74.460 280.785 ;
        RECT 104.050 280.405 106.910 280.785 ;
        RECT 0.240 279.380 0.620 279.760 ;
        RECT 4.160 279.380 4.540 279.760 ;
        RECT 6.700 279.645 9.560 280.025 ;
        RECT 39.150 279.645 42.010 280.025 ;
        RECT 71.600 279.645 74.460 280.025 ;
        RECT 104.050 279.645 106.910 280.025 ;
        RECT 29.380 278.655 29.760 278.705 ;
        RECT 37.560 278.655 37.940 278.705 ;
        RECT 29.380 278.375 37.940 278.655 ;
        RECT 29.380 278.325 29.760 278.375 ;
        RECT 37.560 278.325 37.940 278.375 ;
        RECT 61.830 278.655 62.210 278.705 ;
        RECT 70.010 278.655 70.390 278.705 ;
        RECT 61.830 278.375 70.390 278.655 ;
        RECT 61.830 278.325 62.210 278.375 ;
        RECT 70.010 278.325 70.390 278.375 ;
        RECT 94.280 278.655 94.660 278.705 ;
        RECT 102.460 278.655 102.840 278.705 ;
        RECT 94.280 278.375 102.840 278.655 ;
        RECT 94.280 278.325 94.660 278.375 ;
        RECT 102.460 278.325 102.840 278.375 ;
        RECT 126.730 278.655 127.110 278.705 ;
        RECT 134.910 278.655 135.290 278.705 ;
        RECT 126.730 278.375 135.290 278.655 ;
        RECT 126.730 278.325 127.110 278.375 ;
        RECT 134.910 278.325 135.290 278.375 ;
        RECT 6.700 277.765 9.560 278.145 ;
        RECT 39.150 277.765 42.010 278.145 ;
        RECT 71.600 277.765 74.460 278.145 ;
        RECT 104.050 277.765 106.910 278.145 ;
        RECT 137.355 277.880 137.735 278.260 ;
        RECT 139.395 277.880 139.775 278.260 ;
        RECT 141.180 277.880 141.560 278.260 ;
        RECT 28.100 276.815 28.480 276.865 ;
        RECT 37.560 276.815 37.940 276.865 ;
        RECT 0.240 276.380 0.620 276.760 ;
        RECT 4.160 276.380 4.540 276.760 ;
        RECT 28.100 276.535 37.940 276.815 ;
        RECT 28.100 276.485 28.480 276.535 ;
        RECT 37.560 276.485 37.940 276.535 ;
        RECT 60.550 276.815 60.930 276.865 ;
        RECT 70.010 276.815 70.390 276.865 ;
        RECT 60.550 276.535 70.390 276.815 ;
        RECT 60.550 276.485 60.930 276.535 ;
        RECT 70.010 276.485 70.390 276.535 ;
        RECT 93.000 276.815 93.380 276.865 ;
        RECT 102.460 276.815 102.840 276.865 ;
        RECT 93.000 276.535 102.840 276.815 ;
        RECT 93.000 276.485 93.380 276.535 ;
        RECT 102.460 276.485 102.840 276.535 ;
        RECT 125.450 276.815 125.830 276.865 ;
        RECT 134.910 276.815 135.290 276.865 ;
        RECT 125.450 276.535 135.290 276.815 ;
        RECT 125.450 276.485 125.830 276.535 ;
        RECT 134.910 276.485 135.290 276.535 ;
        RECT 6.700 275.925 9.560 276.305 ;
        RECT 39.150 275.925 42.010 276.305 ;
        RECT 71.600 275.925 74.460 276.305 ;
        RECT 104.050 275.925 106.910 276.305 ;
        RECT 6.700 275.205 9.560 275.585 ;
        RECT 39.150 275.205 42.010 275.585 ;
        RECT 71.600 275.205 74.460 275.585 ;
        RECT 104.050 275.205 106.910 275.585 ;
        RECT 28.740 274.975 29.120 275.025 ;
        RECT 37.560 274.975 37.940 275.025 ;
        RECT 28.740 274.695 37.940 274.975 ;
        RECT 28.740 274.645 29.120 274.695 ;
        RECT 37.560 274.645 37.940 274.695 ;
        RECT 61.190 274.975 61.570 275.025 ;
        RECT 70.010 274.975 70.390 275.025 ;
        RECT 61.190 274.695 70.390 274.975 ;
        RECT 61.190 274.645 61.570 274.695 ;
        RECT 70.010 274.645 70.390 274.695 ;
        RECT 93.640 274.975 94.020 275.025 ;
        RECT 102.460 274.975 102.840 275.025 ;
        RECT 93.640 274.695 102.840 274.975 ;
        RECT 93.640 274.645 94.020 274.695 ;
        RECT 102.460 274.645 102.840 274.695 ;
        RECT 126.090 274.975 126.470 275.025 ;
        RECT 134.910 274.975 135.290 275.025 ;
        RECT 126.090 274.695 135.290 274.975 ;
        RECT 126.090 274.645 126.470 274.695 ;
        RECT 134.910 274.645 135.290 274.695 ;
        RECT 0.240 272.995 0.620 273.375 ;
        RECT 4.160 272.995 4.540 273.375 ;
        RECT 6.700 273.365 9.560 273.745 ;
        RECT 39.150 273.365 42.010 273.745 ;
        RECT 71.600 273.365 74.460 273.745 ;
        RECT 104.050 273.365 106.910 273.745 ;
        RECT 30.020 273.135 30.400 273.185 ;
        RECT 37.560 273.135 37.940 273.185 ;
        RECT 30.020 272.855 37.940 273.135 ;
        RECT 30.020 272.805 30.400 272.855 ;
        RECT 37.560 272.805 37.940 272.855 ;
        RECT 62.470 273.135 62.850 273.185 ;
        RECT 70.010 273.135 70.390 273.185 ;
        RECT 62.470 272.855 70.390 273.135 ;
        RECT 62.470 272.805 62.850 272.855 ;
        RECT 70.010 272.805 70.390 272.855 ;
        RECT 94.920 273.135 95.300 273.185 ;
        RECT 102.460 273.135 102.840 273.185 ;
        RECT 94.920 272.855 102.840 273.135 ;
        RECT 94.920 272.805 95.300 272.855 ;
        RECT 102.460 272.805 102.840 272.855 ;
        RECT 127.370 273.135 127.750 273.185 ;
        RECT 134.910 273.135 135.290 273.185 ;
        RECT 127.370 272.855 135.290 273.135 ;
        RECT 127.370 272.805 127.750 272.855 ;
        RECT 134.910 272.805 135.290 272.855 ;
        RECT 6.700 271.480 9.560 271.860 ;
        RECT 39.150 271.480 42.010 271.860 ;
        RECT 71.600 271.480 74.460 271.860 ;
        RECT 104.050 271.480 106.910 271.860 ;
        RECT 137.355 271.495 137.735 271.875 ;
        RECT 139.395 271.495 139.775 271.875 ;
        RECT 141.180 271.495 141.560 271.875 ;
        RECT 6.700 270.720 9.560 271.100 ;
        RECT 39.150 270.720 42.010 271.100 ;
        RECT 71.600 270.720 74.460 271.100 ;
        RECT 104.050 270.720 106.910 271.100 ;
        RECT 31.300 270.490 31.680 270.540 ;
        RECT 37.560 270.490 37.940 270.540 ;
        RECT 0.240 269.995 0.620 270.375 ;
        RECT 4.160 269.995 4.540 270.375 ;
        RECT 31.300 270.210 37.940 270.490 ;
        RECT 31.300 270.160 31.680 270.210 ;
        RECT 37.560 270.160 37.940 270.210 ;
        RECT 63.750 270.490 64.130 270.540 ;
        RECT 70.010 270.490 70.390 270.540 ;
        RECT 63.750 270.210 70.390 270.490 ;
        RECT 63.750 270.160 64.130 270.210 ;
        RECT 70.010 270.160 70.390 270.210 ;
        RECT 96.200 270.490 96.580 270.540 ;
        RECT 102.460 270.490 102.840 270.540 ;
        RECT 96.200 270.210 102.840 270.490 ;
        RECT 96.200 270.160 96.580 270.210 ;
        RECT 102.460 270.160 102.840 270.210 ;
        RECT 128.650 270.490 129.030 270.540 ;
        RECT 134.910 270.490 135.290 270.540 ;
        RECT 128.650 270.210 135.290 270.490 ;
        RECT 128.650 270.160 129.030 270.210 ;
        RECT 134.910 270.160 135.290 270.210 ;
        RECT 6.700 268.880 9.560 269.260 ;
        RECT 39.150 268.880 42.010 269.260 ;
        RECT 71.600 268.880 74.460 269.260 ;
        RECT 104.050 268.880 106.910 269.260 ;
        RECT 32.580 268.650 32.960 268.700 ;
        RECT 37.560 268.650 37.940 268.700 ;
        RECT 32.580 268.370 37.940 268.650 ;
        RECT 32.580 268.320 32.960 268.370 ;
        RECT 37.560 268.320 37.940 268.370 ;
        RECT 65.030 268.650 65.410 268.700 ;
        RECT 70.010 268.650 70.390 268.700 ;
        RECT 65.030 268.370 70.390 268.650 ;
        RECT 65.030 268.320 65.410 268.370 ;
        RECT 70.010 268.320 70.390 268.370 ;
        RECT 97.480 268.650 97.860 268.700 ;
        RECT 102.460 268.650 102.840 268.700 ;
        RECT 97.480 268.370 102.840 268.650 ;
        RECT 97.480 268.320 97.860 268.370 ;
        RECT 102.460 268.320 102.840 268.370 ;
        RECT 129.930 268.650 130.310 268.700 ;
        RECT 134.910 268.650 135.290 268.700 ;
        RECT 129.930 268.370 135.290 268.650 ;
        RECT 137.355 268.495 137.735 268.875 ;
        RECT 139.395 268.495 139.775 268.875 ;
        RECT 141.180 268.495 141.560 268.875 ;
        RECT 129.930 268.320 130.310 268.370 ;
        RECT 134.910 268.320 135.290 268.370 ;
        RECT 0.240 266.995 0.620 267.375 ;
        RECT 4.160 266.995 4.540 267.375 ;
        RECT 6.700 267.040 9.560 267.420 ;
        RECT 39.150 267.040 42.010 267.420 ;
        RECT 71.600 267.040 74.460 267.420 ;
        RECT 104.050 267.040 106.910 267.420 ;
        RECT 33.860 266.810 34.240 266.860 ;
        RECT 37.560 266.810 37.940 266.860 ;
        RECT 33.860 266.530 37.940 266.810 ;
        RECT 33.860 266.480 34.240 266.530 ;
        RECT 37.560 266.480 37.940 266.530 ;
        RECT 66.310 266.810 66.690 266.860 ;
        RECT 70.010 266.810 70.390 266.860 ;
        RECT 66.310 266.530 70.390 266.810 ;
        RECT 66.310 266.480 66.690 266.530 ;
        RECT 70.010 266.480 70.390 266.530 ;
        RECT 98.760 266.810 99.140 266.860 ;
        RECT 102.460 266.810 102.840 266.860 ;
        RECT 98.760 266.530 102.840 266.810 ;
        RECT 98.760 266.480 99.140 266.530 ;
        RECT 102.460 266.480 102.840 266.530 ;
        RECT 131.210 266.810 131.590 266.860 ;
        RECT 134.910 266.810 135.290 266.860 ;
        RECT 131.210 266.530 135.290 266.810 ;
        RECT 131.210 266.480 131.590 266.530 ;
        RECT 134.910 266.480 135.290 266.530 ;
        RECT 6.700 265.155 9.560 265.535 ;
        RECT 39.150 265.155 42.010 265.535 ;
        RECT 71.600 265.155 74.460 265.535 ;
        RECT 104.050 265.155 106.910 265.535 ;
        RECT 137.355 265.495 137.735 265.875 ;
        RECT 139.395 265.495 139.775 265.875 ;
        RECT 141.180 265.495 141.560 265.875 ;
        RECT 6.700 264.395 9.560 264.775 ;
        RECT 39.150 264.395 42.010 264.775 ;
        RECT 71.600 264.395 74.460 264.775 ;
        RECT 104.050 264.395 106.910 264.775 ;
        RECT 0.240 263.995 0.620 264.375 ;
        RECT 4.160 263.995 4.540 264.375 ;
        RECT 35.140 264.165 35.520 264.215 ;
        RECT 37.560 264.165 37.940 264.215 ;
        RECT 35.140 263.885 37.940 264.165 ;
        RECT 35.140 263.835 35.520 263.885 ;
        RECT 37.560 263.835 37.940 263.885 ;
        RECT 67.590 264.165 67.970 264.215 ;
        RECT 70.010 264.165 70.390 264.215 ;
        RECT 67.590 263.885 70.390 264.165 ;
        RECT 67.590 263.835 67.970 263.885 ;
        RECT 70.010 263.835 70.390 263.885 ;
        RECT 100.040 264.165 100.420 264.215 ;
        RECT 102.460 264.165 102.840 264.215 ;
        RECT 100.040 263.885 102.840 264.165 ;
        RECT 100.040 263.835 100.420 263.885 ;
        RECT 102.460 263.835 102.840 263.885 ;
        RECT 132.490 264.165 132.870 264.215 ;
        RECT 134.910 264.165 135.290 264.215 ;
        RECT 132.490 263.885 135.290 264.165 ;
        RECT 132.490 263.835 132.870 263.885 ;
        RECT 134.910 263.835 135.290 263.885 ;
        RECT 6.700 262.555 9.560 262.935 ;
        RECT 39.150 262.555 42.010 262.935 ;
        RECT 71.600 262.555 74.460 262.935 ;
        RECT 104.050 262.555 106.910 262.935 ;
        RECT 137.355 262.495 137.735 262.875 ;
        RECT 139.395 262.495 139.775 262.875 ;
        RECT 141.180 262.495 141.560 262.875 ;
        RECT 36.420 262.325 36.800 262.375 ;
        RECT 37.560 262.325 37.940 262.375 ;
        RECT 36.420 262.045 37.940 262.325 ;
        RECT 36.420 261.995 36.800 262.045 ;
        RECT 37.560 261.995 37.940 262.045 ;
        RECT 68.870 262.325 69.250 262.375 ;
        RECT 70.010 262.325 70.390 262.375 ;
        RECT 68.870 262.045 70.390 262.325 ;
        RECT 68.870 261.995 69.250 262.045 ;
        RECT 70.010 261.995 70.390 262.045 ;
        RECT 101.320 262.325 101.700 262.375 ;
        RECT 102.460 262.325 102.840 262.375 ;
        RECT 101.320 262.045 102.840 262.325 ;
        RECT 101.320 261.995 101.700 262.045 ;
        RECT 102.460 261.995 102.840 262.045 ;
        RECT 133.770 262.325 134.150 262.375 ;
        RECT 134.910 262.325 135.290 262.375 ;
        RECT 133.770 262.045 135.290 262.325 ;
        RECT 133.770 261.995 134.150 262.045 ;
        RECT 134.910 261.995 135.290 262.045 ;
        RECT 0.240 260.995 0.620 261.375 ;
        RECT 4.160 260.995 4.540 261.375 ;
        RECT 6.700 260.715 9.560 261.095 ;
        RECT 39.150 260.715 42.010 261.095 ;
        RECT 71.600 260.715 74.460 261.095 ;
        RECT 104.050 260.715 106.910 261.095 ;
        RECT 37.560 260.155 38.080 260.535 ;
        RECT 70.010 260.155 70.530 260.535 ;
        RECT 102.460 260.155 102.980 260.535 ;
        RECT 134.910 260.155 135.430 260.535 ;
        RECT 137.355 259.495 137.735 259.875 ;
        RECT 139.395 259.495 139.775 259.875 ;
        RECT 141.180 259.495 141.560 259.875 ;
        RECT 0.240 257.995 0.620 258.375 ;
        RECT 4.160 257.995 4.540 258.375 ;
        RECT 0.240 254.995 0.620 255.375 ;
        RECT 137.355 253.495 137.735 253.875 ;
        RECT 139.395 253.495 139.775 253.875 ;
        RECT 141.180 253.495 141.560 253.875 ;
        RECT 0.240 251.995 0.620 252.375 ;
        RECT 4.160 251.995 4.540 252.375 ;
        RECT 37.060 251.590 37.940 251.970 ;
        RECT 69.510 251.590 70.390 251.970 ;
        RECT 101.960 251.590 102.840 251.970 ;
        RECT 134.410 251.590 135.290 251.970 ;
        RECT 6.700 251.030 9.560 251.410 ;
        RECT 39.150 251.030 42.010 251.410 ;
        RECT 71.600 251.030 74.460 251.410 ;
        RECT 104.050 251.030 106.910 251.410 ;
        RECT 137.355 250.495 137.735 250.875 ;
        RECT 139.395 250.495 139.775 250.875 ;
        RECT 141.180 250.495 141.560 250.875 ;
        RECT 35.780 250.080 36.160 250.130 ;
        RECT 37.560 250.080 37.940 250.130 ;
        RECT 35.780 249.800 37.940 250.080 ;
        RECT 35.780 249.750 36.160 249.800 ;
        RECT 37.560 249.750 37.940 249.800 ;
        RECT 68.230 250.080 68.610 250.130 ;
        RECT 70.010 250.080 70.390 250.130 ;
        RECT 68.230 249.800 70.390 250.080 ;
        RECT 68.230 249.750 68.610 249.800 ;
        RECT 70.010 249.750 70.390 249.800 ;
        RECT 100.680 250.080 101.060 250.130 ;
        RECT 102.460 250.080 102.840 250.130 ;
        RECT 100.680 249.800 102.840 250.080 ;
        RECT 100.680 249.750 101.060 249.800 ;
        RECT 102.460 249.750 102.840 249.800 ;
        RECT 133.130 250.080 133.510 250.130 ;
        RECT 134.910 250.080 135.290 250.130 ;
        RECT 133.130 249.800 135.290 250.080 ;
        RECT 133.130 249.750 133.510 249.800 ;
        RECT 134.910 249.750 135.290 249.800 ;
        RECT 0.240 248.995 0.620 249.375 ;
        RECT 4.160 248.995 4.540 249.375 ;
        RECT 6.700 249.190 9.560 249.570 ;
        RECT 39.150 249.190 42.010 249.570 ;
        RECT 71.600 249.190 74.460 249.570 ;
        RECT 104.050 249.190 106.910 249.570 ;
        RECT 34.500 248.235 34.880 248.285 ;
        RECT 37.560 248.235 37.940 248.285 ;
        RECT 34.500 247.955 37.940 248.235 ;
        RECT 34.500 247.905 34.880 247.955 ;
        RECT 37.560 247.905 37.940 247.955 ;
        RECT 66.950 248.235 67.330 248.285 ;
        RECT 70.010 248.235 70.390 248.285 ;
        RECT 66.950 247.955 70.390 248.235 ;
        RECT 66.950 247.905 67.330 247.955 ;
        RECT 70.010 247.905 70.390 247.955 ;
        RECT 99.400 248.235 99.780 248.285 ;
        RECT 102.460 248.235 102.840 248.285 ;
        RECT 99.400 247.955 102.840 248.235 ;
        RECT 99.400 247.905 99.780 247.955 ;
        RECT 102.460 247.905 102.840 247.955 ;
        RECT 131.850 248.235 132.230 248.285 ;
        RECT 134.910 248.235 135.290 248.285 ;
        RECT 131.850 247.955 135.290 248.235 ;
        RECT 131.850 247.905 132.230 247.955 ;
        RECT 134.910 247.905 135.290 247.955 ;
        RECT 6.700 247.345 9.560 247.725 ;
        RECT 39.150 247.345 42.010 247.725 ;
        RECT 71.600 247.345 74.460 247.725 ;
        RECT 104.050 247.345 106.910 247.725 ;
        RECT 137.355 247.495 137.735 247.875 ;
        RECT 139.395 247.495 139.775 247.875 ;
        RECT 141.180 247.495 141.560 247.875 ;
        RECT 6.700 246.585 9.560 246.965 ;
        RECT 39.150 246.585 42.010 246.965 ;
        RECT 71.600 246.585 74.460 246.965 ;
        RECT 104.050 246.585 106.910 246.965 ;
        RECT 0.240 245.995 0.620 246.375 ;
        RECT 4.160 245.995 4.540 246.375 ;
        RECT 33.220 245.595 33.600 245.645 ;
        RECT 37.560 245.595 37.940 245.645 ;
        RECT 33.220 245.315 37.940 245.595 ;
        RECT 33.220 245.265 33.600 245.315 ;
        RECT 37.560 245.265 37.940 245.315 ;
        RECT 65.670 245.595 66.050 245.645 ;
        RECT 70.010 245.595 70.390 245.645 ;
        RECT 65.670 245.315 70.390 245.595 ;
        RECT 65.670 245.265 66.050 245.315 ;
        RECT 70.010 245.265 70.390 245.315 ;
        RECT 98.120 245.595 98.500 245.645 ;
        RECT 102.460 245.595 102.840 245.645 ;
        RECT 98.120 245.315 102.840 245.595 ;
        RECT 98.120 245.265 98.500 245.315 ;
        RECT 102.460 245.265 102.840 245.315 ;
        RECT 130.570 245.595 130.950 245.645 ;
        RECT 134.910 245.595 135.290 245.645 ;
        RECT 130.570 245.315 135.290 245.595 ;
        RECT 130.570 245.265 130.950 245.315 ;
        RECT 134.910 245.265 135.290 245.315 ;
        RECT 6.700 244.705 9.560 245.085 ;
        RECT 39.150 244.705 42.010 245.085 ;
        RECT 71.600 244.705 74.460 245.085 ;
        RECT 104.050 244.705 106.910 245.085 ;
        RECT 137.355 244.495 137.735 244.875 ;
        RECT 139.395 244.495 139.775 244.875 ;
        RECT 141.180 244.495 141.560 244.875 ;
        RECT 31.940 243.755 32.320 243.805 ;
        RECT 37.560 243.755 37.940 243.805 ;
        RECT 31.940 243.475 37.940 243.755 ;
        RECT 31.940 243.425 32.320 243.475 ;
        RECT 37.560 243.425 37.940 243.475 ;
        RECT 64.390 243.755 64.770 243.805 ;
        RECT 70.010 243.755 70.390 243.805 ;
        RECT 64.390 243.475 70.390 243.755 ;
        RECT 64.390 243.425 64.770 243.475 ;
        RECT 70.010 243.425 70.390 243.475 ;
        RECT 96.840 243.755 97.220 243.805 ;
        RECT 102.460 243.755 102.840 243.805 ;
        RECT 96.840 243.475 102.840 243.755 ;
        RECT 96.840 243.425 97.220 243.475 ;
        RECT 102.460 243.425 102.840 243.475 ;
        RECT 129.290 243.755 129.670 243.805 ;
        RECT 134.910 243.755 135.290 243.805 ;
        RECT 129.290 243.475 135.290 243.755 ;
        RECT 129.290 243.425 129.670 243.475 ;
        RECT 134.910 243.425 135.290 243.475 ;
        RECT 0.240 242.995 0.620 243.375 ;
        RECT 4.160 242.995 4.540 243.375 ;
        RECT 6.700 242.865 9.560 243.245 ;
        RECT 39.150 242.865 42.010 243.245 ;
        RECT 71.600 242.865 74.460 243.245 ;
        RECT 104.050 242.865 106.910 243.245 ;
        RECT 30.660 241.910 31.040 241.960 ;
        RECT 37.560 241.910 37.940 241.960 ;
        RECT 30.660 241.630 37.940 241.910 ;
        RECT 30.660 241.580 31.040 241.630 ;
        RECT 37.560 241.580 37.940 241.630 ;
        RECT 63.110 241.910 63.490 241.960 ;
        RECT 70.010 241.910 70.390 241.960 ;
        RECT 63.110 241.630 70.390 241.910 ;
        RECT 63.110 241.580 63.490 241.630 ;
        RECT 70.010 241.580 70.390 241.630 ;
        RECT 95.560 241.910 95.940 241.960 ;
        RECT 102.460 241.910 102.840 241.960 ;
        RECT 95.560 241.630 102.840 241.910 ;
        RECT 95.560 241.580 95.940 241.630 ;
        RECT 102.460 241.580 102.840 241.630 ;
        RECT 128.010 241.910 128.390 241.960 ;
        RECT 134.910 241.910 135.290 241.960 ;
        RECT 128.010 241.630 135.290 241.910 ;
        RECT 128.010 241.580 128.390 241.630 ;
        RECT 134.910 241.580 135.290 241.630 ;
        RECT 137.355 241.495 137.735 241.875 ;
        RECT 139.395 241.495 139.775 241.875 ;
        RECT 141.180 241.495 141.560 241.875 ;
        RECT 6.700 241.020 9.560 241.400 ;
        RECT 39.150 241.020 42.010 241.400 ;
        RECT 71.600 241.020 74.460 241.400 ;
        RECT 104.050 241.020 106.910 241.400 ;
        RECT 0.240 239.995 0.620 240.375 ;
        RECT 4.160 239.995 4.540 240.375 ;
        RECT 6.700 240.260 9.560 240.640 ;
        RECT 39.150 240.260 42.010 240.640 ;
        RECT 71.600 240.260 74.460 240.640 ;
        RECT 104.050 240.260 106.910 240.640 ;
        RECT 29.380 239.270 29.760 239.320 ;
        RECT 37.560 239.270 37.940 239.320 ;
        RECT 29.380 238.990 37.940 239.270 ;
        RECT 29.380 238.940 29.760 238.990 ;
        RECT 37.560 238.940 37.940 238.990 ;
        RECT 61.830 239.270 62.210 239.320 ;
        RECT 70.010 239.270 70.390 239.320 ;
        RECT 61.830 238.990 70.390 239.270 ;
        RECT 61.830 238.940 62.210 238.990 ;
        RECT 70.010 238.940 70.390 238.990 ;
        RECT 94.280 239.270 94.660 239.320 ;
        RECT 102.460 239.270 102.840 239.320 ;
        RECT 94.280 238.990 102.840 239.270 ;
        RECT 94.280 238.940 94.660 238.990 ;
        RECT 102.460 238.940 102.840 238.990 ;
        RECT 126.730 239.270 127.110 239.320 ;
        RECT 134.910 239.270 135.290 239.320 ;
        RECT 126.730 238.990 135.290 239.270 ;
        RECT 126.730 238.940 127.110 238.990 ;
        RECT 134.910 238.940 135.290 238.990 ;
        RECT 6.700 238.380 9.560 238.760 ;
        RECT 39.150 238.380 42.010 238.760 ;
        RECT 71.600 238.380 74.460 238.760 ;
        RECT 104.050 238.380 106.910 238.760 ;
        RECT 137.355 238.495 137.735 238.875 ;
        RECT 139.395 238.495 139.775 238.875 ;
        RECT 141.180 238.495 141.560 238.875 ;
        RECT 28.100 237.430 28.480 237.480 ;
        RECT 37.560 237.430 37.940 237.480 ;
        RECT 0.240 236.995 0.620 237.375 ;
        RECT 4.160 236.995 4.540 237.375 ;
        RECT 28.100 237.150 37.940 237.430 ;
        RECT 28.100 237.100 28.480 237.150 ;
        RECT 37.560 237.100 37.940 237.150 ;
        RECT 60.550 237.430 60.930 237.480 ;
        RECT 70.010 237.430 70.390 237.480 ;
        RECT 60.550 237.150 70.390 237.430 ;
        RECT 60.550 237.100 60.930 237.150 ;
        RECT 70.010 237.100 70.390 237.150 ;
        RECT 93.000 237.430 93.380 237.480 ;
        RECT 102.460 237.430 102.840 237.480 ;
        RECT 93.000 237.150 102.840 237.430 ;
        RECT 93.000 237.100 93.380 237.150 ;
        RECT 102.460 237.100 102.840 237.150 ;
        RECT 125.450 237.430 125.830 237.480 ;
        RECT 134.910 237.430 135.290 237.480 ;
        RECT 125.450 237.150 135.290 237.430 ;
        RECT 125.450 237.100 125.830 237.150 ;
        RECT 134.910 237.100 135.290 237.150 ;
        RECT 6.700 236.540 9.560 236.920 ;
        RECT 39.150 236.540 42.010 236.920 ;
        RECT 71.600 236.540 74.460 236.920 ;
        RECT 104.050 236.540 106.910 236.920 ;
        RECT 6.700 235.820 9.560 236.200 ;
        RECT 39.150 235.820 42.010 236.200 ;
        RECT 71.600 235.820 74.460 236.200 ;
        RECT 104.050 235.820 106.910 236.200 ;
        RECT 28.740 235.590 29.120 235.640 ;
        RECT 37.560 235.590 37.940 235.640 ;
        RECT 28.740 235.310 37.940 235.590 ;
        RECT 28.740 235.260 29.120 235.310 ;
        RECT 37.560 235.260 37.940 235.310 ;
        RECT 61.190 235.590 61.570 235.640 ;
        RECT 70.010 235.590 70.390 235.640 ;
        RECT 61.190 235.310 70.390 235.590 ;
        RECT 61.190 235.260 61.570 235.310 ;
        RECT 70.010 235.260 70.390 235.310 ;
        RECT 93.640 235.590 94.020 235.640 ;
        RECT 102.460 235.590 102.840 235.640 ;
        RECT 93.640 235.310 102.840 235.590 ;
        RECT 93.640 235.260 94.020 235.310 ;
        RECT 102.460 235.260 102.840 235.310 ;
        RECT 126.090 235.590 126.470 235.640 ;
        RECT 134.910 235.590 135.290 235.640 ;
        RECT 126.090 235.310 135.290 235.590 ;
        RECT 126.090 235.260 126.470 235.310 ;
        RECT 134.910 235.260 135.290 235.310 ;
        RECT 0.240 233.610 0.620 233.990 ;
        RECT 4.160 233.610 4.540 233.990 ;
        RECT 6.700 233.980 9.560 234.360 ;
        RECT 39.150 233.980 42.010 234.360 ;
        RECT 71.600 233.980 74.460 234.360 ;
        RECT 104.050 233.980 106.910 234.360 ;
        RECT 30.020 233.750 30.400 233.800 ;
        RECT 37.560 233.750 37.940 233.800 ;
        RECT 30.020 233.470 37.940 233.750 ;
        RECT 30.020 233.420 30.400 233.470 ;
        RECT 37.560 233.420 37.940 233.470 ;
        RECT 62.470 233.750 62.850 233.800 ;
        RECT 70.010 233.750 70.390 233.800 ;
        RECT 62.470 233.470 70.390 233.750 ;
        RECT 62.470 233.420 62.850 233.470 ;
        RECT 70.010 233.420 70.390 233.470 ;
        RECT 94.920 233.750 95.300 233.800 ;
        RECT 102.460 233.750 102.840 233.800 ;
        RECT 94.920 233.470 102.840 233.750 ;
        RECT 94.920 233.420 95.300 233.470 ;
        RECT 102.460 233.420 102.840 233.470 ;
        RECT 127.370 233.750 127.750 233.800 ;
        RECT 134.910 233.750 135.290 233.800 ;
        RECT 127.370 233.470 135.290 233.750 ;
        RECT 127.370 233.420 127.750 233.470 ;
        RECT 134.910 233.420 135.290 233.470 ;
        RECT 6.700 232.095 9.560 232.475 ;
        RECT 39.150 232.095 42.010 232.475 ;
        RECT 71.600 232.095 74.460 232.475 ;
        RECT 104.050 232.095 106.910 232.475 ;
        RECT 137.355 232.110 137.735 232.490 ;
        RECT 139.395 232.110 139.775 232.490 ;
        RECT 141.180 232.110 141.560 232.490 ;
        RECT 6.700 231.335 9.560 231.715 ;
        RECT 39.150 231.335 42.010 231.715 ;
        RECT 71.600 231.335 74.460 231.715 ;
        RECT 104.050 231.335 106.910 231.715 ;
        RECT 31.300 231.105 31.680 231.155 ;
        RECT 37.560 231.105 37.940 231.155 ;
        RECT 0.240 230.610 0.620 230.990 ;
        RECT 4.160 230.610 4.540 230.990 ;
        RECT 31.300 230.825 37.940 231.105 ;
        RECT 31.300 230.775 31.680 230.825 ;
        RECT 37.560 230.775 37.940 230.825 ;
        RECT 63.750 231.105 64.130 231.155 ;
        RECT 70.010 231.105 70.390 231.155 ;
        RECT 63.750 230.825 70.390 231.105 ;
        RECT 63.750 230.775 64.130 230.825 ;
        RECT 70.010 230.775 70.390 230.825 ;
        RECT 96.200 231.105 96.580 231.155 ;
        RECT 102.460 231.105 102.840 231.155 ;
        RECT 96.200 230.825 102.840 231.105 ;
        RECT 96.200 230.775 96.580 230.825 ;
        RECT 102.460 230.775 102.840 230.825 ;
        RECT 128.650 231.105 129.030 231.155 ;
        RECT 134.910 231.105 135.290 231.155 ;
        RECT 128.650 230.825 135.290 231.105 ;
        RECT 128.650 230.775 129.030 230.825 ;
        RECT 134.910 230.775 135.290 230.825 ;
        RECT 6.700 229.495 9.560 229.875 ;
        RECT 39.150 229.495 42.010 229.875 ;
        RECT 71.600 229.495 74.460 229.875 ;
        RECT 104.050 229.495 106.910 229.875 ;
        RECT 32.580 229.265 32.960 229.315 ;
        RECT 37.560 229.265 37.940 229.315 ;
        RECT 32.580 228.985 37.940 229.265 ;
        RECT 32.580 228.935 32.960 228.985 ;
        RECT 37.560 228.935 37.940 228.985 ;
        RECT 65.030 229.265 65.410 229.315 ;
        RECT 70.010 229.265 70.390 229.315 ;
        RECT 65.030 228.985 70.390 229.265 ;
        RECT 65.030 228.935 65.410 228.985 ;
        RECT 70.010 228.935 70.390 228.985 ;
        RECT 97.480 229.265 97.860 229.315 ;
        RECT 102.460 229.265 102.840 229.315 ;
        RECT 97.480 228.985 102.840 229.265 ;
        RECT 97.480 228.935 97.860 228.985 ;
        RECT 102.460 228.935 102.840 228.985 ;
        RECT 129.930 229.265 130.310 229.315 ;
        RECT 134.910 229.265 135.290 229.315 ;
        RECT 129.930 228.985 135.290 229.265 ;
        RECT 137.355 229.110 137.735 229.490 ;
        RECT 139.395 229.110 139.775 229.490 ;
        RECT 141.180 229.110 141.560 229.490 ;
        RECT 129.930 228.935 130.310 228.985 ;
        RECT 134.910 228.935 135.290 228.985 ;
        RECT 0.240 227.610 0.620 227.990 ;
        RECT 4.160 227.610 4.540 227.990 ;
        RECT 6.700 227.655 9.560 228.035 ;
        RECT 39.150 227.655 42.010 228.035 ;
        RECT 71.600 227.655 74.460 228.035 ;
        RECT 104.050 227.655 106.910 228.035 ;
        RECT 33.860 227.425 34.240 227.475 ;
        RECT 37.560 227.425 37.940 227.475 ;
        RECT 33.860 227.145 37.940 227.425 ;
        RECT 33.860 227.095 34.240 227.145 ;
        RECT 37.560 227.095 37.940 227.145 ;
        RECT 66.310 227.425 66.690 227.475 ;
        RECT 70.010 227.425 70.390 227.475 ;
        RECT 66.310 227.145 70.390 227.425 ;
        RECT 66.310 227.095 66.690 227.145 ;
        RECT 70.010 227.095 70.390 227.145 ;
        RECT 98.760 227.425 99.140 227.475 ;
        RECT 102.460 227.425 102.840 227.475 ;
        RECT 98.760 227.145 102.840 227.425 ;
        RECT 98.760 227.095 99.140 227.145 ;
        RECT 102.460 227.095 102.840 227.145 ;
        RECT 131.210 227.425 131.590 227.475 ;
        RECT 134.910 227.425 135.290 227.475 ;
        RECT 131.210 227.145 135.290 227.425 ;
        RECT 131.210 227.095 131.590 227.145 ;
        RECT 134.910 227.095 135.290 227.145 ;
        RECT 6.700 225.770 9.560 226.150 ;
        RECT 39.150 225.770 42.010 226.150 ;
        RECT 71.600 225.770 74.460 226.150 ;
        RECT 104.050 225.770 106.910 226.150 ;
        RECT 137.355 226.110 137.735 226.490 ;
        RECT 139.395 226.110 139.775 226.490 ;
        RECT 141.180 226.110 141.560 226.490 ;
        RECT 6.700 225.010 9.560 225.390 ;
        RECT 39.150 225.010 42.010 225.390 ;
        RECT 71.600 225.010 74.460 225.390 ;
        RECT 104.050 225.010 106.910 225.390 ;
        RECT 0.240 224.610 0.620 224.990 ;
        RECT 4.160 224.610 4.540 224.990 ;
        RECT 35.140 224.780 35.520 224.830 ;
        RECT 37.560 224.780 37.940 224.830 ;
        RECT 35.140 224.500 37.940 224.780 ;
        RECT 35.140 224.450 35.520 224.500 ;
        RECT 37.560 224.450 37.940 224.500 ;
        RECT 67.590 224.780 67.970 224.830 ;
        RECT 70.010 224.780 70.390 224.830 ;
        RECT 67.590 224.500 70.390 224.780 ;
        RECT 67.590 224.450 67.970 224.500 ;
        RECT 70.010 224.450 70.390 224.500 ;
        RECT 100.040 224.780 100.420 224.830 ;
        RECT 102.460 224.780 102.840 224.830 ;
        RECT 100.040 224.500 102.840 224.780 ;
        RECT 100.040 224.450 100.420 224.500 ;
        RECT 102.460 224.450 102.840 224.500 ;
        RECT 132.490 224.780 132.870 224.830 ;
        RECT 134.910 224.780 135.290 224.830 ;
        RECT 132.490 224.500 135.290 224.780 ;
        RECT 132.490 224.450 132.870 224.500 ;
        RECT 134.910 224.450 135.290 224.500 ;
        RECT 6.700 223.170 9.560 223.550 ;
        RECT 39.150 223.170 42.010 223.550 ;
        RECT 71.600 223.170 74.460 223.550 ;
        RECT 104.050 223.170 106.910 223.550 ;
        RECT 137.355 223.110 137.735 223.490 ;
        RECT 139.395 223.110 139.775 223.490 ;
        RECT 141.180 223.110 141.560 223.490 ;
        RECT 36.420 222.940 36.800 222.990 ;
        RECT 37.560 222.940 37.940 222.990 ;
        RECT 36.420 222.660 37.940 222.940 ;
        RECT 36.420 222.610 36.800 222.660 ;
        RECT 37.560 222.610 37.940 222.660 ;
        RECT 68.870 222.940 69.250 222.990 ;
        RECT 70.010 222.940 70.390 222.990 ;
        RECT 68.870 222.660 70.390 222.940 ;
        RECT 68.870 222.610 69.250 222.660 ;
        RECT 70.010 222.610 70.390 222.660 ;
        RECT 101.320 222.940 101.700 222.990 ;
        RECT 102.460 222.940 102.840 222.990 ;
        RECT 101.320 222.660 102.840 222.940 ;
        RECT 101.320 222.610 101.700 222.660 ;
        RECT 102.460 222.610 102.840 222.660 ;
        RECT 133.770 222.940 134.150 222.990 ;
        RECT 134.910 222.940 135.290 222.990 ;
        RECT 133.770 222.660 135.290 222.940 ;
        RECT 133.770 222.610 134.150 222.660 ;
        RECT 134.910 222.610 135.290 222.660 ;
        RECT 0.240 221.610 0.620 221.990 ;
        RECT 4.160 221.610 4.540 221.990 ;
        RECT 6.700 221.330 9.560 221.710 ;
        RECT 39.150 221.330 42.010 221.710 ;
        RECT 71.600 221.330 74.460 221.710 ;
        RECT 104.050 221.330 106.910 221.710 ;
        RECT 37.560 220.770 38.080 221.150 ;
        RECT 70.010 220.770 70.530 221.150 ;
        RECT 102.460 220.770 102.980 221.150 ;
        RECT 134.910 220.770 135.430 221.150 ;
        RECT 137.355 220.110 137.735 220.490 ;
        RECT 139.395 220.110 139.775 220.490 ;
        RECT 141.180 220.110 141.560 220.490 ;
        RECT 0.240 218.610 0.620 218.990 ;
        RECT 4.160 218.610 4.540 218.990 ;
        RECT 0.240 215.610 0.620 215.990 ;
        RECT 137.355 214.110 137.735 214.490 ;
        RECT 139.395 214.110 139.775 214.490 ;
        RECT 141.180 214.110 141.560 214.490 ;
        RECT 0.240 212.610 0.620 212.990 ;
        RECT 4.160 212.610 4.540 212.990 ;
        RECT 37.060 212.205 37.940 212.585 ;
        RECT 69.510 212.205 70.390 212.585 ;
        RECT 101.960 212.205 102.840 212.585 ;
        RECT 134.410 212.205 135.290 212.585 ;
        RECT 6.700 211.645 9.560 212.025 ;
        RECT 39.150 211.645 42.010 212.025 ;
        RECT 71.600 211.645 74.460 212.025 ;
        RECT 104.050 211.645 106.910 212.025 ;
        RECT 137.355 211.110 137.735 211.490 ;
        RECT 139.395 211.110 139.775 211.490 ;
        RECT 141.180 211.110 141.560 211.490 ;
        RECT 35.780 210.695 36.160 210.745 ;
        RECT 37.560 210.695 37.940 210.745 ;
        RECT 35.780 210.415 37.940 210.695 ;
        RECT 35.780 210.365 36.160 210.415 ;
        RECT 37.560 210.365 37.940 210.415 ;
        RECT 68.230 210.695 68.610 210.745 ;
        RECT 70.010 210.695 70.390 210.745 ;
        RECT 68.230 210.415 70.390 210.695 ;
        RECT 68.230 210.365 68.610 210.415 ;
        RECT 70.010 210.365 70.390 210.415 ;
        RECT 100.680 210.695 101.060 210.745 ;
        RECT 102.460 210.695 102.840 210.745 ;
        RECT 100.680 210.415 102.840 210.695 ;
        RECT 100.680 210.365 101.060 210.415 ;
        RECT 102.460 210.365 102.840 210.415 ;
        RECT 133.130 210.695 133.510 210.745 ;
        RECT 134.910 210.695 135.290 210.745 ;
        RECT 133.130 210.415 135.290 210.695 ;
        RECT 133.130 210.365 133.510 210.415 ;
        RECT 134.910 210.365 135.290 210.415 ;
        RECT 0.240 209.610 0.620 209.990 ;
        RECT 4.160 209.610 4.540 209.990 ;
        RECT 6.700 209.805 9.560 210.185 ;
        RECT 39.150 209.805 42.010 210.185 ;
        RECT 71.600 209.805 74.460 210.185 ;
        RECT 104.050 209.805 106.910 210.185 ;
        RECT 34.500 208.850 34.880 208.900 ;
        RECT 37.560 208.850 37.940 208.900 ;
        RECT 34.500 208.570 37.940 208.850 ;
        RECT 34.500 208.520 34.880 208.570 ;
        RECT 37.560 208.520 37.940 208.570 ;
        RECT 66.950 208.850 67.330 208.900 ;
        RECT 70.010 208.850 70.390 208.900 ;
        RECT 66.950 208.570 70.390 208.850 ;
        RECT 66.950 208.520 67.330 208.570 ;
        RECT 70.010 208.520 70.390 208.570 ;
        RECT 99.400 208.850 99.780 208.900 ;
        RECT 102.460 208.850 102.840 208.900 ;
        RECT 99.400 208.570 102.840 208.850 ;
        RECT 99.400 208.520 99.780 208.570 ;
        RECT 102.460 208.520 102.840 208.570 ;
        RECT 131.850 208.850 132.230 208.900 ;
        RECT 134.910 208.850 135.290 208.900 ;
        RECT 131.850 208.570 135.290 208.850 ;
        RECT 131.850 208.520 132.230 208.570 ;
        RECT 134.910 208.520 135.290 208.570 ;
        RECT 6.700 207.960 9.560 208.340 ;
        RECT 39.150 207.960 42.010 208.340 ;
        RECT 71.600 207.960 74.460 208.340 ;
        RECT 104.050 207.960 106.910 208.340 ;
        RECT 137.355 208.110 137.735 208.490 ;
        RECT 139.395 208.110 139.775 208.490 ;
        RECT 141.180 208.110 141.560 208.490 ;
        RECT 6.700 207.200 9.560 207.580 ;
        RECT 39.150 207.200 42.010 207.580 ;
        RECT 71.600 207.200 74.460 207.580 ;
        RECT 104.050 207.200 106.910 207.580 ;
        RECT 0.240 206.610 0.620 206.990 ;
        RECT 4.160 206.610 4.540 206.990 ;
        RECT 33.220 206.210 33.600 206.260 ;
        RECT 37.560 206.210 37.940 206.260 ;
        RECT 33.220 205.930 37.940 206.210 ;
        RECT 33.220 205.880 33.600 205.930 ;
        RECT 37.560 205.880 37.940 205.930 ;
        RECT 65.670 206.210 66.050 206.260 ;
        RECT 70.010 206.210 70.390 206.260 ;
        RECT 65.670 205.930 70.390 206.210 ;
        RECT 65.670 205.880 66.050 205.930 ;
        RECT 70.010 205.880 70.390 205.930 ;
        RECT 98.120 206.210 98.500 206.260 ;
        RECT 102.460 206.210 102.840 206.260 ;
        RECT 98.120 205.930 102.840 206.210 ;
        RECT 98.120 205.880 98.500 205.930 ;
        RECT 102.460 205.880 102.840 205.930 ;
        RECT 130.570 206.210 130.950 206.260 ;
        RECT 134.910 206.210 135.290 206.260 ;
        RECT 130.570 205.930 135.290 206.210 ;
        RECT 130.570 205.880 130.950 205.930 ;
        RECT 134.910 205.880 135.290 205.930 ;
        RECT 6.700 205.320 9.560 205.700 ;
        RECT 39.150 205.320 42.010 205.700 ;
        RECT 71.600 205.320 74.460 205.700 ;
        RECT 104.050 205.320 106.910 205.700 ;
        RECT 137.355 205.110 137.735 205.490 ;
        RECT 139.395 205.110 139.775 205.490 ;
        RECT 141.180 205.110 141.560 205.490 ;
        RECT 31.940 204.370 32.320 204.420 ;
        RECT 37.560 204.370 37.940 204.420 ;
        RECT 31.940 204.090 37.940 204.370 ;
        RECT 31.940 204.040 32.320 204.090 ;
        RECT 37.560 204.040 37.940 204.090 ;
        RECT 64.390 204.370 64.770 204.420 ;
        RECT 70.010 204.370 70.390 204.420 ;
        RECT 64.390 204.090 70.390 204.370 ;
        RECT 64.390 204.040 64.770 204.090 ;
        RECT 70.010 204.040 70.390 204.090 ;
        RECT 96.840 204.370 97.220 204.420 ;
        RECT 102.460 204.370 102.840 204.420 ;
        RECT 96.840 204.090 102.840 204.370 ;
        RECT 96.840 204.040 97.220 204.090 ;
        RECT 102.460 204.040 102.840 204.090 ;
        RECT 129.290 204.370 129.670 204.420 ;
        RECT 134.910 204.370 135.290 204.420 ;
        RECT 129.290 204.090 135.290 204.370 ;
        RECT 129.290 204.040 129.670 204.090 ;
        RECT 134.910 204.040 135.290 204.090 ;
        RECT 0.240 203.610 0.620 203.990 ;
        RECT 4.160 203.610 4.540 203.990 ;
        RECT 6.700 203.480 9.560 203.860 ;
        RECT 39.150 203.480 42.010 203.860 ;
        RECT 71.600 203.480 74.460 203.860 ;
        RECT 104.050 203.480 106.910 203.860 ;
        RECT 30.660 202.525 31.040 202.575 ;
        RECT 37.560 202.525 37.940 202.575 ;
        RECT 30.660 202.245 37.940 202.525 ;
        RECT 30.660 202.195 31.040 202.245 ;
        RECT 37.560 202.195 37.940 202.245 ;
        RECT 63.110 202.525 63.490 202.575 ;
        RECT 70.010 202.525 70.390 202.575 ;
        RECT 63.110 202.245 70.390 202.525 ;
        RECT 63.110 202.195 63.490 202.245 ;
        RECT 70.010 202.195 70.390 202.245 ;
        RECT 95.560 202.525 95.940 202.575 ;
        RECT 102.460 202.525 102.840 202.575 ;
        RECT 95.560 202.245 102.840 202.525 ;
        RECT 95.560 202.195 95.940 202.245 ;
        RECT 102.460 202.195 102.840 202.245 ;
        RECT 128.010 202.525 128.390 202.575 ;
        RECT 134.910 202.525 135.290 202.575 ;
        RECT 128.010 202.245 135.290 202.525 ;
        RECT 128.010 202.195 128.390 202.245 ;
        RECT 134.910 202.195 135.290 202.245 ;
        RECT 137.355 202.110 137.735 202.490 ;
        RECT 139.395 202.110 139.775 202.490 ;
        RECT 141.180 202.110 141.560 202.490 ;
        RECT 6.700 201.635 9.560 202.015 ;
        RECT 39.150 201.635 42.010 202.015 ;
        RECT 71.600 201.635 74.460 202.015 ;
        RECT 104.050 201.635 106.910 202.015 ;
        RECT 0.240 200.610 0.620 200.990 ;
        RECT 4.160 200.610 4.540 200.990 ;
        RECT 6.700 200.875 9.560 201.255 ;
        RECT 39.150 200.875 42.010 201.255 ;
        RECT 71.600 200.875 74.460 201.255 ;
        RECT 104.050 200.875 106.910 201.255 ;
        RECT 29.380 199.885 29.760 199.935 ;
        RECT 37.560 199.885 37.940 199.935 ;
        RECT 29.380 199.605 37.940 199.885 ;
        RECT 29.380 199.555 29.760 199.605 ;
        RECT 37.560 199.555 37.940 199.605 ;
        RECT 61.830 199.885 62.210 199.935 ;
        RECT 70.010 199.885 70.390 199.935 ;
        RECT 61.830 199.605 70.390 199.885 ;
        RECT 61.830 199.555 62.210 199.605 ;
        RECT 70.010 199.555 70.390 199.605 ;
        RECT 94.280 199.885 94.660 199.935 ;
        RECT 102.460 199.885 102.840 199.935 ;
        RECT 94.280 199.605 102.840 199.885 ;
        RECT 94.280 199.555 94.660 199.605 ;
        RECT 102.460 199.555 102.840 199.605 ;
        RECT 126.730 199.885 127.110 199.935 ;
        RECT 134.910 199.885 135.290 199.935 ;
        RECT 126.730 199.605 135.290 199.885 ;
        RECT 126.730 199.555 127.110 199.605 ;
        RECT 134.910 199.555 135.290 199.605 ;
        RECT 6.700 198.995 9.560 199.375 ;
        RECT 39.150 198.995 42.010 199.375 ;
        RECT 71.600 198.995 74.460 199.375 ;
        RECT 104.050 198.995 106.910 199.375 ;
        RECT 137.355 199.110 137.735 199.490 ;
        RECT 139.395 199.110 139.775 199.490 ;
        RECT 141.180 199.110 141.560 199.490 ;
        RECT 28.100 198.045 28.480 198.095 ;
        RECT 37.560 198.045 37.940 198.095 ;
        RECT 0.240 197.610 0.620 197.990 ;
        RECT 4.160 197.610 4.540 197.990 ;
        RECT 28.100 197.765 37.940 198.045 ;
        RECT 28.100 197.715 28.480 197.765 ;
        RECT 37.560 197.715 37.940 197.765 ;
        RECT 60.550 198.045 60.930 198.095 ;
        RECT 70.010 198.045 70.390 198.095 ;
        RECT 60.550 197.765 70.390 198.045 ;
        RECT 60.550 197.715 60.930 197.765 ;
        RECT 70.010 197.715 70.390 197.765 ;
        RECT 93.000 198.045 93.380 198.095 ;
        RECT 102.460 198.045 102.840 198.095 ;
        RECT 93.000 197.765 102.840 198.045 ;
        RECT 93.000 197.715 93.380 197.765 ;
        RECT 102.460 197.715 102.840 197.765 ;
        RECT 125.450 198.045 125.830 198.095 ;
        RECT 134.910 198.045 135.290 198.095 ;
        RECT 125.450 197.765 135.290 198.045 ;
        RECT 125.450 197.715 125.830 197.765 ;
        RECT 134.910 197.715 135.290 197.765 ;
        RECT 6.700 197.155 9.560 197.535 ;
        RECT 39.150 197.155 42.010 197.535 ;
        RECT 71.600 197.155 74.460 197.535 ;
        RECT 104.050 197.155 106.910 197.535 ;
        RECT 6.700 196.435 9.560 196.815 ;
        RECT 39.150 196.435 42.010 196.815 ;
        RECT 71.600 196.435 74.460 196.815 ;
        RECT 104.050 196.435 106.910 196.815 ;
        RECT 28.740 196.205 29.120 196.255 ;
        RECT 37.560 196.205 37.940 196.255 ;
        RECT 28.740 195.925 37.940 196.205 ;
        RECT 28.740 195.875 29.120 195.925 ;
        RECT 37.560 195.875 37.940 195.925 ;
        RECT 61.190 196.205 61.570 196.255 ;
        RECT 70.010 196.205 70.390 196.255 ;
        RECT 61.190 195.925 70.390 196.205 ;
        RECT 61.190 195.875 61.570 195.925 ;
        RECT 70.010 195.875 70.390 195.925 ;
        RECT 93.640 196.205 94.020 196.255 ;
        RECT 102.460 196.205 102.840 196.255 ;
        RECT 93.640 195.925 102.840 196.205 ;
        RECT 93.640 195.875 94.020 195.925 ;
        RECT 102.460 195.875 102.840 195.925 ;
        RECT 126.090 196.205 126.470 196.255 ;
        RECT 134.910 196.205 135.290 196.255 ;
        RECT 126.090 195.925 135.290 196.205 ;
        RECT 126.090 195.875 126.470 195.925 ;
        RECT 134.910 195.875 135.290 195.925 ;
        RECT 0.240 194.225 0.620 194.605 ;
        RECT 4.160 194.225 4.540 194.605 ;
        RECT 6.700 194.595 9.560 194.975 ;
        RECT 39.150 194.595 42.010 194.975 ;
        RECT 71.600 194.595 74.460 194.975 ;
        RECT 104.050 194.595 106.910 194.975 ;
        RECT 30.020 194.365 30.400 194.415 ;
        RECT 37.560 194.365 37.940 194.415 ;
        RECT 30.020 194.085 37.940 194.365 ;
        RECT 30.020 194.035 30.400 194.085 ;
        RECT 37.560 194.035 37.940 194.085 ;
        RECT 62.470 194.365 62.850 194.415 ;
        RECT 70.010 194.365 70.390 194.415 ;
        RECT 62.470 194.085 70.390 194.365 ;
        RECT 62.470 194.035 62.850 194.085 ;
        RECT 70.010 194.035 70.390 194.085 ;
        RECT 94.920 194.365 95.300 194.415 ;
        RECT 102.460 194.365 102.840 194.415 ;
        RECT 94.920 194.085 102.840 194.365 ;
        RECT 94.920 194.035 95.300 194.085 ;
        RECT 102.460 194.035 102.840 194.085 ;
        RECT 127.370 194.365 127.750 194.415 ;
        RECT 134.910 194.365 135.290 194.415 ;
        RECT 127.370 194.085 135.290 194.365 ;
        RECT 127.370 194.035 127.750 194.085 ;
        RECT 134.910 194.035 135.290 194.085 ;
        RECT 6.700 192.710 9.560 193.090 ;
        RECT 39.150 192.710 42.010 193.090 ;
        RECT 71.600 192.710 74.460 193.090 ;
        RECT 104.050 192.710 106.910 193.090 ;
        RECT 137.355 192.725 137.735 193.105 ;
        RECT 139.395 192.725 139.775 193.105 ;
        RECT 141.180 192.725 141.560 193.105 ;
        RECT 6.700 191.950 9.560 192.330 ;
        RECT 39.150 191.950 42.010 192.330 ;
        RECT 71.600 191.950 74.460 192.330 ;
        RECT 104.050 191.950 106.910 192.330 ;
        RECT 31.300 191.720 31.680 191.770 ;
        RECT 37.560 191.720 37.940 191.770 ;
        RECT 0.240 191.225 0.620 191.605 ;
        RECT 4.160 191.225 4.540 191.605 ;
        RECT 31.300 191.440 37.940 191.720 ;
        RECT 31.300 191.390 31.680 191.440 ;
        RECT 37.560 191.390 37.940 191.440 ;
        RECT 63.750 191.720 64.130 191.770 ;
        RECT 70.010 191.720 70.390 191.770 ;
        RECT 63.750 191.440 70.390 191.720 ;
        RECT 63.750 191.390 64.130 191.440 ;
        RECT 70.010 191.390 70.390 191.440 ;
        RECT 96.200 191.720 96.580 191.770 ;
        RECT 102.460 191.720 102.840 191.770 ;
        RECT 96.200 191.440 102.840 191.720 ;
        RECT 96.200 191.390 96.580 191.440 ;
        RECT 102.460 191.390 102.840 191.440 ;
        RECT 128.650 191.720 129.030 191.770 ;
        RECT 134.910 191.720 135.290 191.770 ;
        RECT 128.650 191.440 135.290 191.720 ;
        RECT 128.650 191.390 129.030 191.440 ;
        RECT 134.910 191.390 135.290 191.440 ;
        RECT 6.700 190.110 9.560 190.490 ;
        RECT 39.150 190.110 42.010 190.490 ;
        RECT 71.600 190.110 74.460 190.490 ;
        RECT 104.050 190.110 106.910 190.490 ;
        RECT 32.580 189.880 32.960 189.930 ;
        RECT 37.560 189.880 37.940 189.930 ;
        RECT 32.580 189.600 37.940 189.880 ;
        RECT 32.580 189.550 32.960 189.600 ;
        RECT 37.560 189.550 37.940 189.600 ;
        RECT 65.030 189.880 65.410 189.930 ;
        RECT 70.010 189.880 70.390 189.930 ;
        RECT 65.030 189.600 70.390 189.880 ;
        RECT 65.030 189.550 65.410 189.600 ;
        RECT 70.010 189.550 70.390 189.600 ;
        RECT 97.480 189.880 97.860 189.930 ;
        RECT 102.460 189.880 102.840 189.930 ;
        RECT 97.480 189.600 102.840 189.880 ;
        RECT 97.480 189.550 97.860 189.600 ;
        RECT 102.460 189.550 102.840 189.600 ;
        RECT 129.930 189.880 130.310 189.930 ;
        RECT 134.910 189.880 135.290 189.930 ;
        RECT 129.930 189.600 135.290 189.880 ;
        RECT 137.355 189.725 137.735 190.105 ;
        RECT 139.395 189.725 139.775 190.105 ;
        RECT 141.180 189.725 141.560 190.105 ;
        RECT 129.930 189.550 130.310 189.600 ;
        RECT 134.910 189.550 135.290 189.600 ;
        RECT 0.240 188.225 0.620 188.605 ;
        RECT 4.160 188.225 4.540 188.605 ;
        RECT 6.700 188.270 9.560 188.650 ;
        RECT 39.150 188.270 42.010 188.650 ;
        RECT 71.600 188.270 74.460 188.650 ;
        RECT 104.050 188.270 106.910 188.650 ;
        RECT 33.860 188.040 34.240 188.090 ;
        RECT 37.560 188.040 37.940 188.090 ;
        RECT 33.860 187.760 37.940 188.040 ;
        RECT 33.860 187.710 34.240 187.760 ;
        RECT 37.560 187.710 37.940 187.760 ;
        RECT 66.310 188.040 66.690 188.090 ;
        RECT 70.010 188.040 70.390 188.090 ;
        RECT 66.310 187.760 70.390 188.040 ;
        RECT 66.310 187.710 66.690 187.760 ;
        RECT 70.010 187.710 70.390 187.760 ;
        RECT 98.760 188.040 99.140 188.090 ;
        RECT 102.460 188.040 102.840 188.090 ;
        RECT 98.760 187.760 102.840 188.040 ;
        RECT 98.760 187.710 99.140 187.760 ;
        RECT 102.460 187.710 102.840 187.760 ;
        RECT 131.210 188.040 131.590 188.090 ;
        RECT 134.910 188.040 135.290 188.090 ;
        RECT 131.210 187.760 135.290 188.040 ;
        RECT 131.210 187.710 131.590 187.760 ;
        RECT 134.910 187.710 135.290 187.760 ;
        RECT 6.700 186.385 9.560 186.765 ;
        RECT 39.150 186.385 42.010 186.765 ;
        RECT 71.600 186.385 74.460 186.765 ;
        RECT 104.050 186.385 106.910 186.765 ;
        RECT 137.355 186.725 137.735 187.105 ;
        RECT 139.395 186.725 139.775 187.105 ;
        RECT 141.180 186.725 141.560 187.105 ;
        RECT 6.700 185.625 9.560 186.005 ;
        RECT 39.150 185.625 42.010 186.005 ;
        RECT 71.600 185.625 74.460 186.005 ;
        RECT 104.050 185.625 106.910 186.005 ;
        RECT 0.240 185.225 0.620 185.605 ;
        RECT 4.160 185.225 4.540 185.605 ;
        RECT 35.140 185.395 35.520 185.445 ;
        RECT 37.560 185.395 37.940 185.445 ;
        RECT 35.140 185.115 37.940 185.395 ;
        RECT 35.140 185.065 35.520 185.115 ;
        RECT 37.560 185.065 37.940 185.115 ;
        RECT 67.590 185.395 67.970 185.445 ;
        RECT 70.010 185.395 70.390 185.445 ;
        RECT 67.590 185.115 70.390 185.395 ;
        RECT 67.590 185.065 67.970 185.115 ;
        RECT 70.010 185.065 70.390 185.115 ;
        RECT 100.040 185.395 100.420 185.445 ;
        RECT 102.460 185.395 102.840 185.445 ;
        RECT 100.040 185.115 102.840 185.395 ;
        RECT 100.040 185.065 100.420 185.115 ;
        RECT 102.460 185.065 102.840 185.115 ;
        RECT 132.490 185.395 132.870 185.445 ;
        RECT 134.910 185.395 135.290 185.445 ;
        RECT 132.490 185.115 135.290 185.395 ;
        RECT 132.490 185.065 132.870 185.115 ;
        RECT 134.910 185.065 135.290 185.115 ;
        RECT 6.700 183.785 9.560 184.165 ;
        RECT 39.150 183.785 42.010 184.165 ;
        RECT 71.600 183.785 74.460 184.165 ;
        RECT 104.050 183.785 106.910 184.165 ;
        RECT 137.355 183.725 137.735 184.105 ;
        RECT 139.395 183.725 139.775 184.105 ;
        RECT 141.180 183.725 141.560 184.105 ;
        RECT 36.420 183.555 36.800 183.605 ;
        RECT 37.560 183.555 37.940 183.605 ;
        RECT 36.420 183.275 37.940 183.555 ;
        RECT 36.420 183.225 36.800 183.275 ;
        RECT 37.560 183.225 37.940 183.275 ;
        RECT 68.870 183.555 69.250 183.605 ;
        RECT 70.010 183.555 70.390 183.605 ;
        RECT 68.870 183.275 70.390 183.555 ;
        RECT 68.870 183.225 69.250 183.275 ;
        RECT 70.010 183.225 70.390 183.275 ;
        RECT 101.320 183.555 101.700 183.605 ;
        RECT 102.460 183.555 102.840 183.605 ;
        RECT 101.320 183.275 102.840 183.555 ;
        RECT 101.320 183.225 101.700 183.275 ;
        RECT 102.460 183.225 102.840 183.275 ;
        RECT 133.770 183.555 134.150 183.605 ;
        RECT 134.910 183.555 135.290 183.605 ;
        RECT 133.770 183.275 135.290 183.555 ;
        RECT 133.770 183.225 134.150 183.275 ;
        RECT 134.910 183.225 135.290 183.275 ;
        RECT 0.240 182.225 0.620 182.605 ;
        RECT 4.160 182.225 4.540 182.605 ;
        RECT 6.700 181.945 9.560 182.325 ;
        RECT 39.150 181.945 42.010 182.325 ;
        RECT 71.600 181.945 74.460 182.325 ;
        RECT 104.050 181.945 106.910 182.325 ;
        RECT 37.560 181.385 38.080 181.765 ;
        RECT 70.010 181.385 70.530 181.765 ;
        RECT 102.460 181.385 102.980 181.765 ;
        RECT 134.910 181.385 135.430 181.765 ;
        RECT 137.355 180.725 137.735 181.105 ;
        RECT 139.395 180.725 139.775 181.105 ;
        RECT 141.180 180.725 141.560 181.105 ;
        RECT 0.240 179.225 0.620 179.605 ;
        RECT 4.160 179.225 4.540 179.605 ;
        RECT 0.240 176.225 0.620 176.605 ;
        RECT 137.355 174.725 137.735 175.105 ;
        RECT 139.395 174.725 139.775 175.105 ;
        RECT 141.180 174.725 141.560 175.105 ;
        RECT 0.240 173.225 0.620 173.605 ;
        RECT 4.160 173.225 4.540 173.605 ;
        RECT 37.060 172.820 37.940 173.200 ;
        RECT 69.510 172.820 70.390 173.200 ;
        RECT 101.960 172.820 102.840 173.200 ;
        RECT 134.410 172.820 135.290 173.200 ;
        RECT 6.700 172.260 9.560 172.640 ;
        RECT 39.150 172.260 42.010 172.640 ;
        RECT 71.600 172.260 74.460 172.640 ;
        RECT 104.050 172.260 106.910 172.640 ;
        RECT 137.355 171.725 137.735 172.105 ;
        RECT 139.395 171.725 139.775 172.105 ;
        RECT 141.180 171.725 141.560 172.105 ;
        RECT 35.780 171.310 36.160 171.360 ;
        RECT 37.560 171.310 37.940 171.360 ;
        RECT 35.780 171.030 37.940 171.310 ;
        RECT 35.780 170.980 36.160 171.030 ;
        RECT 37.560 170.980 37.940 171.030 ;
        RECT 68.230 171.310 68.610 171.360 ;
        RECT 70.010 171.310 70.390 171.360 ;
        RECT 68.230 171.030 70.390 171.310 ;
        RECT 68.230 170.980 68.610 171.030 ;
        RECT 70.010 170.980 70.390 171.030 ;
        RECT 100.680 171.310 101.060 171.360 ;
        RECT 102.460 171.310 102.840 171.360 ;
        RECT 100.680 171.030 102.840 171.310 ;
        RECT 100.680 170.980 101.060 171.030 ;
        RECT 102.460 170.980 102.840 171.030 ;
        RECT 133.130 171.310 133.510 171.360 ;
        RECT 134.910 171.310 135.290 171.360 ;
        RECT 133.130 171.030 135.290 171.310 ;
        RECT 133.130 170.980 133.510 171.030 ;
        RECT 134.910 170.980 135.290 171.030 ;
        RECT 0.240 170.225 0.620 170.605 ;
        RECT 4.160 170.225 4.540 170.605 ;
        RECT 6.700 170.420 9.560 170.800 ;
        RECT 39.150 170.420 42.010 170.800 ;
        RECT 71.600 170.420 74.460 170.800 ;
        RECT 104.050 170.420 106.910 170.800 ;
        RECT 34.500 169.465 34.880 169.515 ;
        RECT 37.560 169.465 37.940 169.515 ;
        RECT 34.500 169.185 37.940 169.465 ;
        RECT 34.500 169.135 34.880 169.185 ;
        RECT 37.560 169.135 37.940 169.185 ;
        RECT 66.950 169.465 67.330 169.515 ;
        RECT 70.010 169.465 70.390 169.515 ;
        RECT 66.950 169.185 70.390 169.465 ;
        RECT 66.950 169.135 67.330 169.185 ;
        RECT 70.010 169.135 70.390 169.185 ;
        RECT 99.400 169.465 99.780 169.515 ;
        RECT 102.460 169.465 102.840 169.515 ;
        RECT 99.400 169.185 102.840 169.465 ;
        RECT 99.400 169.135 99.780 169.185 ;
        RECT 102.460 169.135 102.840 169.185 ;
        RECT 131.850 169.465 132.230 169.515 ;
        RECT 134.910 169.465 135.290 169.515 ;
        RECT 131.850 169.185 135.290 169.465 ;
        RECT 131.850 169.135 132.230 169.185 ;
        RECT 134.910 169.135 135.290 169.185 ;
        RECT 6.700 168.575 9.560 168.955 ;
        RECT 39.150 168.575 42.010 168.955 ;
        RECT 71.600 168.575 74.460 168.955 ;
        RECT 104.050 168.575 106.910 168.955 ;
        RECT 137.355 168.725 137.735 169.105 ;
        RECT 139.395 168.725 139.775 169.105 ;
        RECT 141.180 168.725 141.560 169.105 ;
        RECT 6.700 167.815 9.560 168.195 ;
        RECT 39.150 167.815 42.010 168.195 ;
        RECT 71.600 167.815 74.460 168.195 ;
        RECT 104.050 167.815 106.910 168.195 ;
        RECT 0.240 167.225 0.620 167.605 ;
        RECT 4.160 167.225 4.540 167.605 ;
        RECT 33.220 166.825 33.600 166.875 ;
        RECT 37.560 166.825 37.940 166.875 ;
        RECT 33.220 166.545 37.940 166.825 ;
        RECT 33.220 166.495 33.600 166.545 ;
        RECT 37.560 166.495 37.940 166.545 ;
        RECT 65.670 166.825 66.050 166.875 ;
        RECT 70.010 166.825 70.390 166.875 ;
        RECT 65.670 166.545 70.390 166.825 ;
        RECT 65.670 166.495 66.050 166.545 ;
        RECT 70.010 166.495 70.390 166.545 ;
        RECT 98.120 166.825 98.500 166.875 ;
        RECT 102.460 166.825 102.840 166.875 ;
        RECT 98.120 166.545 102.840 166.825 ;
        RECT 98.120 166.495 98.500 166.545 ;
        RECT 102.460 166.495 102.840 166.545 ;
        RECT 130.570 166.825 130.950 166.875 ;
        RECT 134.910 166.825 135.290 166.875 ;
        RECT 130.570 166.545 135.290 166.825 ;
        RECT 130.570 166.495 130.950 166.545 ;
        RECT 134.910 166.495 135.290 166.545 ;
        RECT 6.700 165.935 9.560 166.315 ;
        RECT 39.150 165.935 42.010 166.315 ;
        RECT 71.600 165.935 74.460 166.315 ;
        RECT 104.050 165.935 106.910 166.315 ;
        RECT 137.355 165.725 137.735 166.105 ;
        RECT 139.395 165.725 139.775 166.105 ;
        RECT 141.180 165.725 141.560 166.105 ;
        RECT 31.940 164.985 32.320 165.035 ;
        RECT 37.560 164.985 37.940 165.035 ;
        RECT 31.940 164.705 37.940 164.985 ;
        RECT 31.940 164.655 32.320 164.705 ;
        RECT 37.560 164.655 37.940 164.705 ;
        RECT 64.390 164.985 64.770 165.035 ;
        RECT 70.010 164.985 70.390 165.035 ;
        RECT 64.390 164.705 70.390 164.985 ;
        RECT 64.390 164.655 64.770 164.705 ;
        RECT 70.010 164.655 70.390 164.705 ;
        RECT 96.840 164.985 97.220 165.035 ;
        RECT 102.460 164.985 102.840 165.035 ;
        RECT 96.840 164.705 102.840 164.985 ;
        RECT 96.840 164.655 97.220 164.705 ;
        RECT 102.460 164.655 102.840 164.705 ;
        RECT 129.290 164.985 129.670 165.035 ;
        RECT 134.910 164.985 135.290 165.035 ;
        RECT 129.290 164.705 135.290 164.985 ;
        RECT 129.290 164.655 129.670 164.705 ;
        RECT 134.910 164.655 135.290 164.705 ;
        RECT 0.240 164.225 0.620 164.605 ;
        RECT 4.160 164.225 4.540 164.605 ;
        RECT 6.700 164.095 9.560 164.475 ;
        RECT 39.150 164.095 42.010 164.475 ;
        RECT 71.600 164.095 74.460 164.475 ;
        RECT 104.050 164.095 106.910 164.475 ;
        RECT 30.660 163.140 31.040 163.190 ;
        RECT 37.560 163.140 37.940 163.190 ;
        RECT 30.660 162.860 37.940 163.140 ;
        RECT 30.660 162.810 31.040 162.860 ;
        RECT 37.560 162.810 37.940 162.860 ;
        RECT 63.110 163.140 63.490 163.190 ;
        RECT 70.010 163.140 70.390 163.190 ;
        RECT 63.110 162.860 70.390 163.140 ;
        RECT 63.110 162.810 63.490 162.860 ;
        RECT 70.010 162.810 70.390 162.860 ;
        RECT 95.560 163.140 95.940 163.190 ;
        RECT 102.460 163.140 102.840 163.190 ;
        RECT 95.560 162.860 102.840 163.140 ;
        RECT 95.560 162.810 95.940 162.860 ;
        RECT 102.460 162.810 102.840 162.860 ;
        RECT 128.010 163.140 128.390 163.190 ;
        RECT 134.910 163.140 135.290 163.190 ;
        RECT 128.010 162.860 135.290 163.140 ;
        RECT 128.010 162.810 128.390 162.860 ;
        RECT 134.910 162.810 135.290 162.860 ;
        RECT 137.355 162.725 137.735 163.105 ;
        RECT 139.395 162.725 139.775 163.105 ;
        RECT 141.180 162.725 141.560 163.105 ;
        RECT 6.700 162.250 9.560 162.630 ;
        RECT 39.150 162.250 42.010 162.630 ;
        RECT 71.600 162.250 74.460 162.630 ;
        RECT 104.050 162.250 106.910 162.630 ;
        RECT 0.240 161.225 0.620 161.605 ;
        RECT 4.160 161.225 4.540 161.605 ;
        RECT 6.700 161.490 9.560 161.870 ;
        RECT 39.150 161.490 42.010 161.870 ;
        RECT 71.600 161.490 74.460 161.870 ;
        RECT 104.050 161.490 106.910 161.870 ;
        RECT 29.380 160.500 29.760 160.550 ;
        RECT 37.560 160.500 37.940 160.550 ;
        RECT 29.380 160.220 37.940 160.500 ;
        RECT 29.380 160.170 29.760 160.220 ;
        RECT 37.560 160.170 37.940 160.220 ;
        RECT 61.830 160.500 62.210 160.550 ;
        RECT 70.010 160.500 70.390 160.550 ;
        RECT 61.830 160.220 70.390 160.500 ;
        RECT 61.830 160.170 62.210 160.220 ;
        RECT 70.010 160.170 70.390 160.220 ;
        RECT 94.280 160.500 94.660 160.550 ;
        RECT 102.460 160.500 102.840 160.550 ;
        RECT 94.280 160.220 102.840 160.500 ;
        RECT 94.280 160.170 94.660 160.220 ;
        RECT 102.460 160.170 102.840 160.220 ;
        RECT 126.730 160.500 127.110 160.550 ;
        RECT 134.910 160.500 135.290 160.550 ;
        RECT 126.730 160.220 135.290 160.500 ;
        RECT 126.730 160.170 127.110 160.220 ;
        RECT 134.910 160.170 135.290 160.220 ;
        RECT 6.700 159.610 9.560 159.990 ;
        RECT 39.150 159.610 42.010 159.990 ;
        RECT 71.600 159.610 74.460 159.990 ;
        RECT 104.050 159.610 106.910 159.990 ;
        RECT 137.355 159.725 137.735 160.105 ;
        RECT 139.395 159.725 139.775 160.105 ;
        RECT 141.180 159.725 141.560 160.105 ;
        RECT 28.100 158.660 28.480 158.710 ;
        RECT 37.560 158.660 37.940 158.710 ;
        RECT 0.240 158.225 0.620 158.605 ;
        RECT 4.160 158.225 4.540 158.605 ;
        RECT 28.100 158.380 37.940 158.660 ;
        RECT 28.100 158.330 28.480 158.380 ;
        RECT 37.560 158.330 37.940 158.380 ;
        RECT 60.550 158.660 60.930 158.710 ;
        RECT 70.010 158.660 70.390 158.710 ;
        RECT 60.550 158.380 70.390 158.660 ;
        RECT 60.550 158.330 60.930 158.380 ;
        RECT 70.010 158.330 70.390 158.380 ;
        RECT 93.000 158.660 93.380 158.710 ;
        RECT 102.460 158.660 102.840 158.710 ;
        RECT 93.000 158.380 102.840 158.660 ;
        RECT 93.000 158.330 93.380 158.380 ;
        RECT 102.460 158.330 102.840 158.380 ;
        RECT 125.450 158.660 125.830 158.710 ;
        RECT 134.910 158.660 135.290 158.710 ;
        RECT 125.450 158.380 135.290 158.660 ;
        RECT 125.450 158.330 125.830 158.380 ;
        RECT 134.910 158.330 135.290 158.380 ;
        RECT 6.700 157.770 9.560 158.150 ;
        RECT 39.150 157.770 42.010 158.150 ;
        RECT 71.600 157.770 74.460 158.150 ;
        RECT 104.050 157.770 106.910 158.150 ;
        RECT 6.700 157.050 9.560 157.430 ;
        RECT 39.150 157.050 42.010 157.430 ;
        RECT 71.600 157.050 74.460 157.430 ;
        RECT 104.050 157.050 106.910 157.430 ;
        RECT 28.740 156.820 29.120 156.870 ;
        RECT 37.560 156.820 37.940 156.870 ;
        RECT 28.740 156.540 37.940 156.820 ;
        RECT 28.740 156.490 29.120 156.540 ;
        RECT 37.560 156.490 37.940 156.540 ;
        RECT 61.190 156.820 61.570 156.870 ;
        RECT 70.010 156.820 70.390 156.870 ;
        RECT 61.190 156.540 70.390 156.820 ;
        RECT 61.190 156.490 61.570 156.540 ;
        RECT 70.010 156.490 70.390 156.540 ;
        RECT 93.640 156.820 94.020 156.870 ;
        RECT 102.460 156.820 102.840 156.870 ;
        RECT 93.640 156.540 102.840 156.820 ;
        RECT 93.640 156.490 94.020 156.540 ;
        RECT 102.460 156.490 102.840 156.540 ;
        RECT 126.090 156.820 126.470 156.870 ;
        RECT 134.910 156.820 135.290 156.870 ;
        RECT 126.090 156.540 135.290 156.820 ;
        RECT 126.090 156.490 126.470 156.540 ;
        RECT 134.910 156.490 135.290 156.540 ;
        RECT 0.240 154.840 0.620 155.220 ;
        RECT 4.160 154.840 4.540 155.220 ;
        RECT 6.700 155.210 9.560 155.590 ;
        RECT 39.150 155.210 42.010 155.590 ;
        RECT 71.600 155.210 74.460 155.590 ;
        RECT 104.050 155.210 106.910 155.590 ;
        RECT 30.020 154.980 30.400 155.030 ;
        RECT 37.560 154.980 37.940 155.030 ;
        RECT 30.020 154.700 37.940 154.980 ;
        RECT 30.020 154.650 30.400 154.700 ;
        RECT 37.560 154.650 37.940 154.700 ;
        RECT 62.470 154.980 62.850 155.030 ;
        RECT 70.010 154.980 70.390 155.030 ;
        RECT 62.470 154.700 70.390 154.980 ;
        RECT 62.470 154.650 62.850 154.700 ;
        RECT 70.010 154.650 70.390 154.700 ;
        RECT 94.920 154.980 95.300 155.030 ;
        RECT 102.460 154.980 102.840 155.030 ;
        RECT 94.920 154.700 102.840 154.980 ;
        RECT 94.920 154.650 95.300 154.700 ;
        RECT 102.460 154.650 102.840 154.700 ;
        RECT 127.370 154.980 127.750 155.030 ;
        RECT 134.910 154.980 135.290 155.030 ;
        RECT 127.370 154.700 135.290 154.980 ;
        RECT 127.370 154.650 127.750 154.700 ;
        RECT 134.910 154.650 135.290 154.700 ;
        RECT 6.700 153.325 9.560 153.705 ;
        RECT 39.150 153.325 42.010 153.705 ;
        RECT 71.600 153.325 74.460 153.705 ;
        RECT 104.050 153.325 106.910 153.705 ;
        RECT 137.355 153.340 137.735 153.720 ;
        RECT 139.395 153.340 139.775 153.720 ;
        RECT 141.180 153.340 141.560 153.720 ;
        RECT 6.700 152.565 9.560 152.945 ;
        RECT 39.150 152.565 42.010 152.945 ;
        RECT 71.600 152.565 74.460 152.945 ;
        RECT 104.050 152.565 106.910 152.945 ;
        RECT 31.300 152.335 31.680 152.385 ;
        RECT 37.560 152.335 37.940 152.385 ;
        RECT 0.240 151.840 0.620 152.220 ;
        RECT 4.160 151.840 4.540 152.220 ;
        RECT 31.300 152.055 37.940 152.335 ;
        RECT 31.300 152.005 31.680 152.055 ;
        RECT 37.560 152.005 37.940 152.055 ;
        RECT 63.750 152.335 64.130 152.385 ;
        RECT 70.010 152.335 70.390 152.385 ;
        RECT 63.750 152.055 70.390 152.335 ;
        RECT 63.750 152.005 64.130 152.055 ;
        RECT 70.010 152.005 70.390 152.055 ;
        RECT 96.200 152.335 96.580 152.385 ;
        RECT 102.460 152.335 102.840 152.385 ;
        RECT 96.200 152.055 102.840 152.335 ;
        RECT 96.200 152.005 96.580 152.055 ;
        RECT 102.460 152.005 102.840 152.055 ;
        RECT 128.650 152.335 129.030 152.385 ;
        RECT 134.910 152.335 135.290 152.385 ;
        RECT 128.650 152.055 135.290 152.335 ;
        RECT 128.650 152.005 129.030 152.055 ;
        RECT 134.910 152.005 135.290 152.055 ;
        RECT 6.700 150.725 9.560 151.105 ;
        RECT 39.150 150.725 42.010 151.105 ;
        RECT 71.600 150.725 74.460 151.105 ;
        RECT 104.050 150.725 106.910 151.105 ;
        RECT 32.580 150.495 32.960 150.545 ;
        RECT 37.560 150.495 37.940 150.545 ;
        RECT 32.580 150.215 37.940 150.495 ;
        RECT 32.580 150.165 32.960 150.215 ;
        RECT 37.560 150.165 37.940 150.215 ;
        RECT 65.030 150.495 65.410 150.545 ;
        RECT 70.010 150.495 70.390 150.545 ;
        RECT 65.030 150.215 70.390 150.495 ;
        RECT 65.030 150.165 65.410 150.215 ;
        RECT 70.010 150.165 70.390 150.215 ;
        RECT 97.480 150.495 97.860 150.545 ;
        RECT 102.460 150.495 102.840 150.545 ;
        RECT 97.480 150.215 102.840 150.495 ;
        RECT 97.480 150.165 97.860 150.215 ;
        RECT 102.460 150.165 102.840 150.215 ;
        RECT 129.930 150.495 130.310 150.545 ;
        RECT 134.910 150.495 135.290 150.545 ;
        RECT 129.930 150.215 135.290 150.495 ;
        RECT 137.355 150.340 137.735 150.720 ;
        RECT 139.395 150.340 139.775 150.720 ;
        RECT 141.180 150.340 141.560 150.720 ;
        RECT 129.930 150.165 130.310 150.215 ;
        RECT 134.910 150.165 135.290 150.215 ;
        RECT 0.240 148.840 0.620 149.220 ;
        RECT 4.160 148.840 4.540 149.220 ;
        RECT 6.700 148.885 9.560 149.265 ;
        RECT 39.150 148.885 42.010 149.265 ;
        RECT 71.600 148.885 74.460 149.265 ;
        RECT 104.050 148.885 106.910 149.265 ;
        RECT 33.860 148.655 34.240 148.705 ;
        RECT 37.560 148.655 37.940 148.705 ;
        RECT 33.860 148.375 37.940 148.655 ;
        RECT 33.860 148.325 34.240 148.375 ;
        RECT 37.560 148.325 37.940 148.375 ;
        RECT 66.310 148.655 66.690 148.705 ;
        RECT 70.010 148.655 70.390 148.705 ;
        RECT 66.310 148.375 70.390 148.655 ;
        RECT 66.310 148.325 66.690 148.375 ;
        RECT 70.010 148.325 70.390 148.375 ;
        RECT 98.760 148.655 99.140 148.705 ;
        RECT 102.460 148.655 102.840 148.705 ;
        RECT 98.760 148.375 102.840 148.655 ;
        RECT 98.760 148.325 99.140 148.375 ;
        RECT 102.460 148.325 102.840 148.375 ;
        RECT 131.210 148.655 131.590 148.705 ;
        RECT 134.910 148.655 135.290 148.705 ;
        RECT 131.210 148.375 135.290 148.655 ;
        RECT 131.210 148.325 131.590 148.375 ;
        RECT 134.910 148.325 135.290 148.375 ;
        RECT 6.700 147.000 9.560 147.380 ;
        RECT 39.150 147.000 42.010 147.380 ;
        RECT 71.600 147.000 74.460 147.380 ;
        RECT 104.050 147.000 106.910 147.380 ;
        RECT 137.355 147.340 137.735 147.720 ;
        RECT 139.395 147.340 139.775 147.720 ;
        RECT 141.180 147.340 141.560 147.720 ;
        RECT 6.700 146.240 9.560 146.620 ;
        RECT 39.150 146.240 42.010 146.620 ;
        RECT 71.600 146.240 74.460 146.620 ;
        RECT 104.050 146.240 106.910 146.620 ;
        RECT 0.240 145.840 0.620 146.220 ;
        RECT 4.160 145.840 4.540 146.220 ;
        RECT 35.140 146.010 35.520 146.060 ;
        RECT 37.560 146.010 37.940 146.060 ;
        RECT 35.140 145.730 37.940 146.010 ;
        RECT 35.140 145.680 35.520 145.730 ;
        RECT 37.560 145.680 37.940 145.730 ;
        RECT 67.590 146.010 67.970 146.060 ;
        RECT 70.010 146.010 70.390 146.060 ;
        RECT 67.590 145.730 70.390 146.010 ;
        RECT 67.590 145.680 67.970 145.730 ;
        RECT 70.010 145.680 70.390 145.730 ;
        RECT 100.040 146.010 100.420 146.060 ;
        RECT 102.460 146.010 102.840 146.060 ;
        RECT 100.040 145.730 102.840 146.010 ;
        RECT 100.040 145.680 100.420 145.730 ;
        RECT 102.460 145.680 102.840 145.730 ;
        RECT 132.490 146.010 132.870 146.060 ;
        RECT 134.910 146.010 135.290 146.060 ;
        RECT 132.490 145.730 135.290 146.010 ;
        RECT 132.490 145.680 132.870 145.730 ;
        RECT 134.910 145.680 135.290 145.730 ;
        RECT 6.700 144.400 9.560 144.780 ;
        RECT 39.150 144.400 42.010 144.780 ;
        RECT 71.600 144.400 74.460 144.780 ;
        RECT 104.050 144.400 106.910 144.780 ;
        RECT 137.355 144.340 137.735 144.720 ;
        RECT 139.395 144.340 139.775 144.720 ;
        RECT 141.180 144.340 141.560 144.720 ;
        RECT 36.420 144.170 36.800 144.220 ;
        RECT 37.560 144.170 37.940 144.220 ;
        RECT 36.420 143.890 37.940 144.170 ;
        RECT 36.420 143.840 36.800 143.890 ;
        RECT 37.560 143.840 37.940 143.890 ;
        RECT 68.870 144.170 69.250 144.220 ;
        RECT 70.010 144.170 70.390 144.220 ;
        RECT 68.870 143.890 70.390 144.170 ;
        RECT 68.870 143.840 69.250 143.890 ;
        RECT 70.010 143.840 70.390 143.890 ;
        RECT 101.320 144.170 101.700 144.220 ;
        RECT 102.460 144.170 102.840 144.220 ;
        RECT 101.320 143.890 102.840 144.170 ;
        RECT 101.320 143.840 101.700 143.890 ;
        RECT 102.460 143.840 102.840 143.890 ;
        RECT 133.770 144.170 134.150 144.220 ;
        RECT 134.910 144.170 135.290 144.220 ;
        RECT 133.770 143.890 135.290 144.170 ;
        RECT 133.770 143.840 134.150 143.890 ;
        RECT 134.910 143.840 135.290 143.890 ;
        RECT 0.240 142.840 0.620 143.220 ;
        RECT 4.160 142.840 4.540 143.220 ;
        RECT 6.700 142.560 9.560 142.940 ;
        RECT 39.150 142.560 42.010 142.940 ;
        RECT 71.600 142.560 74.460 142.940 ;
        RECT 104.050 142.560 106.910 142.940 ;
        RECT 37.560 142.000 38.080 142.380 ;
        RECT 70.010 142.000 70.530 142.380 ;
        RECT 102.460 142.000 102.980 142.380 ;
        RECT 134.910 142.000 135.430 142.380 ;
        RECT 137.355 141.340 137.735 141.720 ;
        RECT 139.395 141.340 139.775 141.720 ;
        RECT 141.180 141.340 141.560 141.720 ;
        RECT 0.240 139.840 0.620 140.220 ;
        RECT 4.160 139.840 4.540 140.220 ;
        RECT 0.240 136.840 0.620 137.220 ;
        RECT 137.355 135.340 137.735 135.720 ;
        RECT 139.395 135.340 139.775 135.720 ;
        RECT 141.180 135.340 141.560 135.720 ;
        RECT 0.240 133.840 0.620 134.220 ;
        RECT 4.160 133.840 4.540 134.220 ;
        RECT 37.060 133.435 37.940 133.815 ;
        RECT 69.510 133.435 70.390 133.815 ;
        RECT 101.960 133.435 102.840 133.815 ;
        RECT 134.410 133.435 135.290 133.815 ;
        RECT 6.700 132.875 9.560 133.255 ;
        RECT 39.150 132.875 42.010 133.255 ;
        RECT 71.600 132.875 74.460 133.255 ;
        RECT 104.050 132.875 106.910 133.255 ;
        RECT 137.355 132.340 137.735 132.720 ;
        RECT 139.395 132.340 139.775 132.720 ;
        RECT 141.180 132.340 141.560 132.720 ;
        RECT 35.780 131.925 36.160 131.975 ;
        RECT 37.560 131.925 37.940 131.975 ;
        RECT 35.780 131.645 37.940 131.925 ;
        RECT 35.780 131.595 36.160 131.645 ;
        RECT 37.560 131.595 37.940 131.645 ;
        RECT 68.230 131.925 68.610 131.975 ;
        RECT 70.010 131.925 70.390 131.975 ;
        RECT 68.230 131.645 70.390 131.925 ;
        RECT 68.230 131.595 68.610 131.645 ;
        RECT 70.010 131.595 70.390 131.645 ;
        RECT 100.680 131.925 101.060 131.975 ;
        RECT 102.460 131.925 102.840 131.975 ;
        RECT 100.680 131.645 102.840 131.925 ;
        RECT 100.680 131.595 101.060 131.645 ;
        RECT 102.460 131.595 102.840 131.645 ;
        RECT 133.130 131.925 133.510 131.975 ;
        RECT 134.910 131.925 135.290 131.975 ;
        RECT 133.130 131.645 135.290 131.925 ;
        RECT 133.130 131.595 133.510 131.645 ;
        RECT 134.910 131.595 135.290 131.645 ;
        RECT 0.240 130.840 0.620 131.220 ;
        RECT 4.160 130.840 4.540 131.220 ;
        RECT 6.700 131.035 9.560 131.415 ;
        RECT 39.150 131.035 42.010 131.415 ;
        RECT 71.600 131.035 74.460 131.415 ;
        RECT 104.050 131.035 106.910 131.415 ;
        RECT 34.500 130.080 34.880 130.130 ;
        RECT 37.560 130.080 37.940 130.130 ;
        RECT 34.500 129.800 37.940 130.080 ;
        RECT 34.500 129.750 34.880 129.800 ;
        RECT 37.560 129.750 37.940 129.800 ;
        RECT 66.950 130.080 67.330 130.130 ;
        RECT 70.010 130.080 70.390 130.130 ;
        RECT 66.950 129.800 70.390 130.080 ;
        RECT 66.950 129.750 67.330 129.800 ;
        RECT 70.010 129.750 70.390 129.800 ;
        RECT 99.400 130.080 99.780 130.130 ;
        RECT 102.460 130.080 102.840 130.130 ;
        RECT 99.400 129.800 102.840 130.080 ;
        RECT 99.400 129.750 99.780 129.800 ;
        RECT 102.460 129.750 102.840 129.800 ;
        RECT 131.850 130.080 132.230 130.130 ;
        RECT 134.910 130.080 135.290 130.130 ;
        RECT 131.850 129.800 135.290 130.080 ;
        RECT 131.850 129.750 132.230 129.800 ;
        RECT 134.910 129.750 135.290 129.800 ;
        RECT 6.700 129.190 9.560 129.570 ;
        RECT 39.150 129.190 42.010 129.570 ;
        RECT 71.600 129.190 74.460 129.570 ;
        RECT 104.050 129.190 106.910 129.570 ;
        RECT 137.355 129.340 137.735 129.720 ;
        RECT 139.395 129.340 139.775 129.720 ;
        RECT 141.180 129.340 141.560 129.720 ;
        RECT 6.700 128.430 9.560 128.810 ;
        RECT 39.150 128.430 42.010 128.810 ;
        RECT 71.600 128.430 74.460 128.810 ;
        RECT 104.050 128.430 106.910 128.810 ;
        RECT 0.240 127.840 0.620 128.220 ;
        RECT 4.160 127.840 4.540 128.220 ;
        RECT 33.220 127.440 33.600 127.490 ;
        RECT 37.560 127.440 37.940 127.490 ;
        RECT 33.220 127.160 37.940 127.440 ;
        RECT 33.220 127.110 33.600 127.160 ;
        RECT 37.560 127.110 37.940 127.160 ;
        RECT 65.670 127.440 66.050 127.490 ;
        RECT 70.010 127.440 70.390 127.490 ;
        RECT 65.670 127.160 70.390 127.440 ;
        RECT 65.670 127.110 66.050 127.160 ;
        RECT 70.010 127.110 70.390 127.160 ;
        RECT 98.120 127.440 98.500 127.490 ;
        RECT 102.460 127.440 102.840 127.490 ;
        RECT 98.120 127.160 102.840 127.440 ;
        RECT 98.120 127.110 98.500 127.160 ;
        RECT 102.460 127.110 102.840 127.160 ;
        RECT 130.570 127.440 130.950 127.490 ;
        RECT 134.910 127.440 135.290 127.490 ;
        RECT 130.570 127.160 135.290 127.440 ;
        RECT 130.570 127.110 130.950 127.160 ;
        RECT 134.910 127.110 135.290 127.160 ;
        RECT 6.700 126.550 9.560 126.930 ;
        RECT 39.150 126.550 42.010 126.930 ;
        RECT 71.600 126.550 74.460 126.930 ;
        RECT 104.050 126.550 106.910 126.930 ;
        RECT 137.355 126.340 137.735 126.720 ;
        RECT 139.395 126.340 139.775 126.720 ;
        RECT 141.180 126.340 141.560 126.720 ;
        RECT 31.940 125.600 32.320 125.650 ;
        RECT 37.560 125.600 37.940 125.650 ;
        RECT 31.940 125.320 37.940 125.600 ;
        RECT 31.940 125.270 32.320 125.320 ;
        RECT 37.560 125.270 37.940 125.320 ;
        RECT 64.390 125.600 64.770 125.650 ;
        RECT 70.010 125.600 70.390 125.650 ;
        RECT 64.390 125.320 70.390 125.600 ;
        RECT 64.390 125.270 64.770 125.320 ;
        RECT 70.010 125.270 70.390 125.320 ;
        RECT 96.840 125.600 97.220 125.650 ;
        RECT 102.460 125.600 102.840 125.650 ;
        RECT 96.840 125.320 102.840 125.600 ;
        RECT 96.840 125.270 97.220 125.320 ;
        RECT 102.460 125.270 102.840 125.320 ;
        RECT 129.290 125.600 129.670 125.650 ;
        RECT 134.910 125.600 135.290 125.650 ;
        RECT 129.290 125.320 135.290 125.600 ;
        RECT 129.290 125.270 129.670 125.320 ;
        RECT 134.910 125.270 135.290 125.320 ;
        RECT 0.240 124.840 0.620 125.220 ;
        RECT 4.160 124.840 4.540 125.220 ;
        RECT 6.700 124.710 9.560 125.090 ;
        RECT 39.150 124.710 42.010 125.090 ;
        RECT 71.600 124.710 74.460 125.090 ;
        RECT 104.050 124.710 106.910 125.090 ;
        RECT 30.660 123.755 31.040 123.805 ;
        RECT 37.560 123.755 37.940 123.805 ;
        RECT 30.660 123.475 37.940 123.755 ;
        RECT 30.660 123.425 31.040 123.475 ;
        RECT 37.560 123.425 37.940 123.475 ;
        RECT 63.110 123.755 63.490 123.805 ;
        RECT 70.010 123.755 70.390 123.805 ;
        RECT 63.110 123.475 70.390 123.755 ;
        RECT 63.110 123.425 63.490 123.475 ;
        RECT 70.010 123.425 70.390 123.475 ;
        RECT 95.560 123.755 95.940 123.805 ;
        RECT 102.460 123.755 102.840 123.805 ;
        RECT 95.560 123.475 102.840 123.755 ;
        RECT 95.560 123.425 95.940 123.475 ;
        RECT 102.460 123.425 102.840 123.475 ;
        RECT 128.010 123.755 128.390 123.805 ;
        RECT 134.910 123.755 135.290 123.805 ;
        RECT 128.010 123.475 135.290 123.755 ;
        RECT 128.010 123.425 128.390 123.475 ;
        RECT 134.910 123.425 135.290 123.475 ;
        RECT 137.355 123.340 137.735 123.720 ;
        RECT 139.395 123.340 139.775 123.720 ;
        RECT 141.180 123.340 141.560 123.720 ;
        RECT 6.700 122.865 9.560 123.245 ;
        RECT 39.150 122.865 42.010 123.245 ;
        RECT 71.600 122.865 74.460 123.245 ;
        RECT 104.050 122.865 106.910 123.245 ;
        RECT 0.240 121.840 0.620 122.220 ;
        RECT 4.160 121.840 4.540 122.220 ;
        RECT 6.700 122.105 9.560 122.485 ;
        RECT 39.150 122.105 42.010 122.485 ;
        RECT 71.600 122.105 74.460 122.485 ;
        RECT 104.050 122.105 106.910 122.485 ;
        RECT 29.380 121.115 29.760 121.165 ;
        RECT 37.560 121.115 37.940 121.165 ;
        RECT 29.380 120.835 37.940 121.115 ;
        RECT 29.380 120.785 29.760 120.835 ;
        RECT 37.560 120.785 37.940 120.835 ;
        RECT 61.830 121.115 62.210 121.165 ;
        RECT 70.010 121.115 70.390 121.165 ;
        RECT 61.830 120.835 70.390 121.115 ;
        RECT 61.830 120.785 62.210 120.835 ;
        RECT 70.010 120.785 70.390 120.835 ;
        RECT 94.280 121.115 94.660 121.165 ;
        RECT 102.460 121.115 102.840 121.165 ;
        RECT 94.280 120.835 102.840 121.115 ;
        RECT 94.280 120.785 94.660 120.835 ;
        RECT 102.460 120.785 102.840 120.835 ;
        RECT 126.730 121.115 127.110 121.165 ;
        RECT 134.910 121.115 135.290 121.165 ;
        RECT 126.730 120.835 135.290 121.115 ;
        RECT 126.730 120.785 127.110 120.835 ;
        RECT 134.910 120.785 135.290 120.835 ;
        RECT 6.700 120.225 9.560 120.605 ;
        RECT 39.150 120.225 42.010 120.605 ;
        RECT 71.600 120.225 74.460 120.605 ;
        RECT 104.050 120.225 106.910 120.605 ;
        RECT 137.355 120.340 137.735 120.720 ;
        RECT 139.395 120.340 139.775 120.720 ;
        RECT 141.180 120.340 141.560 120.720 ;
        RECT 28.100 119.275 28.480 119.325 ;
        RECT 37.560 119.275 37.940 119.325 ;
        RECT 0.240 118.840 0.620 119.220 ;
        RECT 4.160 118.840 4.540 119.220 ;
        RECT 28.100 118.995 37.940 119.275 ;
        RECT 28.100 118.945 28.480 118.995 ;
        RECT 37.560 118.945 37.940 118.995 ;
        RECT 60.550 119.275 60.930 119.325 ;
        RECT 70.010 119.275 70.390 119.325 ;
        RECT 60.550 118.995 70.390 119.275 ;
        RECT 60.550 118.945 60.930 118.995 ;
        RECT 70.010 118.945 70.390 118.995 ;
        RECT 93.000 119.275 93.380 119.325 ;
        RECT 102.460 119.275 102.840 119.325 ;
        RECT 93.000 118.995 102.840 119.275 ;
        RECT 93.000 118.945 93.380 118.995 ;
        RECT 102.460 118.945 102.840 118.995 ;
        RECT 125.450 119.275 125.830 119.325 ;
        RECT 134.910 119.275 135.290 119.325 ;
        RECT 125.450 118.995 135.290 119.275 ;
        RECT 125.450 118.945 125.830 118.995 ;
        RECT 134.910 118.945 135.290 118.995 ;
        RECT 6.700 118.385 9.560 118.765 ;
        RECT 39.150 118.385 42.010 118.765 ;
        RECT 71.600 118.385 74.460 118.765 ;
        RECT 104.050 118.385 106.910 118.765 ;
        RECT 6.700 117.665 9.560 118.045 ;
        RECT 39.150 117.665 42.010 118.045 ;
        RECT 71.600 117.665 74.460 118.045 ;
        RECT 104.050 117.665 106.910 118.045 ;
        RECT 28.740 117.435 29.120 117.485 ;
        RECT 37.560 117.435 37.940 117.485 ;
        RECT 28.740 117.155 37.940 117.435 ;
        RECT 28.740 117.105 29.120 117.155 ;
        RECT 37.560 117.105 37.940 117.155 ;
        RECT 61.190 117.435 61.570 117.485 ;
        RECT 70.010 117.435 70.390 117.485 ;
        RECT 61.190 117.155 70.390 117.435 ;
        RECT 61.190 117.105 61.570 117.155 ;
        RECT 70.010 117.105 70.390 117.155 ;
        RECT 93.640 117.435 94.020 117.485 ;
        RECT 102.460 117.435 102.840 117.485 ;
        RECT 93.640 117.155 102.840 117.435 ;
        RECT 93.640 117.105 94.020 117.155 ;
        RECT 102.460 117.105 102.840 117.155 ;
        RECT 126.090 117.435 126.470 117.485 ;
        RECT 134.910 117.435 135.290 117.485 ;
        RECT 126.090 117.155 135.290 117.435 ;
        RECT 126.090 117.105 126.470 117.155 ;
        RECT 134.910 117.105 135.290 117.155 ;
        RECT 0.240 115.455 0.620 115.835 ;
        RECT 4.160 115.455 4.540 115.835 ;
        RECT 6.700 115.825 9.560 116.205 ;
        RECT 39.150 115.825 42.010 116.205 ;
        RECT 71.600 115.825 74.460 116.205 ;
        RECT 104.050 115.825 106.910 116.205 ;
        RECT 30.020 115.595 30.400 115.645 ;
        RECT 37.560 115.595 37.940 115.645 ;
        RECT 30.020 115.315 37.940 115.595 ;
        RECT 30.020 115.265 30.400 115.315 ;
        RECT 37.560 115.265 37.940 115.315 ;
        RECT 62.470 115.595 62.850 115.645 ;
        RECT 70.010 115.595 70.390 115.645 ;
        RECT 62.470 115.315 70.390 115.595 ;
        RECT 62.470 115.265 62.850 115.315 ;
        RECT 70.010 115.265 70.390 115.315 ;
        RECT 94.920 115.595 95.300 115.645 ;
        RECT 102.460 115.595 102.840 115.645 ;
        RECT 94.920 115.315 102.840 115.595 ;
        RECT 94.920 115.265 95.300 115.315 ;
        RECT 102.460 115.265 102.840 115.315 ;
        RECT 127.370 115.595 127.750 115.645 ;
        RECT 134.910 115.595 135.290 115.645 ;
        RECT 127.370 115.315 135.290 115.595 ;
        RECT 127.370 115.265 127.750 115.315 ;
        RECT 134.910 115.265 135.290 115.315 ;
        RECT 6.700 113.940 9.560 114.320 ;
        RECT 39.150 113.940 42.010 114.320 ;
        RECT 71.600 113.940 74.460 114.320 ;
        RECT 104.050 113.940 106.910 114.320 ;
        RECT 137.355 113.955 137.735 114.335 ;
        RECT 139.395 113.955 139.775 114.335 ;
        RECT 141.180 113.955 141.560 114.335 ;
        RECT 6.700 113.180 9.560 113.560 ;
        RECT 39.150 113.180 42.010 113.560 ;
        RECT 71.600 113.180 74.460 113.560 ;
        RECT 104.050 113.180 106.910 113.560 ;
        RECT 31.300 112.950 31.680 113.000 ;
        RECT 37.560 112.950 37.940 113.000 ;
        RECT 0.240 112.455 0.620 112.835 ;
        RECT 4.160 112.455 4.540 112.835 ;
        RECT 31.300 112.670 37.940 112.950 ;
        RECT 31.300 112.620 31.680 112.670 ;
        RECT 37.560 112.620 37.940 112.670 ;
        RECT 63.750 112.950 64.130 113.000 ;
        RECT 70.010 112.950 70.390 113.000 ;
        RECT 63.750 112.670 70.390 112.950 ;
        RECT 63.750 112.620 64.130 112.670 ;
        RECT 70.010 112.620 70.390 112.670 ;
        RECT 96.200 112.950 96.580 113.000 ;
        RECT 102.460 112.950 102.840 113.000 ;
        RECT 96.200 112.670 102.840 112.950 ;
        RECT 96.200 112.620 96.580 112.670 ;
        RECT 102.460 112.620 102.840 112.670 ;
        RECT 128.650 112.950 129.030 113.000 ;
        RECT 134.910 112.950 135.290 113.000 ;
        RECT 128.650 112.670 135.290 112.950 ;
        RECT 128.650 112.620 129.030 112.670 ;
        RECT 134.910 112.620 135.290 112.670 ;
        RECT 6.700 111.340 9.560 111.720 ;
        RECT 39.150 111.340 42.010 111.720 ;
        RECT 71.600 111.340 74.460 111.720 ;
        RECT 104.050 111.340 106.910 111.720 ;
        RECT 32.580 111.110 32.960 111.160 ;
        RECT 37.560 111.110 37.940 111.160 ;
        RECT 32.580 110.830 37.940 111.110 ;
        RECT 32.580 110.780 32.960 110.830 ;
        RECT 37.560 110.780 37.940 110.830 ;
        RECT 65.030 111.110 65.410 111.160 ;
        RECT 70.010 111.110 70.390 111.160 ;
        RECT 65.030 110.830 70.390 111.110 ;
        RECT 65.030 110.780 65.410 110.830 ;
        RECT 70.010 110.780 70.390 110.830 ;
        RECT 97.480 111.110 97.860 111.160 ;
        RECT 102.460 111.110 102.840 111.160 ;
        RECT 97.480 110.830 102.840 111.110 ;
        RECT 97.480 110.780 97.860 110.830 ;
        RECT 102.460 110.780 102.840 110.830 ;
        RECT 129.930 111.110 130.310 111.160 ;
        RECT 134.910 111.110 135.290 111.160 ;
        RECT 129.930 110.830 135.290 111.110 ;
        RECT 137.355 110.955 137.735 111.335 ;
        RECT 139.395 110.955 139.775 111.335 ;
        RECT 141.180 110.955 141.560 111.335 ;
        RECT 129.930 110.780 130.310 110.830 ;
        RECT 134.910 110.780 135.290 110.830 ;
        RECT 0.240 109.455 0.620 109.835 ;
        RECT 4.160 109.455 4.540 109.835 ;
        RECT 6.700 109.500 9.560 109.880 ;
        RECT 39.150 109.500 42.010 109.880 ;
        RECT 71.600 109.500 74.460 109.880 ;
        RECT 104.050 109.500 106.910 109.880 ;
        RECT 33.860 109.270 34.240 109.320 ;
        RECT 37.560 109.270 37.940 109.320 ;
        RECT 33.860 108.990 37.940 109.270 ;
        RECT 33.860 108.940 34.240 108.990 ;
        RECT 37.560 108.940 37.940 108.990 ;
        RECT 66.310 109.270 66.690 109.320 ;
        RECT 70.010 109.270 70.390 109.320 ;
        RECT 66.310 108.990 70.390 109.270 ;
        RECT 66.310 108.940 66.690 108.990 ;
        RECT 70.010 108.940 70.390 108.990 ;
        RECT 98.760 109.270 99.140 109.320 ;
        RECT 102.460 109.270 102.840 109.320 ;
        RECT 98.760 108.990 102.840 109.270 ;
        RECT 98.760 108.940 99.140 108.990 ;
        RECT 102.460 108.940 102.840 108.990 ;
        RECT 131.210 109.270 131.590 109.320 ;
        RECT 134.910 109.270 135.290 109.320 ;
        RECT 131.210 108.990 135.290 109.270 ;
        RECT 131.210 108.940 131.590 108.990 ;
        RECT 134.910 108.940 135.290 108.990 ;
        RECT 6.700 107.615 9.560 107.995 ;
        RECT 39.150 107.615 42.010 107.995 ;
        RECT 71.600 107.615 74.460 107.995 ;
        RECT 104.050 107.615 106.910 107.995 ;
        RECT 137.355 107.955 137.735 108.335 ;
        RECT 139.395 107.955 139.775 108.335 ;
        RECT 141.180 107.955 141.560 108.335 ;
        RECT 6.700 106.855 9.560 107.235 ;
        RECT 39.150 106.855 42.010 107.235 ;
        RECT 71.600 106.855 74.460 107.235 ;
        RECT 104.050 106.855 106.910 107.235 ;
        RECT 0.240 106.455 0.620 106.835 ;
        RECT 4.160 106.455 4.540 106.835 ;
        RECT 35.140 106.625 35.520 106.675 ;
        RECT 37.560 106.625 37.940 106.675 ;
        RECT 35.140 106.345 37.940 106.625 ;
        RECT 35.140 106.295 35.520 106.345 ;
        RECT 37.560 106.295 37.940 106.345 ;
        RECT 67.590 106.625 67.970 106.675 ;
        RECT 70.010 106.625 70.390 106.675 ;
        RECT 67.590 106.345 70.390 106.625 ;
        RECT 67.590 106.295 67.970 106.345 ;
        RECT 70.010 106.295 70.390 106.345 ;
        RECT 100.040 106.625 100.420 106.675 ;
        RECT 102.460 106.625 102.840 106.675 ;
        RECT 100.040 106.345 102.840 106.625 ;
        RECT 100.040 106.295 100.420 106.345 ;
        RECT 102.460 106.295 102.840 106.345 ;
        RECT 132.490 106.625 132.870 106.675 ;
        RECT 134.910 106.625 135.290 106.675 ;
        RECT 132.490 106.345 135.290 106.625 ;
        RECT 132.490 106.295 132.870 106.345 ;
        RECT 134.910 106.295 135.290 106.345 ;
        RECT 6.700 105.015 9.560 105.395 ;
        RECT 39.150 105.015 42.010 105.395 ;
        RECT 71.600 105.015 74.460 105.395 ;
        RECT 104.050 105.015 106.910 105.395 ;
        RECT 137.355 104.955 137.735 105.335 ;
        RECT 139.395 104.955 139.775 105.335 ;
        RECT 141.180 104.955 141.560 105.335 ;
        RECT 36.420 104.785 36.800 104.835 ;
        RECT 37.560 104.785 37.940 104.835 ;
        RECT 36.420 104.505 37.940 104.785 ;
        RECT 36.420 104.455 36.800 104.505 ;
        RECT 37.560 104.455 37.940 104.505 ;
        RECT 68.870 104.785 69.250 104.835 ;
        RECT 70.010 104.785 70.390 104.835 ;
        RECT 68.870 104.505 70.390 104.785 ;
        RECT 68.870 104.455 69.250 104.505 ;
        RECT 70.010 104.455 70.390 104.505 ;
        RECT 101.320 104.785 101.700 104.835 ;
        RECT 102.460 104.785 102.840 104.835 ;
        RECT 101.320 104.505 102.840 104.785 ;
        RECT 101.320 104.455 101.700 104.505 ;
        RECT 102.460 104.455 102.840 104.505 ;
        RECT 133.770 104.785 134.150 104.835 ;
        RECT 134.910 104.785 135.290 104.835 ;
        RECT 133.770 104.505 135.290 104.785 ;
        RECT 133.770 104.455 134.150 104.505 ;
        RECT 134.910 104.455 135.290 104.505 ;
        RECT 0.240 103.455 0.620 103.835 ;
        RECT 4.160 103.455 4.540 103.835 ;
        RECT 6.700 103.175 9.560 103.555 ;
        RECT 39.150 103.175 42.010 103.555 ;
        RECT 71.600 103.175 74.460 103.555 ;
        RECT 104.050 103.175 106.910 103.555 ;
        RECT 37.560 102.615 38.080 102.995 ;
        RECT 70.010 102.615 70.530 102.995 ;
        RECT 102.460 102.615 102.980 102.995 ;
        RECT 134.910 102.615 135.430 102.995 ;
        RECT 137.355 101.955 137.735 102.335 ;
        RECT 139.395 101.955 139.775 102.335 ;
        RECT 141.180 101.955 141.560 102.335 ;
        RECT 0.240 100.455 0.620 100.835 ;
        RECT 4.160 100.455 4.540 100.835 ;
        RECT 0.240 97.455 0.620 97.835 ;
        RECT 137.355 95.955 137.735 96.335 ;
        RECT 139.395 95.955 139.775 96.335 ;
        RECT 141.180 95.955 141.560 96.335 ;
        RECT 0.240 94.455 0.620 94.835 ;
        RECT 4.160 94.455 4.540 94.835 ;
        RECT 37.060 94.050 37.940 94.430 ;
        RECT 69.510 94.050 70.390 94.430 ;
        RECT 101.960 94.050 102.840 94.430 ;
        RECT 134.410 94.050 135.290 94.430 ;
        RECT 6.700 93.490 9.560 93.870 ;
        RECT 39.150 93.490 42.010 93.870 ;
        RECT 71.600 93.490 74.460 93.870 ;
        RECT 104.050 93.490 106.910 93.870 ;
        RECT 137.355 92.955 137.735 93.335 ;
        RECT 139.395 92.955 139.775 93.335 ;
        RECT 141.180 92.955 141.560 93.335 ;
        RECT 35.780 92.540 36.160 92.590 ;
        RECT 37.560 92.540 37.940 92.590 ;
        RECT 35.780 92.260 37.940 92.540 ;
        RECT 35.780 92.210 36.160 92.260 ;
        RECT 37.560 92.210 37.940 92.260 ;
        RECT 68.230 92.540 68.610 92.590 ;
        RECT 70.010 92.540 70.390 92.590 ;
        RECT 68.230 92.260 70.390 92.540 ;
        RECT 68.230 92.210 68.610 92.260 ;
        RECT 70.010 92.210 70.390 92.260 ;
        RECT 100.680 92.540 101.060 92.590 ;
        RECT 102.460 92.540 102.840 92.590 ;
        RECT 100.680 92.260 102.840 92.540 ;
        RECT 100.680 92.210 101.060 92.260 ;
        RECT 102.460 92.210 102.840 92.260 ;
        RECT 133.130 92.540 133.510 92.590 ;
        RECT 134.910 92.540 135.290 92.590 ;
        RECT 133.130 92.260 135.290 92.540 ;
        RECT 133.130 92.210 133.510 92.260 ;
        RECT 134.910 92.210 135.290 92.260 ;
        RECT 0.240 91.455 0.620 91.835 ;
        RECT 4.160 91.455 4.540 91.835 ;
        RECT 6.700 91.650 9.560 92.030 ;
        RECT 39.150 91.650 42.010 92.030 ;
        RECT 71.600 91.650 74.460 92.030 ;
        RECT 104.050 91.650 106.910 92.030 ;
        RECT 34.500 90.695 34.880 90.745 ;
        RECT 37.560 90.695 37.940 90.745 ;
        RECT 34.500 90.415 37.940 90.695 ;
        RECT 34.500 90.365 34.880 90.415 ;
        RECT 37.560 90.365 37.940 90.415 ;
        RECT 66.950 90.695 67.330 90.745 ;
        RECT 70.010 90.695 70.390 90.745 ;
        RECT 66.950 90.415 70.390 90.695 ;
        RECT 66.950 90.365 67.330 90.415 ;
        RECT 70.010 90.365 70.390 90.415 ;
        RECT 99.400 90.695 99.780 90.745 ;
        RECT 102.460 90.695 102.840 90.745 ;
        RECT 99.400 90.415 102.840 90.695 ;
        RECT 99.400 90.365 99.780 90.415 ;
        RECT 102.460 90.365 102.840 90.415 ;
        RECT 131.850 90.695 132.230 90.745 ;
        RECT 134.910 90.695 135.290 90.745 ;
        RECT 131.850 90.415 135.290 90.695 ;
        RECT 131.850 90.365 132.230 90.415 ;
        RECT 134.910 90.365 135.290 90.415 ;
        RECT 6.700 89.805 9.560 90.185 ;
        RECT 39.150 89.805 42.010 90.185 ;
        RECT 71.600 89.805 74.460 90.185 ;
        RECT 104.050 89.805 106.910 90.185 ;
        RECT 137.355 89.955 137.735 90.335 ;
        RECT 139.395 89.955 139.775 90.335 ;
        RECT 141.180 89.955 141.560 90.335 ;
        RECT 6.700 89.045 9.560 89.425 ;
        RECT 39.150 89.045 42.010 89.425 ;
        RECT 71.600 89.045 74.460 89.425 ;
        RECT 104.050 89.045 106.910 89.425 ;
        RECT 0.240 88.455 0.620 88.835 ;
        RECT 4.160 88.455 4.540 88.835 ;
        RECT 33.220 88.055 33.600 88.105 ;
        RECT 37.560 88.055 37.940 88.105 ;
        RECT 33.220 87.775 37.940 88.055 ;
        RECT 33.220 87.725 33.600 87.775 ;
        RECT 37.560 87.725 37.940 87.775 ;
        RECT 65.670 88.055 66.050 88.105 ;
        RECT 70.010 88.055 70.390 88.105 ;
        RECT 65.670 87.775 70.390 88.055 ;
        RECT 65.670 87.725 66.050 87.775 ;
        RECT 70.010 87.725 70.390 87.775 ;
        RECT 98.120 88.055 98.500 88.105 ;
        RECT 102.460 88.055 102.840 88.105 ;
        RECT 98.120 87.775 102.840 88.055 ;
        RECT 98.120 87.725 98.500 87.775 ;
        RECT 102.460 87.725 102.840 87.775 ;
        RECT 130.570 88.055 130.950 88.105 ;
        RECT 134.910 88.055 135.290 88.105 ;
        RECT 130.570 87.775 135.290 88.055 ;
        RECT 130.570 87.725 130.950 87.775 ;
        RECT 134.910 87.725 135.290 87.775 ;
        RECT 6.700 87.165 9.560 87.545 ;
        RECT 39.150 87.165 42.010 87.545 ;
        RECT 71.600 87.165 74.460 87.545 ;
        RECT 104.050 87.165 106.910 87.545 ;
        RECT 137.355 86.955 137.735 87.335 ;
        RECT 139.395 86.955 139.775 87.335 ;
        RECT 141.180 86.955 141.560 87.335 ;
        RECT 31.940 86.215 32.320 86.265 ;
        RECT 37.560 86.215 37.940 86.265 ;
        RECT 31.940 85.935 37.940 86.215 ;
        RECT 31.940 85.885 32.320 85.935 ;
        RECT 37.560 85.885 37.940 85.935 ;
        RECT 64.390 86.215 64.770 86.265 ;
        RECT 70.010 86.215 70.390 86.265 ;
        RECT 64.390 85.935 70.390 86.215 ;
        RECT 64.390 85.885 64.770 85.935 ;
        RECT 70.010 85.885 70.390 85.935 ;
        RECT 96.840 86.215 97.220 86.265 ;
        RECT 102.460 86.215 102.840 86.265 ;
        RECT 96.840 85.935 102.840 86.215 ;
        RECT 96.840 85.885 97.220 85.935 ;
        RECT 102.460 85.885 102.840 85.935 ;
        RECT 129.290 86.215 129.670 86.265 ;
        RECT 134.910 86.215 135.290 86.265 ;
        RECT 129.290 85.935 135.290 86.215 ;
        RECT 129.290 85.885 129.670 85.935 ;
        RECT 134.910 85.885 135.290 85.935 ;
        RECT 0.240 85.455 0.620 85.835 ;
        RECT 4.160 85.455 4.540 85.835 ;
        RECT 6.700 85.325 9.560 85.705 ;
        RECT 39.150 85.325 42.010 85.705 ;
        RECT 71.600 85.325 74.460 85.705 ;
        RECT 104.050 85.325 106.910 85.705 ;
        RECT 30.660 84.370 31.040 84.420 ;
        RECT 37.560 84.370 37.940 84.420 ;
        RECT 30.660 84.090 37.940 84.370 ;
        RECT 30.660 84.040 31.040 84.090 ;
        RECT 37.560 84.040 37.940 84.090 ;
        RECT 63.110 84.370 63.490 84.420 ;
        RECT 70.010 84.370 70.390 84.420 ;
        RECT 63.110 84.090 70.390 84.370 ;
        RECT 63.110 84.040 63.490 84.090 ;
        RECT 70.010 84.040 70.390 84.090 ;
        RECT 95.560 84.370 95.940 84.420 ;
        RECT 102.460 84.370 102.840 84.420 ;
        RECT 95.560 84.090 102.840 84.370 ;
        RECT 95.560 84.040 95.940 84.090 ;
        RECT 102.460 84.040 102.840 84.090 ;
        RECT 128.010 84.370 128.390 84.420 ;
        RECT 134.910 84.370 135.290 84.420 ;
        RECT 128.010 84.090 135.290 84.370 ;
        RECT 128.010 84.040 128.390 84.090 ;
        RECT 134.910 84.040 135.290 84.090 ;
        RECT 137.355 83.955 137.735 84.335 ;
        RECT 139.395 83.955 139.775 84.335 ;
        RECT 141.180 83.955 141.560 84.335 ;
        RECT 6.700 83.480 9.560 83.860 ;
        RECT 39.150 83.480 42.010 83.860 ;
        RECT 71.600 83.480 74.460 83.860 ;
        RECT 104.050 83.480 106.910 83.860 ;
        RECT 0.240 82.455 0.620 82.835 ;
        RECT 4.160 82.455 4.540 82.835 ;
        RECT 6.700 82.720 9.560 83.100 ;
        RECT 39.150 82.720 42.010 83.100 ;
        RECT 71.600 82.720 74.460 83.100 ;
        RECT 104.050 82.720 106.910 83.100 ;
        RECT 29.380 81.730 29.760 81.780 ;
        RECT 37.560 81.730 37.940 81.780 ;
        RECT 29.380 81.450 37.940 81.730 ;
        RECT 29.380 81.400 29.760 81.450 ;
        RECT 37.560 81.400 37.940 81.450 ;
        RECT 61.830 81.730 62.210 81.780 ;
        RECT 70.010 81.730 70.390 81.780 ;
        RECT 61.830 81.450 70.390 81.730 ;
        RECT 61.830 81.400 62.210 81.450 ;
        RECT 70.010 81.400 70.390 81.450 ;
        RECT 94.280 81.730 94.660 81.780 ;
        RECT 102.460 81.730 102.840 81.780 ;
        RECT 94.280 81.450 102.840 81.730 ;
        RECT 94.280 81.400 94.660 81.450 ;
        RECT 102.460 81.400 102.840 81.450 ;
        RECT 126.730 81.730 127.110 81.780 ;
        RECT 134.910 81.730 135.290 81.780 ;
        RECT 126.730 81.450 135.290 81.730 ;
        RECT 126.730 81.400 127.110 81.450 ;
        RECT 134.910 81.400 135.290 81.450 ;
        RECT 6.700 80.840 9.560 81.220 ;
        RECT 39.150 80.840 42.010 81.220 ;
        RECT 71.600 80.840 74.460 81.220 ;
        RECT 104.050 80.840 106.910 81.220 ;
        RECT 137.355 80.955 137.735 81.335 ;
        RECT 139.395 80.955 139.775 81.335 ;
        RECT 141.180 80.955 141.560 81.335 ;
        RECT 28.100 79.890 28.480 79.940 ;
        RECT 37.560 79.890 37.940 79.940 ;
        RECT 0.240 79.455 0.620 79.835 ;
        RECT 4.160 79.455 4.540 79.835 ;
        RECT 28.100 79.610 37.940 79.890 ;
        RECT 28.100 79.560 28.480 79.610 ;
        RECT 37.560 79.560 37.940 79.610 ;
        RECT 60.550 79.890 60.930 79.940 ;
        RECT 70.010 79.890 70.390 79.940 ;
        RECT 60.550 79.610 70.390 79.890 ;
        RECT 60.550 79.560 60.930 79.610 ;
        RECT 70.010 79.560 70.390 79.610 ;
        RECT 93.000 79.890 93.380 79.940 ;
        RECT 102.460 79.890 102.840 79.940 ;
        RECT 93.000 79.610 102.840 79.890 ;
        RECT 93.000 79.560 93.380 79.610 ;
        RECT 102.460 79.560 102.840 79.610 ;
        RECT 125.450 79.890 125.830 79.940 ;
        RECT 134.910 79.890 135.290 79.940 ;
        RECT 125.450 79.610 135.290 79.890 ;
        RECT 125.450 79.560 125.830 79.610 ;
        RECT 134.910 79.560 135.290 79.610 ;
        RECT 6.700 79.000 9.560 79.380 ;
        RECT 39.150 79.000 42.010 79.380 ;
        RECT 71.600 79.000 74.460 79.380 ;
        RECT 104.050 79.000 106.910 79.380 ;
        RECT 6.700 78.280 9.560 78.660 ;
        RECT 39.150 78.280 42.010 78.660 ;
        RECT 71.600 78.280 74.460 78.660 ;
        RECT 104.050 78.280 106.910 78.660 ;
        RECT 28.740 78.050 29.120 78.100 ;
        RECT 37.560 78.050 37.940 78.100 ;
        RECT 28.740 77.770 37.940 78.050 ;
        RECT 28.740 77.720 29.120 77.770 ;
        RECT 37.560 77.720 37.940 77.770 ;
        RECT 61.190 78.050 61.570 78.100 ;
        RECT 70.010 78.050 70.390 78.100 ;
        RECT 61.190 77.770 70.390 78.050 ;
        RECT 61.190 77.720 61.570 77.770 ;
        RECT 70.010 77.720 70.390 77.770 ;
        RECT 93.640 78.050 94.020 78.100 ;
        RECT 102.460 78.050 102.840 78.100 ;
        RECT 93.640 77.770 102.840 78.050 ;
        RECT 93.640 77.720 94.020 77.770 ;
        RECT 102.460 77.720 102.840 77.770 ;
        RECT 126.090 78.050 126.470 78.100 ;
        RECT 134.910 78.050 135.290 78.100 ;
        RECT 126.090 77.770 135.290 78.050 ;
        RECT 126.090 77.720 126.470 77.770 ;
        RECT 134.910 77.720 135.290 77.770 ;
        RECT 0.240 76.070 0.620 76.450 ;
        RECT 4.160 76.070 4.540 76.450 ;
        RECT 6.700 76.440 9.560 76.820 ;
        RECT 39.150 76.440 42.010 76.820 ;
        RECT 71.600 76.440 74.460 76.820 ;
        RECT 104.050 76.440 106.910 76.820 ;
        RECT 30.020 76.210 30.400 76.260 ;
        RECT 37.560 76.210 37.940 76.260 ;
        RECT 30.020 75.930 37.940 76.210 ;
        RECT 30.020 75.880 30.400 75.930 ;
        RECT 37.560 75.880 37.940 75.930 ;
        RECT 62.470 76.210 62.850 76.260 ;
        RECT 70.010 76.210 70.390 76.260 ;
        RECT 62.470 75.930 70.390 76.210 ;
        RECT 62.470 75.880 62.850 75.930 ;
        RECT 70.010 75.880 70.390 75.930 ;
        RECT 94.920 76.210 95.300 76.260 ;
        RECT 102.460 76.210 102.840 76.260 ;
        RECT 94.920 75.930 102.840 76.210 ;
        RECT 94.920 75.880 95.300 75.930 ;
        RECT 102.460 75.880 102.840 75.930 ;
        RECT 127.370 76.210 127.750 76.260 ;
        RECT 134.910 76.210 135.290 76.260 ;
        RECT 127.370 75.930 135.290 76.210 ;
        RECT 127.370 75.880 127.750 75.930 ;
        RECT 134.910 75.880 135.290 75.930 ;
        RECT 6.700 74.555 9.560 74.935 ;
        RECT 39.150 74.555 42.010 74.935 ;
        RECT 71.600 74.555 74.460 74.935 ;
        RECT 104.050 74.555 106.910 74.935 ;
        RECT 137.355 74.570 137.735 74.950 ;
        RECT 139.395 74.570 139.775 74.950 ;
        RECT 141.180 74.570 141.560 74.950 ;
        RECT 6.700 73.795 9.560 74.175 ;
        RECT 39.150 73.795 42.010 74.175 ;
        RECT 71.600 73.795 74.460 74.175 ;
        RECT 104.050 73.795 106.910 74.175 ;
        RECT 31.300 73.565 31.680 73.615 ;
        RECT 37.560 73.565 37.940 73.615 ;
        RECT 0.240 73.070 0.620 73.450 ;
        RECT 4.160 73.070 4.540 73.450 ;
        RECT 31.300 73.285 37.940 73.565 ;
        RECT 31.300 73.235 31.680 73.285 ;
        RECT 37.560 73.235 37.940 73.285 ;
        RECT 63.750 73.565 64.130 73.615 ;
        RECT 70.010 73.565 70.390 73.615 ;
        RECT 63.750 73.285 70.390 73.565 ;
        RECT 63.750 73.235 64.130 73.285 ;
        RECT 70.010 73.235 70.390 73.285 ;
        RECT 96.200 73.565 96.580 73.615 ;
        RECT 102.460 73.565 102.840 73.615 ;
        RECT 96.200 73.285 102.840 73.565 ;
        RECT 96.200 73.235 96.580 73.285 ;
        RECT 102.460 73.235 102.840 73.285 ;
        RECT 128.650 73.565 129.030 73.615 ;
        RECT 134.910 73.565 135.290 73.615 ;
        RECT 128.650 73.285 135.290 73.565 ;
        RECT 128.650 73.235 129.030 73.285 ;
        RECT 134.910 73.235 135.290 73.285 ;
        RECT 6.700 71.955 9.560 72.335 ;
        RECT 39.150 71.955 42.010 72.335 ;
        RECT 71.600 71.955 74.460 72.335 ;
        RECT 104.050 71.955 106.910 72.335 ;
        RECT 32.580 71.725 32.960 71.775 ;
        RECT 37.560 71.725 37.940 71.775 ;
        RECT 32.580 71.445 37.940 71.725 ;
        RECT 32.580 71.395 32.960 71.445 ;
        RECT 37.560 71.395 37.940 71.445 ;
        RECT 65.030 71.725 65.410 71.775 ;
        RECT 70.010 71.725 70.390 71.775 ;
        RECT 65.030 71.445 70.390 71.725 ;
        RECT 65.030 71.395 65.410 71.445 ;
        RECT 70.010 71.395 70.390 71.445 ;
        RECT 97.480 71.725 97.860 71.775 ;
        RECT 102.460 71.725 102.840 71.775 ;
        RECT 97.480 71.445 102.840 71.725 ;
        RECT 97.480 71.395 97.860 71.445 ;
        RECT 102.460 71.395 102.840 71.445 ;
        RECT 129.930 71.725 130.310 71.775 ;
        RECT 134.910 71.725 135.290 71.775 ;
        RECT 129.930 71.445 135.290 71.725 ;
        RECT 137.355 71.570 137.735 71.950 ;
        RECT 139.395 71.570 139.775 71.950 ;
        RECT 141.180 71.570 141.560 71.950 ;
        RECT 129.930 71.395 130.310 71.445 ;
        RECT 134.910 71.395 135.290 71.445 ;
        RECT 0.240 70.070 0.620 70.450 ;
        RECT 4.160 70.070 4.540 70.450 ;
        RECT 6.700 70.115 9.560 70.495 ;
        RECT 39.150 70.115 42.010 70.495 ;
        RECT 71.600 70.115 74.460 70.495 ;
        RECT 104.050 70.115 106.910 70.495 ;
        RECT 33.860 69.885 34.240 69.935 ;
        RECT 37.560 69.885 37.940 69.935 ;
        RECT 33.860 69.605 37.940 69.885 ;
        RECT 33.860 69.555 34.240 69.605 ;
        RECT 37.560 69.555 37.940 69.605 ;
        RECT 66.310 69.885 66.690 69.935 ;
        RECT 70.010 69.885 70.390 69.935 ;
        RECT 66.310 69.605 70.390 69.885 ;
        RECT 66.310 69.555 66.690 69.605 ;
        RECT 70.010 69.555 70.390 69.605 ;
        RECT 98.760 69.885 99.140 69.935 ;
        RECT 102.460 69.885 102.840 69.935 ;
        RECT 98.760 69.605 102.840 69.885 ;
        RECT 98.760 69.555 99.140 69.605 ;
        RECT 102.460 69.555 102.840 69.605 ;
        RECT 131.210 69.885 131.590 69.935 ;
        RECT 134.910 69.885 135.290 69.935 ;
        RECT 131.210 69.605 135.290 69.885 ;
        RECT 131.210 69.555 131.590 69.605 ;
        RECT 134.910 69.555 135.290 69.605 ;
        RECT 6.700 68.230 9.560 68.610 ;
        RECT 39.150 68.230 42.010 68.610 ;
        RECT 71.600 68.230 74.460 68.610 ;
        RECT 104.050 68.230 106.910 68.610 ;
        RECT 137.355 68.570 137.735 68.950 ;
        RECT 139.395 68.570 139.775 68.950 ;
        RECT 141.180 68.570 141.560 68.950 ;
        RECT 6.700 67.470 9.560 67.850 ;
        RECT 39.150 67.470 42.010 67.850 ;
        RECT 71.600 67.470 74.460 67.850 ;
        RECT 104.050 67.470 106.910 67.850 ;
        RECT 0.240 67.070 0.620 67.450 ;
        RECT 4.160 67.070 4.540 67.450 ;
        RECT 35.140 67.240 35.520 67.290 ;
        RECT 37.560 67.240 37.940 67.290 ;
        RECT 35.140 66.960 37.940 67.240 ;
        RECT 35.140 66.910 35.520 66.960 ;
        RECT 37.560 66.910 37.940 66.960 ;
        RECT 67.590 67.240 67.970 67.290 ;
        RECT 70.010 67.240 70.390 67.290 ;
        RECT 67.590 66.960 70.390 67.240 ;
        RECT 67.590 66.910 67.970 66.960 ;
        RECT 70.010 66.910 70.390 66.960 ;
        RECT 100.040 67.240 100.420 67.290 ;
        RECT 102.460 67.240 102.840 67.290 ;
        RECT 100.040 66.960 102.840 67.240 ;
        RECT 100.040 66.910 100.420 66.960 ;
        RECT 102.460 66.910 102.840 66.960 ;
        RECT 132.490 67.240 132.870 67.290 ;
        RECT 134.910 67.240 135.290 67.290 ;
        RECT 132.490 66.960 135.290 67.240 ;
        RECT 132.490 66.910 132.870 66.960 ;
        RECT 134.910 66.910 135.290 66.960 ;
        RECT 6.700 65.630 9.560 66.010 ;
        RECT 39.150 65.630 42.010 66.010 ;
        RECT 71.600 65.630 74.460 66.010 ;
        RECT 104.050 65.630 106.910 66.010 ;
        RECT 137.355 65.570 137.735 65.950 ;
        RECT 139.395 65.570 139.775 65.950 ;
        RECT 141.180 65.570 141.560 65.950 ;
        RECT 36.420 65.400 36.800 65.450 ;
        RECT 37.560 65.400 37.940 65.450 ;
        RECT 36.420 65.120 37.940 65.400 ;
        RECT 36.420 65.070 36.800 65.120 ;
        RECT 37.560 65.070 37.940 65.120 ;
        RECT 68.870 65.400 69.250 65.450 ;
        RECT 70.010 65.400 70.390 65.450 ;
        RECT 68.870 65.120 70.390 65.400 ;
        RECT 68.870 65.070 69.250 65.120 ;
        RECT 70.010 65.070 70.390 65.120 ;
        RECT 101.320 65.400 101.700 65.450 ;
        RECT 102.460 65.400 102.840 65.450 ;
        RECT 101.320 65.120 102.840 65.400 ;
        RECT 101.320 65.070 101.700 65.120 ;
        RECT 102.460 65.070 102.840 65.120 ;
        RECT 133.770 65.400 134.150 65.450 ;
        RECT 134.910 65.400 135.290 65.450 ;
        RECT 133.770 65.120 135.290 65.400 ;
        RECT 133.770 65.070 134.150 65.120 ;
        RECT 134.910 65.070 135.290 65.120 ;
        RECT 0.240 64.070 0.620 64.450 ;
        RECT 4.160 64.070 4.540 64.450 ;
        RECT 6.700 63.790 9.560 64.170 ;
        RECT 39.150 63.790 42.010 64.170 ;
        RECT 71.600 63.790 74.460 64.170 ;
        RECT 104.050 63.790 106.910 64.170 ;
        RECT 37.560 63.230 38.080 63.610 ;
        RECT 70.010 63.230 70.530 63.610 ;
        RECT 102.460 63.230 102.980 63.610 ;
        RECT 134.910 63.230 135.430 63.610 ;
        RECT 137.355 62.570 137.735 62.950 ;
        RECT 139.395 62.570 139.775 62.950 ;
        RECT 141.180 62.570 141.560 62.950 ;
        RECT 0.240 61.070 0.620 61.450 ;
        RECT 4.160 61.070 4.540 61.450 ;
        RECT 0.240 58.070 0.620 58.450 ;
        RECT 137.355 56.570 137.735 56.950 ;
        RECT 139.395 56.570 139.775 56.950 ;
        RECT 141.180 56.570 141.560 56.950 ;
        RECT 0.240 55.070 0.620 55.450 ;
        RECT 4.160 55.070 4.540 55.450 ;
        RECT 37.060 54.665 37.940 55.045 ;
        RECT 69.510 54.665 70.390 55.045 ;
        RECT 101.960 54.665 102.840 55.045 ;
        RECT 134.410 54.665 135.290 55.045 ;
        RECT 6.700 54.105 9.560 54.485 ;
        RECT 39.150 54.105 42.010 54.485 ;
        RECT 71.600 54.105 74.460 54.485 ;
        RECT 104.050 54.105 106.910 54.485 ;
        RECT 137.355 53.570 137.735 53.950 ;
        RECT 139.395 53.570 139.775 53.950 ;
        RECT 141.180 53.570 141.560 53.950 ;
        RECT 35.780 53.155 36.160 53.205 ;
        RECT 37.560 53.155 37.940 53.205 ;
        RECT 35.780 52.875 37.940 53.155 ;
        RECT 35.780 52.825 36.160 52.875 ;
        RECT 37.560 52.825 37.940 52.875 ;
        RECT 68.230 53.155 68.610 53.205 ;
        RECT 70.010 53.155 70.390 53.205 ;
        RECT 68.230 52.875 70.390 53.155 ;
        RECT 68.230 52.825 68.610 52.875 ;
        RECT 70.010 52.825 70.390 52.875 ;
        RECT 100.680 53.155 101.060 53.205 ;
        RECT 102.460 53.155 102.840 53.205 ;
        RECT 100.680 52.875 102.840 53.155 ;
        RECT 100.680 52.825 101.060 52.875 ;
        RECT 102.460 52.825 102.840 52.875 ;
        RECT 133.130 53.155 133.510 53.205 ;
        RECT 134.910 53.155 135.290 53.205 ;
        RECT 133.130 52.875 135.290 53.155 ;
        RECT 133.130 52.825 133.510 52.875 ;
        RECT 134.910 52.825 135.290 52.875 ;
        RECT 0.240 52.070 0.620 52.450 ;
        RECT 4.160 52.070 4.540 52.450 ;
        RECT 6.700 52.265 9.560 52.645 ;
        RECT 39.150 52.265 42.010 52.645 ;
        RECT 71.600 52.265 74.460 52.645 ;
        RECT 104.050 52.265 106.910 52.645 ;
        RECT 34.500 51.310 34.880 51.360 ;
        RECT 37.560 51.310 37.940 51.360 ;
        RECT 34.500 51.030 37.940 51.310 ;
        RECT 34.500 50.980 34.880 51.030 ;
        RECT 37.560 50.980 37.940 51.030 ;
        RECT 66.950 51.310 67.330 51.360 ;
        RECT 70.010 51.310 70.390 51.360 ;
        RECT 66.950 51.030 70.390 51.310 ;
        RECT 66.950 50.980 67.330 51.030 ;
        RECT 70.010 50.980 70.390 51.030 ;
        RECT 99.400 51.310 99.780 51.360 ;
        RECT 102.460 51.310 102.840 51.360 ;
        RECT 99.400 51.030 102.840 51.310 ;
        RECT 99.400 50.980 99.780 51.030 ;
        RECT 102.460 50.980 102.840 51.030 ;
        RECT 131.850 51.310 132.230 51.360 ;
        RECT 134.910 51.310 135.290 51.360 ;
        RECT 131.850 51.030 135.290 51.310 ;
        RECT 131.850 50.980 132.230 51.030 ;
        RECT 134.910 50.980 135.290 51.030 ;
        RECT 6.700 50.420 9.560 50.800 ;
        RECT 39.150 50.420 42.010 50.800 ;
        RECT 71.600 50.420 74.460 50.800 ;
        RECT 104.050 50.420 106.910 50.800 ;
        RECT 137.355 50.570 137.735 50.950 ;
        RECT 139.395 50.570 139.775 50.950 ;
        RECT 141.180 50.570 141.560 50.950 ;
        RECT 6.700 49.660 9.560 50.040 ;
        RECT 39.150 49.660 42.010 50.040 ;
        RECT 71.600 49.660 74.460 50.040 ;
        RECT 104.050 49.660 106.910 50.040 ;
        RECT 0.240 49.070 0.620 49.450 ;
        RECT 4.160 49.070 4.540 49.450 ;
        RECT 33.220 48.670 33.600 48.720 ;
        RECT 37.560 48.670 37.940 48.720 ;
        RECT 33.220 48.390 37.940 48.670 ;
        RECT 33.220 48.340 33.600 48.390 ;
        RECT 37.560 48.340 37.940 48.390 ;
        RECT 65.670 48.670 66.050 48.720 ;
        RECT 70.010 48.670 70.390 48.720 ;
        RECT 65.670 48.390 70.390 48.670 ;
        RECT 65.670 48.340 66.050 48.390 ;
        RECT 70.010 48.340 70.390 48.390 ;
        RECT 98.120 48.670 98.500 48.720 ;
        RECT 102.460 48.670 102.840 48.720 ;
        RECT 98.120 48.390 102.840 48.670 ;
        RECT 98.120 48.340 98.500 48.390 ;
        RECT 102.460 48.340 102.840 48.390 ;
        RECT 130.570 48.670 130.950 48.720 ;
        RECT 134.910 48.670 135.290 48.720 ;
        RECT 130.570 48.390 135.290 48.670 ;
        RECT 130.570 48.340 130.950 48.390 ;
        RECT 134.910 48.340 135.290 48.390 ;
        RECT 6.700 47.780 9.560 48.160 ;
        RECT 39.150 47.780 42.010 48.160 ;
        RECT 71.600 47.780 74.460 48.160 ;
        RECT 104.050 47.780 106.910 48.160 ;
        RECT 137.355 47.570 137.735 47.950 ;
        RECT 139.395 47.570 139.775 47.950 ;
        RECT 141.180 47.570 141.560 47.950 ;
        RECT 31.940 46.830 32.320 46.880 ;
        RECT 37.560 46.830 37.940 46.880 ;
        RECT 31.940 46.550 37.940 46.830 ;
        RECT 31.940 46.500 32.320 46.550 ;
        RECT 37.560 46.500 37.940 46.550 ;
        RECT 64.390 46.830 64.770 46.880 ;
        RECT 70.010 46.830 70.390 46.880 ;
        RECT 64.390 46.550 70.390 46.830 ;
        RECT 64.390 46.500 64.770 46.550 ;
        RECT 70.010 46.500 70.390 46.550 ;
        RECT 96.840 46.830 97.220 46.880 ;
        RECT 102.460 46.830 102.840 46.880 ;
        RECT 96.840 46.550 102.840 46.830 ;
        RECT 96.840 46.500 97.220 46.550 ;
        RECT 102.460 46.500 102.840 46.550 ;
        RECT 129.290 46.830 129.670 46.880 ;
        RECT 134.910 46.830 135.290 46.880 ;
        RECT 129.290 46.550 135.290 46.830 ;
        RECT 129.290 46.500 129.670 46.550 ;
        RECT 134.910 46.500 135.290 46.550 ;
        RECT 0.240 46.070 0.620 46.450 ;
        RECT 4.160 46.070 4.540 46.450 ;
        RECT 6.700 45.940 9.560 46.320 ;
        RECT 39.150 45.940 42.010 46.320 ;
        RECT 71.600 45.940 74.460 46.320 ;
        RECT 104.050 45.940 106.910 46.320 ;
        RECT 30.660 44.985 31.040 45.035 ;
        RECT 37.560 44.985 37.940 45.035 ;
        RECT 30.660 44.705 37.940 44.985 ;
        RECT 30.660 44.655 31.040 44.705 ;
        RECT 37.560 44.655 37.940 44.705 ;
        RECT 63.110 44.985 63.490 45.035 ;
        RECT 70.010 44.985 70.390 45.035 ;
        RECT 63.110 44.705 70.390 44.985 ;
        RECT 63.110 44.655 63.490 44.705 ;
        RECT 70.010 44.655 70.390 44.705 ;
        RECT 95.560 44.985 95.940 45.035 ;
        RECT 102.460 44.985 102.840 45.035 ;
        RECT 95.560 44.705 102.840 44.985 ;
        RECT 95.560 44.655 95.940 44.705 ;
        RECT 102.460 44.655 102.840 44.705 ;
        RECT 128.010 44.985 128.390 45.035 ;
        RECT 134.910 44.985 135.290 45.035 ;
        RECT 128.010 44.705 135.290 44.985 ;
        RECT 128.010 44.655 128.390 44.705 ;
        RECT 134.910 44.655 135.290 44.705 ;
        RECT 137.355 44.570 137.735 44.950 ;
        RECT 139.395 44.570 139.775 44.950 ;
        RECT 141.180 44.570 141.560 44.950 ;
        RECT 6.700 44.095 9.560 44.475 ;
        RECT 39.150 44.095 42.010 44.475 ;
        RECT 71.600 44.095 74.460 44.475 ;
        RECT 104.050 44.095 106.910 44.475 ;
        RECT 0.240 43.070 0.620 43.450 ;
        RECT 4.160 43.070 4.540 43.450 ;
        RECT 6.700 43.335 9.560 43.715 ;
        RECT 39.150 43.335 42.010 43.715 ;
        RECT 71.600 43.335 74.460 43.715 ;
        RECT 104.050 43.335 106.910 43.715 ;
        RECT 29.380 42.345 29.760 42.395 ;
        RECT 37.560 42.345 37.940 42.395 ;
        RECT 29.380 42.065 37.940 42.345 ;
        RECT 29.380 42.015 29.760 42.065 ;
        RECT 37.560 42.015 37.940 42.065 ;
        RECT 61.830 42.345 62.210 42.395 ;
        RECT 70.010 42.345 70.390 42.395 ;
        RECT 61.830 42.065 70.390 42.345 ;
        RECT 61.830 42.015 62.210 42.065 ;
        RECT 70.010 42.015 70.390 42.065 ;
        RECT 94.280 42.345 94.660 42.395 ;
        RECT 102.460 42.345 102.840 42.395 ;
        RECT 94.280 42.065 102.840 42.345 ;
        RECT 94.280 42.015 94.660 42.065 ;
        RECT 102.460 42.015 102.840 42.065 ;
        RECT 126.730 42.345 127.110 42.395 ;
        RECT 134.910 42.345 135.290 42.395 ;
        RECT 126.730 42.065 135.290 42.345 ;
        RECT 126.730 42.015 127.110 42.065 ;
        RECT 134.910 42.015 135.290 42.065 ;
        RECT 6.700 41.455 9.560 41.835 ;
        RECT 39.150 41.455 42.010 41.835 ;
        RECT 71.600 41.455 74.460 41.835 ;
        RECT 104.050 41.455 106.910 41.835 ;
        RECT 137.355 41.570 137.735 41.950 ;
        RECT 139.395 41.570 139.775 41.950 ;
        RECT 141.180 41.570 141.560 41.950 ;
        RECT 28.100 40.505 28.480 40.555 ;
        RECT 37.560 40.505 37.940 40.555 ;
        RECT 0.240 40.070 0.620 40.450 ;
        RECT 4.160 40.070 4.540 40.450 ;
        RECT 28.100 40.225 37.940 40.505 ;
        RECT 28.100 40.175 28.480 40.225 ;
        RECT 37.560 40.175 37.940 40.225 ;
        RECT 60.550 40.505 60.930 40.555 ;
        RECT 70.010 40.505 70.390 40.555 ;
        RECT 60.550 40.225 70.390 40.505 ;
        RECT 60.550 40.175 60.930 40.225 ;
        RECT 70.010 40.175 70.390 40.225 ;
        RECT 93.000 40.505 93.380 40.555 ;
        RECT 102.460 40.505 102.840 40.555 ;
        RECT 93.000 40.225 102.840 40.505 ;
        RECT 93.000 40.175 93.380 40.225 ;
        RECT 102.460 40.175 102.840 40.225 ;
        RECT 125.450 40.505 125.830 40.555 ;
        RECT 134.910 40.505 135.290 40.555 ;
        RECT 125.450 40.225 135.290 40.505 ;
        RECT 125.450 40.175 125.830 40.225 ;
        RECT 134.910 40.175 135.290 40.225 ;
        RECT 6.700 39.615 9.560 39.995 ;
        RECT 39.150 39.615 42.010 39.995 ;
        RECT 71.600 39.615 74.460 39.995 ;
        RECT 104.050 39.615 106.910 39.995 ;
        RECT 6.700 38.895 9.560 39.275 ;
        RECT 39.150 38.895 42.010 39.275 ;
        RECT 71.600 38.895 74.460 39.275 ;
        RECT 104.050 38.895 106.910 39.275 ;
        RECT 28.740 38.665 29.120 38.715 ;
        RECT 37.560 38.665 37.940 38.715 ;
        RECT 28.740 38.385 37.940 38.665 ;
        RECT 28.740 38.335 29.120 38.385 ;
        RECT 37.560 38.335 37.940 38.385 ;
        RECT 61.190 38.665 61.570 38.715 ;
        RECT 70.010 38.665 70.390 38.715 ;
        RECT 61.190 38.385 70.390 38.665 ;
        RECT 61.190 38.335 61.570 38.385 ;
        RECT 70.010 38.335 70.390 38.385 ;
        RECT 93.640 38.665 94.020 38.715 ;
        RECT 102.460 38.665 102.840 38.715 ;
        RECT 93.640 38.385 102.840 38.665 ;
        RECT 93.640 38.335 94.020 38.385 ;
        RECT 102.460 38.335 102.840 38.385 ;
        RECT 126.090 38.665 126.470 38.715 ;
        RECT 134.910 38.665 135.290 38.715 ;
        RECT 126.090 38.385 135.290 38.665 ;
        RECT 126.090 38.335 126.470 38.385 ;
        RECT 134.910 38.335 135.290 38.385 ;
        RECT 0.240 36.685 0.620 37.065 ;
        RECT 4.160 36.685 4.540 37.065 ;
        RECT 6.700 37.055 9.560 37.435 ;
        RECT 39.150 37.055 42.010 37.435 ;
        RECT 71.600 37.055 74.460 37.435 ;
        RECT 104.050 37.055 106.910 37.435 ;
        RECT 30.020 36.825 30.400 36.875 ;
        RECT 37.560 36.825 37.940 36.875 ;
        RECT 30.020 36.545 37.940 36.825 ;
        RECT 30.020 36.495 30.400 36.545 ;
        RECT 37.560 36.495 37.940 36.545 ;
        RECT 62.470 36.825 62.850 36.875 ;
        RECT 70.010 36.825 70.390 36.875 ;
        RECT 62.470 36.545 70.390 36.825 ;
        RECT 62.470 36.495 62.850 36.545 ;
        RECT 70.010 36.495 70.390 36.545 ;
        RECT 94.920 36.825 95.300 36.875 ;
        RECT 102.460 36.825 102.840 36.875 ;
        RECT 94.920 36.545 102.840 36.825 ;
        RECT 94.920 36.495 95.300 36.545 ;
        RECT 102.460 36.495 102.840 36.545 ;
        RECT 127.370 36.825 127.750 36.875 ;
        RECT 134.910 36.825 135.290 36.875 ;
        RECT 127.370 36.545 135.290 36.825 ;
        RECT 127.370 36.495 127.750 36.545 ;
        RECT 134.910 36.495 135.290 36.545 ;
        RECT 6.700 35.170 9.560 35.550 ;
        RECT 39.150 35.170 42.010 35.550 ;
        RECT 71.600 35.170 74.460 35.550 ;
        RECT 104.050 35.170 106.910 35.550 ;
        RECT 137.355 35.185 137.735 35.565 ;
        RECT 139.395 35.185 139.775 35.565 ;
        RECT 141.180 35.185 141.560 35.565 ;
        RECT 6.700 34.410 9.560 34.790 ;
        RECT 39.150 34.410 42.010 34.790 ;
        RECT 71.600 34.410 74.460 34.790 ;
        RECT 104.050 34.410 106.910 34.790 ;
        RECT 31.300 34.180 31.680 34.230 ;
        RECT 37.560 34.180 37.940 34.230 ;
        RECT 0.240 33.685 0.620 34.065 ;
        RECT 4.160 33.685 4.540 34.065 ;
        RECT 31.300 33.900 37.940 34.180 ;
        RECT 31.300 33.850 31.680 33.900 ;
        RECT 37.560 33.850 37.940 33.900 ;
        RECT 63.750 34.180 64.130 34.230 ;
        RECT 70.010 34.180 70.390 34.230 ;
        RECT 63.750 33.900 70.390 34.180 ;
        RECT 63.750 33.850 64.130 33.900 ;
        RECT 70.010 33.850 70.390 33.900 ;
        RECT 96.200 34.180 96.580 34.230 ;
        RECT 102.460 34.180 102.840 34.230 ;
        RECT 96.200 33.900 102.840 34.180 ;
        RECT 96.200 33.850 96.580 33.900 ;
        RECT 102.460 33.850 102.840 33.900 ;
        RECT 128.650 34.180 129.030 34.230 ;
        RECT 134.910 34.180 135.290 34.230 ;
        RECT 128.650 33.900 135.290 34.180 ;
        RECT 128.650 33.850 129.030 33.900 ;
        RECT 134.910 33.850 135.290 33.900 ;
        RECT 6.700 32.570 9.560 32.950 ;
        RECT 39.150 32.570 42.010 32.950 ;
        RECT 71.600 32.570 74.460 32.950 ;
        RECT 104.050 32.570 106.910 32.950 ;
        RECT 32.580 32.340 32.960 32.390 ;
        RECT 37.560 32.340 37.940 32.390 ;
        RECT 32.580 32.060 37.940 32.340 ;
        RECT 32.580 32.010 32.960 32.060 ;
        RECT 37.560 32.010 37.940 32.060 ;
        RECT 65.030 32.340 65.410 32.390 ;
        RECT 70.010 32.340 70.390 32.390 ;
        RECT 65.030 32.060 70.390 32.340 ;
        RECT 65.030 32.010 65.410 32.060 ;
        RECT 70.010 32.010 70.390 32.060 ;
        RECT 97.480 32.340 97.860 32.390 ;
        RECT 102.460 32.340 102.840 32.390 ;
        RECT 97.480 32.060 102.840 32.340 ;
        RECT 97.480 32.010 97.860 32.060 ;
        RECT 102.460 32.010 102.840 32.060 ;
        RECT 129.930 32.340 130.310 32.390 ;
        RECT 134.910 32.340 135.290 32.390 ;
        RECT 129.930 32.060 135.290 32.340 ;
        RECT 137.355 32.185 137.735 32.565 ;
        RECT 139.395 32.185 139.775 32.565 ;
        RECT 141.180 32.185 141.560 32.565 ;
        RECT 129.930 32.010 130.310 32.060 ;
        RECT 134.910 32.010 135.290 32.060 ;
        RECT 0.240 30.685 0.620 31.065 ;
        RECT 4.160 30.685 4.540 31.065 ;
        RECT 6.700 30.730 9.560 31.110 ;
        RECT 39.150 30.730 42.010 31.110 ;
        RECT 71.600 30.730 74.460 31.110 ;
        RECT 104.050 30.730 106.910 31.110 ;
        RECT 33.860 30.500 34.240 30.550 ;
        RECT 37.560 30.500 37.940 30.550 ;
        RECT 33.860 30.220 37.940 30.500 ;
        RECT 33.860 30.170 34.240 30.220 ;
        RECT 37.560 30.170 37.940 30.220 ;
        RECT 66.310 30.500 66.690 30.550 ;
        RECT 70.010 30.500 70.390 30.550 ;
        RECT 66.310 30.220 70.390 30.500 ;
        RECT 66.310 30.170 66.690 30.220 ;
        RECT 70.010 30.170 70.390 30.220 ;
        RECT 98.760 30.500 99.140 30.550 ;
        RECT 102.460 30.500 102.840 30.550 ;
        RECT 98.760 30.220 102.840 30.500 ;
        RECT 98.760 30.170 99.140 30.220 ;
        RECT 102.460 30.170 102.840 30.220 ;
        RECT 131.210 30.500 131.590 30.550 ;
        RECT 134.910 30.500 135.290 30.550 ;
        RECT 131.210 30.220 135.290 30.500 ;
        RECT 131.210 30.170 131.590 30.220 ;
        RECT 134.910 30.170 135.290 30.220 ;
        RECT 6.700 28.845 9.560 29.225 ;
        RECT 39.150 28.845 42.010 29.225 ;
        RECT 71.600 28.845 74.460 29.225 ;
        RECT 104.050 28.845 106.910 29.225 ;
        RECT 137.355 29.185 137.735 29.565 ;
        RECT 139.395 29.185 139.775 29.565 ;
        RECT 141.180 29.185 141.560 29.565 ;
        RECT 6.700 28.085 9.560 28.465 ;
        RECT 39.150 28.085 42.010 28.465 ;
        RECT 71.600 28.085 74.460 28.465 ;
        RECT 104.050 28.085 106.910 28.465 ;
        RECT 0.240 27.685 0.620 28.065 ;
        RECT 4.160 27.685 4.540 28.065 ;
        RECT 35.140 27.855 35.520 27.905 ;
        RECT 37.560 27.855 37.940 27.905 ;
        RECT 35.140 27.575 37.940 27.855 ;
        RECT 35.140 27.525 35.520 27.575 ;
        RECT 37.560 27.525 37.940 27.575 ;
        RECT 67.590 27.855 67.970 27.905 ;
        RECT 70.010 27.855 70.390 27.905 ;
        RECT 67.590 27.575 70.390 27.855 ;
        RECT 67.590 27.525 67.970 27.575 ;
        RECT 70.010 27.525 70.390 27.575 ;
        RECT 100.040 27.855 100.420 27.905 ;
        RECT 102.460 27.855 102.840 27.905 ;
        RECT 100.040 27.575 102.840 27.855 ;
        RECT 100.040 27.525 100.420 27.575 ;
        RECT 102.460 27.525 102.840 27.575 ;
        RECT 132.490 27.855 132.870 27.905 ;
        RECT 134.910 27.855 135.290 27.905 ;
        RECT 132.490 27.575 135.290 27.855 ;
        RECT 132.490 27.525 132.870 27.575 ;
        RECT 134.910 27.525 135.290 27.575 ;
        RECT 6.700 26.245 9.560 26.625 ;
        RECT 39.150 26.245 42.010 26.625 ;
        RECT 71.600 26.245 74.460 26.625 ;
        RECT 104.050 26.245 106.910 26.625 ;
        RECT 137.355 26.185 137.735 26.565 ;
        RECT 139.395 26.185 139.775 26.565 ;
        RECT 141.180 26.185 141.560 26.565 ;
        RECT 36.420 26.015 36.800 26.065 ;
        RECT 37.560 26.015 37.940 26.065 ;
        RECT 36.420 25.735 37.940 26.015 ;
        RECT 36.420 25.685 36.800 25.735 ;
        RECT 37.560 25.685 37.940 25.735 ;
        RECT 68.870 26.015 69.250 26.065 ;
        RECT 70.010 26.015 70.390 26.065 ;
        RECT 68.870 25.735 70.390 26.015 ;
        RECT 68.870 25.685 69.250 25.735 ;
        RECT 70.010 25.685 70.390 25.735 ;
        RECT 101.320 26.015 101.700 26.065 ;
        RECT 102.460 26.015 102.840 26.065 ;
        RECT 101.320 25.735 102.840 26.015 ;
        RECT 101.320 25.685 101.700 25.735 ;
        RECT 102.460 25.685 102.840 25.735 ;
        RECT 133.770 26.015 134.150 26.065 ;
        RECT 134.910 26.015 135.290 26.065 ;
        RECT 133.770 25.735 135.290 26.015 ;
        RECT 133.770 25.685 134.150 25.735 ;
        RECT 134.910 25.685 135.290 25.735 ;
        RECT 0.240 24.685 0.620 25.065 ;
        RECT 4.160 24.685 4.540 25.065 ;
        RECT 6.700 24.405 9.560 24.785 ;
        RECT 39.150 24.405 42.010 24.785 ;
        RECT 71.600 24.405 74.460 24.785 ;
        RECT 104.050 24.405 106.910 24.785 ;
        RECT 37.560 23.845 38.080 24.225 ;
        RECT 70.010 23.845 70.530 24.225 ;
        RECT 102.460 23.845 102.980 24.225 ;
        RECT 134.910 23.845 135.430 24.225 ;
        RECT 137.355 23.185 137.735 23.565 ;
        RECT 139.395 23.185 139.775 23.565 ;
        RECT 141.180 23.185 141.560 23.565 ;
        RECT 0.240 21.685 0.620 22.065 ;
        RECT 4.160 21.685 4.540 22.065 ;
        RECT 0.240 18.685 0.620 19.065 ;
        RECT 137.355 17.185 137.735 17.565 ;
        RECT 139.395 17.185 139.775 17.565 ;
        RECT 141.180 17.185 141.560 17.565 ;
        RECT 0.240 15.685 0.620 16.065 ;
        RECT 4.160 15.685 4.540 16.065 ;
        RECT 37.060 15.280 37.940 15.660 ;
        RECT 69.510 15.280 70.390 15.660 ;
        RECT 101.960 15.280 102.840 15.660 ;
        RECT 134.410 15.280 135.290 15.660 ;
        RECT 6.700 14.720 9.560 15.100 ;
        RECT 39.150 14.720 42.010 15.100 ;
        RECT 71.600 14.720 74.460 15.100 ;
        RECT 104.050 14.720 106.910 15.100 ;
        RECT 137.355 14.185 137.735 14.565 ;
        RECT 139.395 14.185 139.775 14.565 ;
        RECT 141.180 14.185 141.560 14.565 ;
        RECT 35.780 13.770 36.160 13.820 ;
        RECT 37.560 13.770 37.940 13.820 ;
        RECT 35.780 13.490 37.940 13.770 ;
        RECT 35.780 13.440 36.160 13.490 ;
        RECT 37.560 13.440 37.940 13.490 ;
        RECT 68.230 13.770 68.610 13.820 ;
        RECT 70.010 13.770 70.390 13.820 ;
        RECT 68.230 13.490 70.390 13.770 ;
        RECT 68.230 13.440 68.610 13.490 ;
        RECT 70.010 13.440 70.390 13.490 ;
        RECT 100.680 13.770 101.060 13.820 ;
        RECT 102.460 13.770 102.840 13.820 ;
        RECT 100.680 13.490 102.840 13.770 ;
        RECT 100.680 13.440 101.060 13.490 ;
        RECT 102.460 13.440 102.840 13.490 ;
        RECT 133.130 13.770 133.510 13.820 ;
        RECT 134.910 13.770 135.290 13.820 ;
        RECT 133.130 13.490 135.290 13.770 ;
        RECT 133.130 13.440 133.510 13.490 ;
        RECT 134.910 13.440 135.290 13.490 ;
        RECT 0.240 12.685 0.620 13.065 ;
        RECT 4.160 12.685 4.540 13.065 ;
        RECT 6.700 12.880 9.560 13.260 ;
        RECT 39.150 12.880 42.010 13.260 ;
        RECT 71.600 12.880 74.460 13.260 ;
        RECT 104.050 12.880 106.910 13.260 ;
        RECT 34.500 11.925 34.880 11.975 ;
        RECT 37.560 11.925 37.940 11.975 ;
        RECT 34.500 11.645 37.940 11.925 ;
        RECT 34.500 11.595 34.880 11.645 ;
        RECT 37.560 11.595 37.940 11.645 ;
        RECT 66.950 11.925 67.330 11.975 ;
        RECT 70.010 11.925 70.390 11.975 ;
        RECT 66.950 11.645 70.390 11.925 ;
        RECT 66.950 11.595 67.330 11.645 ;
        RECT 70.010 11.595 70.390 11.645 ;
        RECT 99.400 11.925 99.780 11.975 ;
        RECT 102.460 11.925 102.840 11.975 ;
        RECT 99.400 11.645 102.840 11.925 ;
        RECT 99.400 11.595 99.780 11.645 ;
        RECT 102.460 11.595 102.840 11.645 ;
        RECT 131.850 11.925 132.230 11.975 ;
        RECT 134.910 11.925 135.290 11.975 ;
        RECT 131.850 11.645 135.290 11.925 ;
        RECT 131.850 11.595 132.230 11.645 ;
        RECT 134.910 11.595 135.290 11.645 ;
        RECT 6.700 11.035 9.560 11.415 ;
        RECT 39.150 11.035 42.010 11.415 ;
        RECT 71.600 11.035 74.460 11.415 ;
        RECT 104.050 11.035 106.910 11.415 ;
        RECT 137.355 11.185 137.735 11.565 ;
        RECT 139.395 11.185 139.775 11.565 ;
        RECT 141.180 11.185 141.560 11.565 ;
        RECT 6.700 10.275 9.560 10.655 ;
        RECT 39.150 10.275 42.010 10.655 ;
        RECT 71.600 10.275 74.460 10.655 ;
        RECT 104.050 10.275 106.910 10.655 ;
        RECT 0.240 9.685 0.620 10.065 ;
        RECT 4.160 9.685 4.540 10.065 ;
        RECT 33.220 9.285 33.600 9.335 ;
        RECT 37.560 9.285 37.940 9.335 ;
        RECT 33.220 9.005 37.940 9.285 ;
        RECT 33.220 8.955 33.600 9.005 ;
        RECT 37.560 8.955 37.940 9.005 ;
        RECT 65.670 9.285 66.050 9.335 ;
        RECT 70.010 9.285 70.390 9.335 ;
        RECT 65.670 9.005 70.390 9.285 ;
        RECT 65.670 8.955 66.050 9.005 ;
        RECT 70.010 8.955 70.390 9.005 ;
        RECT 98.120 9.285 98.500 9.335 ;
        RECT 102.460 9.285 102.840 9.335 ;
        RECT 98.120 9.005 102.840 9.285 ;
        RECT 98.120 8.955 98.500 9.005 ;
        RECT 102.460 8.955 102.840 9.005 ;
        RECT 130.570 9.285 130.950 9.335 ;
        RECT 134.910 9.285 135.290 9.335 ;
        RECT 130.570 9.005 135.290 9.285 ;
        RECT 130.570 8.955 130.950 9.005 ;
        RECT 134.910 8.955 135.290 9.005 ;
        RECT 6.700 8.395 9.560 8.775 ;
        RECT 39.150 8.395 42.010 8.775 ;
        RECT 71.600 8.395 74.460 8.775 ;
        RECT 104.050 8.395 106.910 8.775 ;
        RECT 137.355 8.185 137.735 8.565 ;
        RECT 139.395 8.185 139.775 8.565 ;
        RECT 141.180 8.185 141.560 8.565 ;
        RECT 31.940 7.445 32.320 7.495 ;
        RECT 37.560 7.445 37.940 7.495 ;
        RECT 31.940 7.165 37.940 7.445 ;
        RECT 31.940 7.115 32.320 7.165 ;
        RECT 37.560 7.115 37.940 7.165 ;
        RECT 64.390 7.445 64.770 7.495 ;
        RECT 70.010 7.445 70.390 7.495 ;
        RECT 64.390 7.165 70.390 7.445 ;
        RECT 64.390 7.115 64.770 7.165 ;
        RECT 70.010 7.115 70.390 7.165 ;
        RECT 96.840 7.445 97.220 7.495 ;
        RECT 102.460 7.445 102.840 7.495 ;
        RECT 96.840 7.165 102.840 7.445 ;
        RECT 96.840 7.115 97.220 7.165 ;
        RECT 102.460 7.115 102.840 7.165 ;
        RECT 129.290 7.445 129.670 7.495 ;
        RECT 134.910 7.445 135.290 7.495 ;
        RECT 129.290 7.165 135.290 7.445 ;
        RECT 129.290 7.115 129.670 7.165 ;
        RECT 134.910 7.115 135.290 7.165 ;
        RECT 0.240 6.685 0.620 7.065 ;
        RECT 4.160 6.685 4.540 7.065 ;
        RECT 6.700 6.555 9.560 6.935 ;
        RECT 39.150 6.555 42.010 6.935 ;
        RECT 71.600 6.555 74.460 6.935 ;
        RECT 104.050 6.555 106.910 6.935 ;
        RECT 30.660 5.600 31.040 5.650 ;
        RECT 37.560 5.600 37.940 5.650 ;
        RECT 30.660 5.320 37.940 5.600 ;
        RECT 30.660 5.270 31.040 5.320 ;
        RECT 37.560 5.270 37.940 5.320 ;
        RECT 63.110 5.600 63.490 5.650 ;
        RECT 70.010 5.600 70.390 5.650 ;
        RECT 63.110 5.320 70.390 5.600 ;
        RECT 63.110 5.270 63.490 5.320 ;
        RECT 70.010 5.270 70.390 5.320 ;
        RECT 95.560 5.600 95.940 5.650 ;
        RECT 102.460 5.600 102.840 5.650 ;
        RECT 95.560 5.320 102.840 5.600 ;
        RECT 95.560 5.270 95.940 5.320 ;
        RECT 102.460 5.270 102.840 5.320 ;
        RECT 128.010 5.600 128.390 5.650 ;
        RECT 134.910 5.600 135.290 5.650 ;
        RECT 128.010 5.320 135.290 5.600 ;
        RECT 128.010 5.270 128.390 5.320 ;
        RECT 134.910 5.270 135.290 5.320 ;
        RECT 137.355 5.185 137.735 5.565 ;
        RECT 139.395 5.185 139.775 5.565 ;
        RECT 141.180 5.185 141.560 5.565 ;
        RECT 6.700 4.710 9.560 5.090 ;
        RECT 39.150 4.710 42.010 5.090 ;
        RECT 71.600 4.710 74.460 5.090 ;
        RECT 104.050 4.710 106.910 5.090 ;
        RECT 0.240 3.685 0.620 4.065 ;
        RECT 4.160 3.685 4.540 4.065 ;
        RECT 6.700 3.950 9.560 4.330 ;
        RECT 39.150 3.950 42.010 4.330 ;
        RECT 71.600 3.950 74.460 4.330 ;
        RECT 104.050 3.950 106.910 4.330 ;
        RECT 29.380 2.960 29.760 3.010 ;
        RECT 37.560 2.960 37.940 3.010 ;
        RECT 29.380 2.680 37.940 2.960 ;
        RECT 29.380 2.630 29.760 2.680 ;
        RECT 37.560 2.630 37.940 2.680 ;
        RECT 61.830 2.960 62.210 3.010 ;
        RECT 70.010 2.960 70.390 3.010 ;
        RECT 61.830 2.680 70.390 2.960 ;
        RECT 61.830 2.630 62.210 2.680 ;
        RECT 70.010 2.630 70.390 2.680 ;
        RECT 94.280 2.960 94.660 3.010 ;
        RECT 102.460 2.960 102.840 3.010 ;
        RECT 94.280 2.680 102.840 2.960 ;
        RECT 94.280 2.630 94.660 2.680 ;
        RECT 102.460 2.630 102.840 2.680 ;
        RECT 126.730 2.960 127.110 3.010 ;
        RECT 134.910 2.960 135.290 3.010 ;
        RECT 126.730 2.680 135.290 2.960 ;
        RECT 126.730 2.630 127.110 2.680 ;
        RECT 134.910 2.630 135.290 2.680 ;
        RECT 6.700 2.070 9.560 2.450 ;
        RECT 39.150 2.070 42.010 2.450 ;
        RECT 71.600 2.070 74.460 2.450 ;
        RECT 104.050 2.070 106.910 2.450 ;
        RECT 137.355 2.185 137.735 2.565 ;
        RECT 139.395 2.185 139.775 2.565 ;
        RECT 141.180 2.185 141.560 2.565 ;
        RECT 28.100 1.120 28.480 1.170 ;
        RECT 37.560 1.120 37.940 1.170 ;
        RECT 0.240 0.685 0.620 1.065 ;
        RECT 4.160 0.685 4.540 1.065 ;
        RECT 28.100 0.840 37.940 1.120 ;
        RECT 28.100 0.790 28.480 0.840 ;
        RECT 37.560 0.790 37.940 0.840 ;
        RECT 60.550 1.120 60.930 1.170 ;
        RECT 70.010 1.120 70.390 1.170 ;
        RECT 60.550 0.840 70.390 1.120 ;
        RECT 60.550 0.790 60.930 0.840 ;
        RECT 70.010 0.790 70.390 0.840 ;
        RECT 93.000 1.120 93.380 1.170 ;
        RECT 102.460 1.120 102.840 1.170 ;
        RECT 93.000 0.840 102.840 1.120 ;
        RECT 93.000 0.790 93.380 0.840 ;
        RECT 102.460 0.790 102.840 0.840 ;
        RECT 125.450 1.120 125.830 1.170 ;
        RECT 134.910 1.120 135.290 1.170 ;
        RECT 125.450 0.840 135.290 1.120 ;
        RECT 125.450 0.790 125.830 0.840 ;
        RECT 134.910 0.790 135.290 0.840 ;
        RECT 6.700 0.230 9.560 0.610 ;
        RECT 39.150 0.230 42.010 0.610 ;
        RECT 71.600 0.230 74.460 0.610 ;
        RECT 104.050 0.230 106.910 0.610 ;
  END
END efuse_array_64x8
END LIBRARY

