module efuse_wb_mem_64x8 (wb_ack_o,
    wb_clk_i,
    wb_cyc_i,
    wb_rst_i,
    wb_stb_i,
    wb_we_i,
    write_disable_i,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o);
 output wb_ack_o;
 input wb_clk_i;
 input wb_cyc_i;
 input wb_rst_i;
 input wb_stb_i;
 input wb_we_i;
 input write_disable_i;
 input [7:0] wb_adr_i;
 input [7:0] wb_dat_i;
 output [7:0] wb_dat_o;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire \bit_sel[0] ;
 wire \bit_sel[10] ;
 wire \bit_sel[11] ;
 wire \bit_sel[12] ;
 wire \bit_sel[13] ;
 wire \bit_sel[14] ;
 wire \bit_sel[15] ;
 wire \bit_sel[16] ;
 wire \bit_sel[17] ;
 wire \bit_sel[18] ;
 wire \bit_sel[19] ;
 wire \bit_sel[1] ;
 wire \bit_sel[20] ;
 wire \bit_sel[21] ;
 wire \bit_sel[22] ;
 wire \bit_sel[23] ;
 wire \bit_sel[24] ;
 wire \bit_sel[25] ;
 wire \bit_sel[26] ;
 wire \bit_sel[27] ;
 wire \bit_sel[28] ;
 wire \bit_sel[29] ;
 wire \bit_sel[2] ;
 wire \bit_sel[30] ;
 wire \bit_sel[31] ;
 wire \bit_sel[32] ;
 wire \bit_sel[33] ;
 wire \bit_sel[34] ;
 wire \bit_sel[35] ;
 wire \bit_sel[36] ;
 wire \bit_sel[37] ;
 wire \bit_sel[38] ;
 wire \bit_sel[39] ;
 wire \bit_sel[3] ;
 wire \bit_sel[40] ;
 wire \bit_sel[41] ;
 wire \bit_sel[42] ;
 wire \bit_sel[43] ;
 wire \bit_sel[44] ;
 wire \bit_sel[45] ;
 wire \bit_sel[46] ;
 wire \bit_sel[47] ;
 wire \bit_sel[48] ;
 wire \bit_sel[49] ;
 wire \bit_sel[4] ;
 wire \bit_sel[50] ;
 wire \bit_sel[51] ;
 wire \bit_sel[52] ;
 wire \bit_sel[53] ;
 wire \bit_sel[54] ;
 wire \bit_sel[55] ;
 wire \bit_sel[56] ;
 wire \bit_sel[57] ;
 wire \bit_sel[58] ;
 wire \bit_sel[59] ;
 wire \bit_sel[5] ;
 wire \bit_sel[60] ;
 wire \bit_sel[61] ;
 wire \bit_sel[62] ;
 wire \bit_sel[63] ;
 wire \bit_sel[6] ;
 wire \bit_sel[7] ;
 wire \bit_sel[8] ;
 wire \bit_sel[9] ;
 wire \bit_sel_reg[0] ;
 wire \bit_sel_reg[10] ;
 wire \bit_sel_reg[11] ;
 wire \bit_sel_reg[12] ;
 wire \bit_sel_reg[13] ;
 wire \bit_sel_reg[14] ;
 wire \bit_sel_reg[15] ;
 wire \bit_sel_reg[16] ;
 wire \bit_sel_reg[17] ;
 wire \bit_sel_reg[18] ;
 wire \bit_sel_reg[19] ;
 wire \bit_sel_reg[1] ;
 wire \bit_sel_reg[20] ;
 wire \bit_sel_reg[21] ;
 wire \bit_sel_reg[22] ;
 wire \bit_sel_reg[23] ;
 wire \bit_sel_reg[24] ;
 wire \bit_sel_reg[25] ;
 wire \bit_sel_reg[26] ;
 wire \bit_sel_reg[27] ;
 wire \bit_sel_reg[28] ;
 wire \bit_sel_reg[29] ;
 wire \bit_sel_reg[2] ;
 wire \bit_sel_reg[30] ;
 wire \bit_sel_reg[31] ;
 wire \bit_sel_reg[32] ;
 wire \bit_sel_reg[33] ;
 wire \bit_sel_reg[34] ;
 wire \bit_sel_reg[35] ;
 wire \bit_sel_reg[36] ;
 wire \bit_sel_reg[37] ;
 wire \bit_sel_reg[38] ;
 wire \bit_sel_reg[39] ;
 wire \bit_sel_reg[3] ;
 wire \bit_sel_reg[40] ;
 wire \bit_sel_reg[41] ;
 wire \bit_sel_reg[42] ;
 wire \bit_sel_reg[43] ;
 wire \bit_sel_reg[44] ;
 wire \bit_sel_reg[45] ;
 wire \bit_sel_reg[46] ;
 wire \bit_sel_reg[47] ;
 wire \bit_sel_reg[48] ;
 wire \bit_sel_reg[49] ;
 wire \bit_sel_reg[4] ;
 wire \bit_sel_reg[50] ;
 wire \bit_sel_reg[51] ;
 wire \bit_sel_reg[52] ;
 wire \bit_sel_reg[53] ;
 wire \bit_sel_reg[54] ;
 wire \bit_sel_reg[55] ;
 wire \bit_sel_reg[56] ;
 wire \bit_sel_reg[57] ;
 wire \bit_sel_reg[58] ;
 wire \bit_sel_reg[59] ;
 wire \bit_sel_reg[5] ;
 wire \bit_sel_reg[60] ;
 wire \bit_sel_reg[61] ;
 wire \bit_sel_reg[62] ;
 wire \bit_sel_reg[63] ;
 wire \bit_sel_reg[6] ;
 wire \bit_sel_reg[7] ;
 wire \bit_sel_reg[8] ;
 wire \bit_sel_reg[9] ;
 wire \col_prog_n[0] ;
 wire \col_prog_n[1] ;
 wire \col_prog_n[2] ;
 wire \col_prog_n[3] ;
 wire \col_prog_n[4] ;
 wire \col_prog_n[5] ;
 wire \col_prog_n[6] ;
 wire \col_prog_n[7] ;
 wire \col_prog_n_reg[0] ;
 wire \col_prog_n_reg[1] ;
 wire \col_prog_n_reg[2] ;
 wire \col_prog_n_reg[3] ;
 wire \col_prog_n_reg[4] ;
 wire \col_prog_n_reg[5] ;
 wire \col_prog_n_reg[6] ;
 wire \col_prog_n_reg[7] ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \efuse_out[0] ;
 wire \efuse_out[1] ;
 wire \efuse_out[2] ;
 wire \efuse_out[3] ;
 wire \efuse_out[4] ;
 wire \efuse_out[5] ;
 wire \efuse_out[6] ;
 wire \efuse_out[7] ;
 wire preset_n;
 wire preset_n_reg;
 wire sense;
 wire sense_reg;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _369_ (.I(preset_n_reg),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _370_ (.I(\col_prog_n_reg[7] ),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _371_ (.I(\state[3] ),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _372_ (.I(\col_prog_n_reg[6] ),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _373_ (.I(\col_prog_n_reg[5] ),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _374_ (.I(\col_prog_n_reg[4] ),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _375_ (.I(\col_prog_n_reg[3] ),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _376_ (.I(\col_prog_n_reg[2] ),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _377_ (.I(\col_prog_n_reg[1] ),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _378_ (.I(\col_prog_n_reg[0] ),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _379_ (.I(net29),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _380_ (.I(\state[1] ),
    .ZN(_194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _381_ (.I(\state[0] ),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _382_ (.I(\counter[4] ),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _383_ (.I(\counter[7] ),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _384_ (.I(net26),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _385_ (.I(net28),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _386_ (.I(net16),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _387_ (.I(net12),
    .ZN(_200_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _388_ (.I(net11),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _389_ (.I(net14),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _390_ (.I(net15),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _391_ (.A1(net17),
    .A2(net27),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _392_ (.A1(net29),
    .A2(_195_),
    .A3(net28),
    .A4(_204_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _393_ (.A1(_195_),
    .A2(_000_),
    .Z(_205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _394_ (.A1(\state[2] ),
    .A2(_205_),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _395_ (.A1(_183_),
    .A2(_000_),
    .B(_206_),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _396_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .A3(\counter[2] ),
    .Z(_207_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _397_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .A3(\counter[3] ),
    .A4(\counter[2] ),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _398_ (.A1(\counter[5] ),
    .A2(\counter[4] ),
    .A3(\counter[7] ),
    .A4(\counter[6] ),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _399_ (.A1(_208_),
    .A2(_209_),
    .ZN(_210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _400_ (.A1(\counter[9] ),
    .A2(\counter[8] ),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _401_ (.A1(_208_),
    .A2(_209_),
    .A3(_211_),
    .ZN(_212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _402_ (.A1(\state[3] ),
    .A2(_212_),
    .Z(_213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _403_ (.A1(\state[3] ),
    .A2(_212_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _404_ (.A1(_184_),
    .A2(_185_),
    .B1(net25),
    .B2(_213_),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _405_ (.A1(_185_),
    .A2(_186_),
    .B1(net24),
    .B2(_213_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _406_ (.A1(_185_),
    .A2(_187_),
    .B1(net23),
    .B2(_213_),
    .ZN(_179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _407_ (.A1(_185_),
    .A2(_188_),
    .B1(net22),
    .B2(_213_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _408_ (.A1(_185_),
    .A2(_189_),
    .B1(net21),
    .B2(_213_),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _409_ (.A1(_185_),
    .A2(_190_),
    .B1(net20),
    .B2(_213_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _410_ (.A1(_185_),
    .A2(_191_),
    .B1(net19),
    .B2(_213_),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _411_ (.A1(_185_),
    .A2(_192_),
    .B1(net18),
    .B2(_213_),
    .ZN(_174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _412_ (.A1(\state[2] ),
    .A2(\state[0] ),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _413_ (.I(_215_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _414_ (.A1(\bit_sel_reg[63] ),
    .A2(net42),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _415_ (.A1(net12),
    .A2(net11),
    .ZN(_218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _416_ (.A1(net12),
    .A2(net11),
    .A3(net13),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _417_ (.I(_219_),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _418_ (.A1(net14),
    .A2(net15),
    .A3(_220_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _419_ (.A1(net29),
    .A2(_198_),
    .A3(_204_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _420_ (.A1(\state[0] ),
    .A2(_222_),
    .ZN(_223_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _421_ (.A1(\state[2] ),
    .A2(_222_),
    .B(_216_),
    .C(net16),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _422_ (.A1(_221_),
    .A2(net41),
    .B(_217_),
    .ZN(_173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _423_ (.A1(\bit_sel_reg[62] ),
    .A2(net42),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _424_ (.A1(net12),
    .A2(_201_),
    .A3(net13),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _425_ (.A1(_202_),
    .A2(_203_),
    .A3(_226_),
    .Z(_227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _426_ (.A1(net40),
    .A2(_227_),
    .B(_225_),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _427_ (.A1(\bit_sel_reg[61] ),
    .A2(net42),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _428_ (.A1(_200_),
    .A2(net11),
    .A3(net13),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _429_ (.A1(_202_),
    .A2(_203_),
    .A3(_229_),
    .Z(_230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _430_ (.A1(net41),
    .A2(_230_),
    .B(_228_),
    .ZN(_171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _431_ (.A1(\bit_sel_reg[60] ),
    .A2(net42),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _432_ (.A1(net12),
    .A2(net11),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _433_ (.A1(net13),
    .A2(net14),
    .A3(net15),
    .A4(_232_),
    .ZN(_233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _434_ (.A1(net41),
    .A2(_233_),
    .B(_231_),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _435_ (.A1(\bit_sel_reg[59] ),
    .A2(net43),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _436_ (.A1(net13),
    .A2(_218_),
    .ZN(_235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _437_ (.A1(net14),
    .A2(net15),
    .A3(_235_),
    .ZN(_236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _438_ (.A1(_224_),
    .A2(_236_),
    .B(_234_),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _439_ (.A1(\bit_sel_reg[58] ),
    .A2(net42),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _440_ (.A1(_200_),
    .A2(net11),
    .A3(net13),
    .ZN(_238_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _441_ (.A1(net14),
    .A2(net15),
    .A3(_238_),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _442_ (.A1(net41),
    .A2(_239_),
    .B(_237_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _443_ (.A1(\bit_sel_reg[57] ),
    .A2(net42),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _444_ (.A1(net12),
    .A2(_201_),
    .A3(net13),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _445_ (.A1(net14),
    .A2(net15),
    .A3(_241_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _446_ (.A1(net41),
    .A2(_242_),
    .B(_240_),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _447_ (.A1(\bit_sel_reg[56] ),
    .A2(net42),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _448_ (.A1(net12),
    .A2(net11),
    .A3(net13),
    .ZN(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _449_ (.A1(net14),
    .A2(net15),
    .A3(_244_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _450_ (.A1(net41),
    .A2(_245_),
    .B(_243_),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _451_ (.A1(\bit_sel_reg[55] ),
    .A2(net42),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _452_ (.A1(net14),
    .A2(_219_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _453_ (.A1(net15),
    .A2(_247_),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _454_ (.A1(net41),
    .A2(_248_),
    .B(_246_),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _455_ (.A1(\bit_sel_reg[54] ),
    .A2(net43),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _456_ (.A1(net14),
    .A2(_226_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _457_ (.A1(net15),
    .A2(_250_),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _458_ (.A1(net40),
    .A2(_251_),
    .B(_249_),
    .ZN(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _459_ (.A1(\bit_sel_reg[53] ),
    .A2(net42),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _460_ (.A1(net14),
    .A2(_229_),
    .ZN(_253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _461_ (.A1(net15),
    .A2(_253_),
    .ZN(_254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _462_ (.A1(net41),
    .A2(_254_),
    .B(_252_),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _463_ (.A1(\bit_sel_reg[52] ),
    .A2(net43),
    .ZN(_255_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _464_ (.A1(net13),
    .A2(_202_),
    .A3(_232_),
    .Z(_256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _465_ (.A1(net15),
    .A2(_256_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _466_ (.A1(net40),
    .A2(_257_),
    .B(_255_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _467_ (.A1(\bit_sel_reg[51] ),
    .A2(net42),
    .ZN(_258_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _468_ (.A1(net13),
    .A2(net14),
    .A3(_218_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _469_ (.A1(net15),
    .A2(_259_),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _470_ (.A1(_224_),
    .A2(_260_),
    .B(_258_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _471_ (.A1(\bit_sel_reg[50] ),
    .A2(net42),
    .ZN(_261_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _472_ (.A1(_202_),
    .A2(_238_),
    .Z(_262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _473_ (.A1(net15),
    .A2(_262_),
    .ZN(_263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _474_ (.A1(net41),
    .A2(_263_),
    .B(_261_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _475_ (.A1(\bit_sel_reg[49] ),
    .A2(net42),
    .ZN(_264_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _476_ (.A1(_202_),
    .A2(_241_),
    .Z(_265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _477_ (.A1(net15),
    .A2(_265_),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _478_ (.A1(net41),
    .A2(_266_),
    .B(_264_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _479_ (.A1(\bit_sel_reg[48] ),
    .A2(net42),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _480_ (.A1(_202_),
    .A2(_244_),
    .Z(_268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _481_ (.A1(net15),
    .A2(_268_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _482_ (.A1(net41),
    .A2(_269_),
    .B(_267_),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _483_ (.A1(\bit_sel_reg[47] ),
    .A2(net43),
    .ZN(_270_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _484_ (.A1(net14),
    .A2(_203_),
    .A3(_220_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _485_ (.A1(net40),
    .A2(_271_),
    .B(_270_),
    .ZN(_157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _486_ (.A1(\bit_sel_reg[46] ),
    .A2(net43),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _487_ (.A1(_202_),
    .A2(net15),
    .A3(_226_),
    .ZN(_273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _488_ (.I(_273_),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _489_ (.A1(net40),
    .A2(_274_),
    .B(_272_),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _490_ (.A1(\bit_sel_reg[45] ),
    .A2(net43),
    .ZN(_275_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _491_ (.A1(_202_),
    .A2(net15),
    .A3(_229_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _492_ (.I(_276_),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _493_ (.A1(net40),
    .A2(_277_),
    .B(_275_),
    .ZN(_155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _494_ (.A1(\bit_sel_reg[44] ),
    .A2(net43),
    .ZN(_278_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _495_ (.A1(net13),
    .A2(net14),
    .A3(_203_),
    .A4(_232_),
    .ZN(_279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _496_ (.A1(net40),
    .A2(_279_),
    .B(_278_),
    .ZN(_154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _497_ (.A1(\bit_sel_reg[43] ),
    .A2(net42),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _498_ (.A1(net14),
    .A2(_203_),
    .A3(_235_),
    .ZN(_281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _499_ (.A1(_224_),
    .A2(_281_),
    .B(_280_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _500_ (.A1(\bit_sel_reg[42] ),
    .A2(net43),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _501_ (.A1(net14),
    .A2(_203_),
    .A3(_238_),
    .ZN(_283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _502_ (.A1(net40),
    .A2(_283_),
    .B(_282_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _503_ (.A1(\bit_sel_reg[41] ),
    .A2(net43),
    .ZN(_284_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _504_ (.A1(net14),
    .A2(_203_),
    .A3(_241_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _505_ (.A1(net40),
    .A2(_285_),
    .B(_284_),
    .ZN(_151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _506_ (.A1(\bit_sel_reg[40] ),
    .A2(net43),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _507_ (.A1(net14),
    .A2(_203_),
    .A3(_244_),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _508_ (.A1(net41),
    .A2(_287_),
    .B(_286_),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _509_ (.A1(\bit_sel_reg[39] ),
    .A2(net43),
    .ZN(_288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _510_ (.A1(_203_),
    .A2(_247_),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _511_ (.A1(net40),
    .A2(_289_),
    .B(_288_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _512_ (.A1(\bit_sel_reg[38] ),
    .A2(net43),
    .ZN(_290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _513_ (.A1(_203_),
    .A2(_250_),
    .ZN(_291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _514_ (.A1(net40),
    .A2(_291_),
    .B(_290_),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _515_ (.A1(\bit_sel_reg[37] ),
    .A2(net42),
    .ZN(_292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _516_ (.A1(_203_),
    .A2(_253_),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _517_ (.A1(net41),
    .A2(_293_),
    .B(_292_),
    .ZN(_147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _518_ (.A1(\bit_sel_reg[36] ),
    .A2(net43),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _519_ (.A1(_203_),
    .A2(_256_),
    .ZN(_295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _520_ (.A1(net40),
    .A2(_295_),
    .B(_294_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _521_ (.A1(\bit_sel_reg[35] ),
    .A2(net43),
    .ZN(_296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _522_ (.A1(_203_),
    .A2(_259_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _523_ (.A1(_224_),
    .A2(_297_),
    .B(_296_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _524_ (.A1(\bit_sel_reg[34] ),
    .A2(net43),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _525_ (.A1(_203_),
    .A2(_262_),
    .ZN(_299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _526_ (.A1(net40),
    .A2(_299_),
    .B(_298_),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _527_ (.A1(\bit_sel_reg[33] ),
    .A2(net43),
    .ZN(_300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _528_ (.A1(_203_),
    .A2(_265_),
    .ZN(_301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _529_ (.A1(net40),
    .A2(_301_),
    .B(_300_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _530_ (.A1(\bit_sel_reg[32] ),
    .A2(net42),
    .ZN(_302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _531_ (.A1(_203_),
    .A2(_268_),
    .ZN(_303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _532_ (.A1(net41),
    .A2(_303_),
    .B(_302_),
    .ZN(_142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _533_ (.A1(\bit_sel_reg[31] ),
    .A2(net42),
    .ZN(_304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _534_ (.A1(\state[2] ),
    .A2(_222_),
    .B(_216_),
    .C(_199_),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _535_ (.A1(_221_),
    .A2(net39),
    .B(_304_),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _536_ (.A1(\bit_sel_reg[30] ),
    .A2(net42),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _537_ (.A1(_227_),
    .A2(net38),
    .B(_306_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _538_ (.A1(\bit_sel_reg[29] ),
    .A2(net42),
    .ZN(_307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _539_ (.A1(_230_),
    .A2(net38),
    .B(_307_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _540_ (.A1(\bit_sel_reg[28] ),
    .A2(net42),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _541_ (.A1(_233_),
    .A2(net38),
    .B(_308_),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _542_ (.A1(\bit_sel_reg[27] ),
    .A2(net43),
    .ZN(_309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _543_ (.A1(_236_),
    .A2(_305_),
    .B(_309_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _544_ (.A1(\bit_sel_reg[26] ),
    .A2(net42),
    .ZN(_310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _545_ (.A1(_239_),
    .A2(net38),
    .B(_310_),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _546_ (.A1(\bit_sel_reg[25] ),
    .A2(net42),
    .ZN(_311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _547_ (.A1(_242_),
    .A2(net38),
    .B(_311_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _548_ (.A1(\bit_sel_reg[24] ),
    .A2(net42),
    .ZN(_312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _549_ (.A1(_245_),
    .A2(net39),
    .B(_312_),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _550_ (.A1(\bit_sel_reg[23] ),
    .A2(net42),
    .ZN(_313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _551_ (.A1(_248_),
    .A2(net39),
    .B(_313_),
    .ZN(_133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _552_ (.A1(\bit_sel_reg[22] ),
    .A2(net43),
    .ZN(_314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _553_ (.A1(_251_),
    .A2(net38),
    .B(_314_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _554_ (.A1(\bit_sel_reg[21] ),
    .A2(net42),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _555_ (.A1(_254_),
    .A2(net38),
    .B(_315_),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _556_ (.A1(\bit_sel_reg[20] ),
    .A2(net43),
    .ZN(_316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _557_ (.A1(_257_),
    .A2(net39),
    .B(_316_),
    .ZN(_130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _558_ (.A1(\bit_sel_reg[19] ),
    .A2(net42),
    .ZN(_317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _559_ (.A1(_260_),
    .A2(_305_),
    .B(_317_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _560_ (.A1(\bit_sel_reg[18] ),
    .A2(net42),
    .ZN(_318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _561_ (.A1(_263_),
    .A2(net38),
    .B(_318_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _562_ (.A1(\bit_sel_reg[17] ),
    .A2(net42),
    .ZN(_319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _563_ (.A1(_266_),
    .A2(net38),
    .B(_319_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _564_ (.A1(\bit_sel_reg[16] ),
    .A2(net42),
    .ZN(_320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _565_ (.A1(_269_),
    .A2(net38),
    .B(_320_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _566_ (.A1(\bit_sel_reg[15] ),
    .A2(net43),
    .ZN(_321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _567_ (.A1(_271_),
    .A2(net39),
    .B(_321_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _568_ (.A1(\bit_sel_reg[14] ),
    .A2(net43),
    .ZN(_322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _569_ (.A1(_274_),
    .A2(net39),
    .B(_322_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _570_ (.A1(\bit_sel_reg[13] ),
    .A2(net43),
    .ZN(_323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _571_ (.A1(_277_),
    .A2(net39),
    .B(_323_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _572_ (.A1(\bit_sel_reg[12] ),
    .A2(net43),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _573_ (.A1(_279_),
    .A2(net39),
    .B(_324_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _574_ (.A1(\bit_sel_reg[11] ),
    .A2(net42),
    .ZN(_325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _575_ (.A1(_281_),
    .A2(_305_),
    .B(_325_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _576_ (.A1(\bit_sel_reg[10] ),
    .A2(net43),
    .ZN(_326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _577_ (.A1(_283_),
    .A2(net39),
    .B(_326_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _578_ (.A1(\bit_sel_reg[9] ),
    .A2(net43),
    .ZN(_327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _579_ (.A1(_285_),
    .A2(net39),
    .B(_327_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _580_ (.A1(\bit_sel_reg[8] ),
    .A2(net43),
    .ZN(_328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _581_ (.A1(_287_),
    .A2(net39),
    .B(_328_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _582_ (.A1(\bit_sel_reg[7] ),
    .A2(net43),
    .ZN(_329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _583_ (.A1(_289_),
    .A2(net39),
    .B(_329_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _584_ (.A1(\bit_sel_reg[6] ),
    .A2(net43),
    .ZN(_330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _585_ (.A1(_291_),
    .A2(net38),
    .B(_330_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _586_ (.A1(\bit_sel_reg[5] ),
    .A2(net42),
    .ZN(_331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _587_ (.A1(_293_),
    .A2(net38),
    .B(_331_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _588_ (.A1(\bit_sel_reg[4] ),
    .A2(net43),
    .ZN(_332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _589_ (.A1(_295_),
    .A2(net39),
    .B(_332_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _590_ (.A1(\bit_sel_reg[3] ),
    .A2(net43),
    .ZN(_333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _591_ (.A1(_297_),
    .A2(net39),
    .B(_333_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _592_ (.A1(\bit_sel_reg[2] ),
    .A2(net43),
    .ZN(_334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _593_ (.A1(_299_),
    .A2(net38),
    .B(_334_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _594_ (.A1(\bit_sel_reg[1] ),
    .A2(net43),
    .ZN(_335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _595_ (.A1(_301_),
    .A2(net38),
    .B(_335_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _596_ (.A1(\bit_sel_reg[0] ),
    .A2(net42),
    .ZN(_336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _597_ (.A1(_303_),
    .A2(net38),
    .B(_336_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _598_ (.A1(\state[3] ),
    .A2(\state[0] ),
    .ZN(_337_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _599_ (.A1(\state[3] ),
    .A2(\state[1] ),
    .A3(\state[0] ),
    .B(_214_),
    .ZN(_338_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _600_ (.A1(\state[3] ),
    .A2(_208_),
    .A3(_209_),
    .A4(_211_),
    .ZN(_339_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _601_ (.A1(\state[3] ),
    .A2(\state[1] ),
    .A3(_195_),
    .ZN(_340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _602_ (.A1(_193_),
    .A2(_338_),
    .B(_340_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _603_ (.A1(sense_reg),
    .A2(_000_),
    .ZN(_341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _604_ (.A1(\state[1] ),
    .A2(_205_),
    .B(_341_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _605_ (.I0(net37),
    .I1(\efuse_out[7] ),
    .S(\state[1] ),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _606_ (.I0(net36),
    .I1(\efuse_out[6] ),
    .S(\state[1] ),
    .Z(_106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _607_ (.I0(net35),
    .I1(\efuse_out[5] ),
    .S(\state[1] ),
    .Z(_105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _608_ (.I0(net34),
    .I1(\efuse_out[4] ),
    .S(\state[1] ),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _609_ (.I0(net33),
    .I1(\efuse_out[3] ),
    .S(\state[1] ),
    .Z(_103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _610_ (.I0(net32),
    .I1(\efuse_out[2] ),
    .S(\state[1] ),
    .Z(_102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _611_ (.I0(net31),
    .I1(\efuse_out[1] ),
    .S(\state[1] ),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _612_ (.I0(net30),
    .I1(\efuse_out[0] ),
    .S(\state[1] ),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _613_ (.A1(net29),
    .A2(_204_),
    .B(\state[0] ),
    .ZN(_342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _614_ (.A1(_194_),
    .A2(_339_),
    .A3(_342_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _615_ (.A1(_214_),
    .A2(_223_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _616_ (.A1(\state[0] ),
    .A2(_198_),
    .B(_337_),
    .C(net26),
    .ZN(_343_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _617_ (.A1(_342_),
    .A2(_343_),
    .Z(_344_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _618_ (.A1(_339_),
    .A2(_342_),
    .A3(_343_),
    .ZN(_345_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _619_ (.A1(_213_),
    .A2(_344_),
    .Z(_346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _620_ (.A1(_213_),
    .A2(_344_),
    .ZN(_347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _621_ (.A1(\counter[0] ),
    .A2(_345_),
    .ZN(_348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _622_ (.A1(\counter[0] ),
    .A2(_347_),
    .B(_348_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _623_ (.A1(\counter[1] ),
    .A2(_345_),
    .ZN(_349_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _624_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .Z(_350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _625_ (.A1(_347_),
    .A2(_350_),
    .B(_349_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _626_ (.A1(\counter[2] ),
    .A2(_345_),
    .ZN(_351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _627_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .B(\counter[2] ),
    .ZN(_352_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _628_ (.A1(_207_),
    .A2(_352_),
    .Z(_353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _629_ (.A1(_347_),
    .A2(_353_),
    .B(_351_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _630_ (.A1(_185_),
    .A2(_208_),
    .ZN(_354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _631_ (.A1(_207_),
    .A2(_345_),
    .B(\counter[3] ),
    .ZN(_355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _632_ (.A1(_345_),
    .A2(_354_),
    .B(_355_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _633_ (.A1(_345_),
    .A2(_354_),
    .B(\counter[4] ),
    .ZN(_356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _634_ (.A1(_196_),
    .A2(_208_),
    .ZN(_357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _635_ (.A1(_347_),
    .A2(_357_),
    .B(_356_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _636_ (.A1(\counter[5] ),
    .A2(_345_),
    .A3(_357_),
    .Z(_358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _637_ (.A1(_185_),
    .A2(_344_),
    .ZN(_359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _638_ (.A1(_345_),
    .A2(_357_),
    .B(\counter[5] ),
    .ZN(_360_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _639_ (.A1(_358_),
    .A2(_359_),
    .A3(_360_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _640_ (.A1(\counter[5] ),
    .A2(\counter[6] ),
    .A3(_357_),
    .B(\state[3] ),
    .ZN(_361_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _641_ (.A1(_339_),
    .A2(_344_),
    .A3(_361_),
    .ZN(_362_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _642_ (.A1(\counter[5] ),
    .A2(_345_),
    .A3(_357_),
    .B(\counter[6] ),
    .ZN(_363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _643_ (.A1(_362_),
    .A2(_363_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _644_ (.A1(\counter[5] ),
    .A2(_197_),
    .A3(\counter[6] ),
    .A4(_357_),
    .ZN(_364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _645_ (.A1(_197_),
    .A2(_362_),
    .B1(_364_),
    .B2(_346_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _646_ (.A1(\counter[8] ),
    .A2(_210_),
    .ZN(_365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _647_ (.A1(_185_),
    .A2(_365_),
    .ZN(_366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _648_ (.A1(_210_),
    .A2(_345_),
    .B(\counter[8] ),
    .ZN(_367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _649_ (.A1(_345_),
    .A2(_366_),
    .B(_367_),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _650_ (.A1(_185_),
    .A2(_344_),
    .B(\counter[9] ),
    .ZN(_368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _651_ (.A1(_346_),
    .A2(_365_),
    .B(_368_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _652_ (.I(net26),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _653_ (.I(net26),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _654_ (.I(net26),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _655_ (.I(net26),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _656_ (.I(net26),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _657_ (.I(net26),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _658_ (.I(net26),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _659_ (.I(net26),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _660_ (.I(net26),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _661_ (.I(net26),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _662_ (.I(net26),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _663_ (.I(net26),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _664_ (.I(net26),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _665_ (.I(net45),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _666_ (.I(net44),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _667_ (.I(net44),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _668_ (.I(net44),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _669_ (.I(net44),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _670_ (.I(net45),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _671_ (.I(net44),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _672_ (.I(net44),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _673_ (.I(net44),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _674_ (.I(net44),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _675_ (.I(net44),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _676_ (.I(net45),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _677_ (.I(net44),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _678_ (.I(net44),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _679_ (.I(net44),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _680_ (.I(net44),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _681_ (.I(net45),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _682_ (.I(net44),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _683_ (.I(net44),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _684_ (.I(net45),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _685_ (.I(net44),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _686_ (.I(net45),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _687_ (.I(net44),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _688_ (.I(net45),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _689_ (.I(net45),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _690_ (.I(net45),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _691_ (.I(net45),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _692_ (.I(net26),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _693_ (.I(net45),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _694_ (.I(net45),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _695_ (.I(net45),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _696_ (.I(net45),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _697_ (.I(net45),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _698_ (.I(net44),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _699_ (.I(net44),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _700_ (.I(net44),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _701_ (.I(net44),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _702_ (.I(net45),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _703_ (.I(net44),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _704_ (.I(net44),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _705_ (.I(net44),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _706_ (.I(net44),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _707_ (.I(net44),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _708_ (.I(net45),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _709_ (.I(net44),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _710_ (.I(net44),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _711_ (.I(net44),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _712_ (.I(net44),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _713_ (.I(net45),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _714_ (.I(net44),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _715_ (.I(net44),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _716_ (.I(net45),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _717_ (.I(net44),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _718_ (.I(net45),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _719_ (.I(net44),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _720_ (.I(net45),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _721_ (.I(net45),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _722_ (.I(net45),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _723_ (.I(net45),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _724_ (.I(net45),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _725_ (.I(net45),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _726_ (.I(net45),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _727_ (.I(net45),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _728_ (.I(net45),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _729_ (.I(net26),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _730_ (.I(net26),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _731_ (.I(net26),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _732_ (.I(net26),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _733_ (.I(net26),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _734_ (.I(net26),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _735_ (.I(net26),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _736_ (.I(net26),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _737_ (.I(net26),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _738_ (.D(_090_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _739_ (.D(_091_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _740_ (.D(_092_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _741_ (.D(_093_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _742_ (.D(_094_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _743_ (.D(_095_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _744_ (.D(_096_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _745_ (.D(_097_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _746_ (.D(_098_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _747_ (.D(_099_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _748_ (.D(_001_),
    .SETN(_003_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _749_ (.D(\state[2] ),
    .RN(_004_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _750_ (.D(_000_),
    .RN(_005_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _751_ (.D(_002_),
    .RN(_006_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _752_ (.D(_100_),
    .RN(_007_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _753_ (.D(_101_),
    .RN(_008_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _754_ (.D(_102_),
    .RN(_009_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _755_ (.D(_103_),
    .RN(_010_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _756_ (.D(_104_),
    .RN(_011_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _757_ (.D(_105_),
    .RN(_012_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _758_ (.D(_106_),
    .RN(_013_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _759_ (.D(_107_),
    .RN(_014_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _760_ (.D(_108_),
    .RN(_015_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(sense_reg));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _761_ (.D(_109_),
    .RN(_016_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _762_ (.D(_110_),
    .RN(_017_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _763_ (.D(_111_),
    .RN(_018_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _764_ (.D(_112_),
    .RN(_019_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _765_ (.D(_113_),
    .RN(_020_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _766_ (.D(_114_),
    .RN(_021_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _767_ (.D(_115_),
    .RN(_022_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _768_ (.D(_116_),
    .RN(_023_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _769_ (.D(_117_),
    .RN(_024_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\bit_sel_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _770_ (.D(_118_),
    .RN(_025_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _771_ (.D(_119_),
    .RN(_026_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _772_ (.D(_120_),
    .RN(_027_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _773_ (.D(_121_),
    .RN(_028_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\bit_sel_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _774_ (.D(_122_),
    .RN(_029_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\bit_sel_reg[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _775_ (.D(_123_),
    .RN(_030_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _776_ (.D(_124_),
    .RN(_031_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _777_ (.D(_125_),
    .RN(_032_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _778_ (.D(_126_),
    .RN(_033_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _779_ (.D(_127_),
    .RN(_034_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _780_ (.D(_128_),
    .RN(_035_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _781_ (.D(_129_),
    .RN(_036_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _782_ (.D(_130_),
    .RN(_037_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _783_ (.D(_131_),
    .RN(_038_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _784_ (.D(_132_),
    .RN(_039_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _785_ (.D(_133_),
    .RN(_040_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _786_ (.D(_134_),
    .RN(_041_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _787_ (.D(_135_),
    .RN(_042_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _788_ (.D(_136_),
    .RN(_043_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _789_ (.D(_137_),
    .RN(_044_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\bit_sel_reg[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _790_ (.D(_138_),
    .RN(_045_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _791_ (.D(_139_),
    .RN(_046_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _792_ (.D(_140_),
    .RN(_047_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _793_ (.D(_141_),
    .RN(_048_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _794_ (.D(_142_),
    .RN(_049_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _795_ (.D(_143_),
    .RN(_050_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _796_ (.D(_144_),
    .RN(_051_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _797_ (.D(_145_),
    .RN(_052_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\bit_sel_reg[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _798_ (.D(_146_),
    .RN(_053_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _799_ (.D(_147_),
    .RN(_054_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _800_ (.D(_148_),
    .RN(_055_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _801_ (.D(_149_),
    .RN(_056_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _802_ (.D(_150_),
    .RN(_057_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _803_ (.D(_151_),
    .RN(_058_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _804_ (.D(_152_),
    .RN(_059_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _805_ (.D(_153_),
    .RN(_060_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\bit_sel_reg[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _806_ (.D(_154_),
    .RN(_061_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\bit_sel_reg[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _807_ (.D(_155_),
    .RN(_062_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _808_ (.D(_156_),
    .RN(_063_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _809_ (.D(_157_),
    .RN(_064_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\bit_sel_reg[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _810_ (.D(_158_),
    .RN(_065_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _811_ (.D(_159_),
    .RN(_066_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _812_ (.D(_160_),
    .RN(_067_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _813_ (.D(_161_),
    .RN(_068_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _814_ (.D(_162_),
    .RN(_069_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _815_ (.D(_163_),
    .RN(_070_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\bit_sel_reg[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _816_ (.D(_164_),
    .RN(_071_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\bit_sel_reg[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _817_ (.D(_165_),
    .RN(_072_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _818_ (.D(_166_),
    .RN(_073_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _819_ (.D(_167_),
    .RN(_074_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _820_ (.D(_168_),
    .RN(_075_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _821_ (.D(_169_),
    .RN(_076_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\bit_sel_reg[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _822_ (.D(_170_),
    .RN(_077_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _823_ (.D(_171_),
    .RN(_078_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\bit_sel_reg[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _824_ (.D(_172_),
    .RN(_079_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\bit_sel_reg[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _825_ (.D(_173_),
    .RN(_080_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\bit_sel_reg[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _826_ (.D(_174_),
    .SETN(_081_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\col_prog_n_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _827_ (.D(_175_),
    .SETN(_082_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\col_prog_n_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _828_ (.D(_176_),
    .SETN(_083_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\col_prog_n_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _829_ (.D(_177_),
    .SETN(_084_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\col_prog_n_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _830_ (.D(_178_),
    .SETN(_085_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\col_prog_n_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _831_ (.D(_179_),
    .SETN(_086_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\col_prog_n_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _832_ (.D(_180_),
    .SETN(_087_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\col_prog_n_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _833_ (.D(_181_),
    .SETN(_088_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\col_prog_n_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _834_ (.D(_182_),
    .SETN(_089_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(preset_n_reg));
 efuse_array_64x8 efuse_array (.PRESET_N(preset_n),
    .SENSE(sense),
    .BIT_SEL({\bit_sel[63] ,
    \bit_sel[62] ,
    \bit_sel[61] ,
    \bit_sel[60] ,
    \bit_sel[59] ,
    \bit_sel[58] ,
    \bit_sel[57] ,
    \bit_sel[56] ,
    \bit_sel[55] ,
    \bit_sel[54] ,
    \bit_sel[53] ,
    \bit_sel[52] ,
    \bit_sel[51] ,
    \bit_sel[50] ,
    \bit_sel[49] ,
    \bit_sel[48] ,
    \bit_sel[47] ,
    \bit_sel[46] ,
    \bit_sel[45] ,
    \bit_sel[44] ,
    \bit_sel[43] ,
    \bit_sel[42] ,
    \bit_sel[41] ,
    \bit_sel[40] ,
    \bit_sel[39] ,
    \bit_sel[38] ,
    \bit_sel[37] ,
    \bit_sel[36] ,
    \bit_sel[35] ,
    \bit_sel[34] ,
    \bit_sel[33] ,
    \bit_sel[32] ,
    \bit_sel[31] ,
    \bit_sel[30] ,
    \bit_sel[29] ,
    \bit_sel[28] ,
    \bit_sel[27] ,
    \bit_sel[26] ,
    \bit_sel[25] ,
    \bit_sel[24] ,
    \bit_sel[23] ,
    \bit_sel[22] ,
    \bit_sel[21] ,
    \bit_sel[20] ,
    \bit_sel[19] ,
    \bit_sel[18] ,
    \bit_sel[17] ,
    \bit_sel[16] ,
    \bit_sel[15] ,
    \bit_sel[14] ,
    \bit_sel[13] ,
    \bit_sel[12] ,
    \bit_sel[11] ,
    \bit_sel[10] ,
    \bit_sel[9] ,
    \bit_sel[8] ,
    \bit_sel[7] ,
    \bit_sel[6] ,
    \bit_sel[5] ,
    \bit_sel[4] ,
    \bit_sel[3] ,
    \bit_sel[2] ,
    \bit_sel[1] ,
    \bit_sel[0] }),
    .COL_PROG_N({\col_prog_n[7] ,
    \col_prog_n[6] ,
    \col_prog_n[5] ,
    \col_prog_n[4] ,
    \col_prog_n[3] ,
    \col_prog_n[2] ,
    \col_prog_n[1] ,
    \col_prog_n[0] }),
    .OUT({\efuse_out[7] ,
    \efuse_out[6] ,
    \efuse_out[5] ,
    \efuse_out[4] ,
    \efuse_out[3] ,
    \efuse_out[2] ,
    \efuse_out[1] ,
    \efuse_out[0] }));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 \genblk1[0].prog_or_keep_cell  (.A1(\col_prog_n_reg[0] ),
    .A2(write_disable_i),
    .Z(\col_prog_n[0] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 \genblk1[1].prog_or_keep_cell  (.A1(\col_prog_n_reg[1] ),
    .A2(write_disable_i),
    .Z(\col_prog_n[1] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 \genblk1[2].prog_or_keep_cell  (.A1(\col_prog_n_reg[2] ),
    .A2(write_disable_i),
    .Z(\col_prog_n[2] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 \genblk1[3].prog_or_keep_cell  (.A1(\col_prog_n_reg[3] ),
    .A2(write_disable_i),
    .Z(\col_prog_n[3] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 \genblk1[4].prog_or_keep_cell  (.A1(\col_prog_n_reg[4] ),
    .A2(write_disable_i),
    .Z(\col_prog_n[4] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 \genblk1[5].prog_or_keep_cell  (.A1(\col_prog_n_reg[5] ),
    .A2(write_disable_i),
    .Z(\col_prog_n[5] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 \genblk1[6].prog_or_keep_cell  (.A1(\col_prog_n_reg[6] ),
    .A2(write_disable_i),
    .Z(\col_prog_n[6] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 \genblk1[7].prog_or_keep_cell  (.A1(\col_prog_n_reg[7] ),
    .A2(write_disable_i),
    .Z(\col_prog_n[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[0].bitsel_buf_keep_cell  (.I(\bit_sel_reg[0] ),
    .Z(\bit_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[10].bitsel_buf_keep_cell  (.I(\bit_sel_reg[10] ),
    .Z(\bit_sel[10] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[11].bitsel_buf_keep_cell  (.I(\bit_sel_reg[11] ),
    .Z(\bit_sel[11] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[12].bitsel_buf_keep_cell  (.I(\bit_sel_reg[12] ),
    .Z(\bit_sel[12] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[13].bitsel_buf_keep_cell  (.I(\bit_sel_reg[13] ),
    .Z(\bit_sel[13] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[14].bitsel_buf_keep_cell  (.I(\bit_sel_reg[14] ),
    .Z(\bit_sel[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[15].bitsel_buf_keep_cell  (.I(\bit_sel_reg[15] ),
    .Z(\bit_sel[15] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[16].bitsel_buf_keep_cell  (.I(\bit_sel_reg[16] ),
    .Z(\bit_sel[16] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[17].bitsel_buf_keep_cell  (.I(\bit_sel_reg[17] ),
    .Z(\bit_sel[17] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[18].bitsel_buf_keep_cell  (.I(\bit_sel_reg[18] ),
    .Z(\bit_sel[18] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[19].bitsel_buf_keep_cell  (.I(\bit_sel_reg[19] ),
    .Z(\bit_sel[19] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[1].bitsel_buf_keep_cell  (.I(\bit_sel_reg[1] ),
    .Z(\bit_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[20].bitsel_buf_keep_cell  (.I(\bit_sel_reg[20] ),
    .Z(\bit_sel[20] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[21].bitsel_buf_keep_cell  (.I(\bit_sel_reg[21] ),
    .Z(\bit_sel[21] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[22].bitsel_buf_keep_cell  (.I(\bit_sel_reg[22] ),
    .Z(\bit_sel[22] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[23].bitsel_buf_keep_cell  (.I(\bit_sel_reg[23] ),
    .Z(\bit_sel[23] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[24].bitsel_buf_keep_cell  (.I(\bit_sel_reg[24] ),
    .Z(\bit_sel[24] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[25].bitsel_buf_keep_cell  (.I(\bit_sel_reg[25] ),
    .Z(\bit_sel[25] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[26].bitsel_buf_keep_cell  (.I(\bit_sel_reg[26] ),
    .Z(\bit_sel[26] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[27].bitsel_buf_keep_cell  (.I(\bit_sel_reg[27] ),
    .Z(\bit_sel[27] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[28].bitsel_buf_keep_cell  (.I(\bit_sel_reg[28] ),
    .Z(\bit_sel[28] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[29].bitsel_buf_keep_cell  (.I(\bit_sel_reg[29] ),
    .Z(\bit_sel[29] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[2].bitsel_buf_keep_cell  (.I(\bit_sel_reg[2] ),
    .Z(\bit_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[30].bitsel_buf_keep_cell  (.I(\bit_sel_reg[30] ),
    .Z(\bit_sel[30] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[31].bitsel_buf_keep_cell  (.I(\bit_sel_reg[31] ),
    .Z(\bit_sel[31] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[32].bitsel_buf_keep_cell  (.I(\bit_sel_reg[32] ),
    .Z(\bit_sel[32] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[33].bitsel_buf_keep_cell  (.I(\bit_sel_reg[33] ),
    .Z(\bit_sel[33] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[34].bitsel_buf_keep_cell  (.I(\bit_sel_reg[34] ),
    .Z(\bit_sel[34] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[35].bitsel_buf_keep_cell  (.I(\bit_sel_reg[35] ),
    .Z(\bit_sel[35] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[36].bitsel_buf_keep_cell  (.I(\bit_sel_reg[36] ),
    .Z(\bit_sel[36] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[37].bitsel_buf_keep_cell  (.I(\bit_sel_reg[37] ),
    .Z(\bit_sel[37] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[38].bitsel_buf_keep_cell  (.I(\bit_sel_reg[38] ),
    .Z(\bit_sel[38] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[39].bitsel_buf_keep_cell  (.I(\bit_sel_reg[39] ),
    .Z(\bit_sel[39] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[3].bitsel_buf_keep_cell  (.I(\bit_sel_reg[3] ),
    .Z(\bit_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[40].bitsel_buf_keep_cell  (.I(\bit_sel_reg[40] ),
    .Z(\bit_sel[40] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[41].bitsel_buf_keep_cell  (.I(\bit_sel_reg[41] ),
    .Z(\bit_sel[41] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[42].bitsel_buf_keep_cell  (.I(\bit_sel_reg[42] ),
    .Z(\bit_sel[42] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[43].bitsel_buf_keep_cell  (.I(\bit_sel_reg[43] ),
    .Z(\bit_sel[43] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[44].bitsel_buf_keep_cell  (.I(\bit_sel_reg[44] ),
    .Z(\bit_sel[44] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[45].bitsel_buf_keep_cell  (.I(\bit_sel_reg[45] ),
    .Z(\bit_sel[45] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[46].bitsel_buf_keep_cell  (.I(\bit_sel_reg[46] ),
    .Z(\bit_sel[46] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[47].bitsel_buf_keep_cell  (.I(\bit_sel_reg[47] ),
    .Z(\bit_sel[47] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[48].bitsel_buf_keep_cell  (.I(\bit_sel_reg[48] ),
    .Z(\bit_sel[48] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[49].bitsel_buf_keep_cell  (.I(\bit_sel_reg[49] ),
    .Z(\bit_sel[49] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[4].bitsel_buf_keep_cell  (.I(\bit_sel_reg[4] ),
    .Z(\bit_sel[4] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[50].bitsel_buf_keep_cell  (.I(\bit_sel_reg[50] ),
    .Z(\bit_sel[50] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[51].bitsel_buf_keep_cell  (.I(\bit_sel_reg[51] ),
    .Z(\bit_sel[51] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[52].bitsel_buf_keep_cell  (.I(\bit_sel_reg[52] ),
    .Z(\bit_sel[52] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[53].bitsel_buf_keep_cell  (.I(\bit_sel_reg[53] ),
    .Z(\bit_sel[53] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[54].bitsel_buf_keep_cell  (.I(\bit_sel_reg[54] ),
    .Z(\bit_sel[54] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[55].bitsel_buf_keep_cell  (.I(\bit_sel_reg[55] ),
    .Z(\bit_sel[55] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[56].bitsel_buf_keep_cell  (.I(\bit_sel_reg[56] ),
    .Z(\bit_sel[56] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[57].bitsel_buf_keep_cell  (.I(\bit_sel_reg[57] ),
    .Z(\bit_sel[57] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[58].bitsel_buf_keep_cell  (.I(\bit_sel_reg[58] ),
    .Z(\bit_sel[58] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[59].bitsel_buf_keep_cell  (.I(\bit_sel_reg[59] ),
    .Z(\bit_sel[59] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[5].bitsel_buf_keep_cell  (.I(\bit_sel_reg[5] ),
    .Z(\bit_sel[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[60].bitsel_buf_keep_cell  (.I(\bit_sel_reg[60] ),
    .Z(\bit_sel[60] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[61].bitsel_buf_keep_cell  (.I(\bit_sel_reg[61] ),
    .Z(\bit_sel[61] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[62].bitsel_buf_keep_cell  (.I(\bit_sel_reg[62] ),
    .Z(\bit_sel[62] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[63].bitsel_buf_keep_cell  (.I(\bit_sel_reg[63] ),
    .Z(\bit_sel[63] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[6].bitsel_buf_keep_cell  (.I(\bit_sel_reg[6] ),
    .Z(\bit_sel[6] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[7].bitsel_buf_keep_cell  (.I(\bit_sel_reg[7] ),
    .Z(\bit_sel[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[8].bitsel_buf_keep_cell  (.I(\bit_sel_reg[8] ),
    .Z(\bit_sel[8] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \genblk2[9].bitsel_buf_keep_cell  (.I(\bit_sel_reg[9] ),
    .Z(\bit_sel[9] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 preset_buf_keep_cell (.I(preset_n_reg),
    .Z(preset_n));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 sense_buf_keep_cell (.I(sense_reg),
    .Z(sense));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_1_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_1_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_1_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_1_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_1_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_1_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_1_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_1_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_1_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_1_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_1_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_1_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_1_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_1_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_1_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_1_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_1_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_1_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_1_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_1_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_1_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_1_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_1_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_1_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_1_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_1_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_1_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_1_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_1_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_1_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_1_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_1_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_1_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_1_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_1_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_1_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_1_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_1_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_1_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_1_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_1_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_1_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_1_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_1_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_1_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_1_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_1_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_1_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_1_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_1_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_1_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_1_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_1_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_1_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_1_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_1_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_1_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_1_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_1_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_1_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_1_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_1_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_1_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_1_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_1_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_1_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_1_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_1_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_1_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_1_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_1_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_1_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_1_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_1_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_1_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_1_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_1_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_1_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_1_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_1_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_1_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_1_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_1_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_1_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_1_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_1_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_1_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_1_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_1_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_1_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_1_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_1_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_1_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_1_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_1_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_1_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_1_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_1_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_1_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_1_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_1_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_1_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_1_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_1_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_1_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_1_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_1_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_1_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_1_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_1_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_1_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_1_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_1_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_1_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_1_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_1_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_1_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_1_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_1_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_1_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_1_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_1_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_1_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_1_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_1_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_1_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_1_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_1_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_1_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_1_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_1_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_1_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_1_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_1_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_1_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_1_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_1_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_1_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_1_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_1_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_1_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_1_Left_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_1_Left_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_1_Left_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_1_Left_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_1_Left_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_1_Left_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_1_Left_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_1_Left_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_1_Left_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_1_Left_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_1_Left_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_1_Left_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_1_Left_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_1_Left_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_1_Left_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_1_Left_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_1_Left_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_1_Left_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_1_Left_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_1_Left_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_1_Left_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_1_Left_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_1_Left_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_1_Left_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Right_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Right_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Right_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Right_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Right_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Right_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Right_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Right_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Right_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Right_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Right_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Right_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Right_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Right_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Right_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Right_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Right_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Right_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Right_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Right_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Right_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Right_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Right_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Right_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Right_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Right_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Right_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Right_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Right_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Right_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Right_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Right_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Right_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Right_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Right_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Right_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Right_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Right_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Right_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Right_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Right_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Right_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Right_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Right_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Right_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Right_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Right_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Right_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Right_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Right_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Right_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Right_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Right_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Right_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Right_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Right_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Right_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Right_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Right_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Right_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Right_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Right_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Right_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Right_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Right_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Right_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Right_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Right_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Right_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Right_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Right_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Right_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Right_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Right_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Right_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Right_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Right_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Right_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Right_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_2_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_2_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_2_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_2_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_2_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_2_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_2_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_2_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_2_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_2_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_2_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_2_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_2_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_2_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_2_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_2_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_2_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_2_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_2_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_2_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_2_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_2_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_2_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_2_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_2_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_2_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_2_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_2_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_2_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_2_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_2_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_2_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_2_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_2_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_2_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_2_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_2_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_2_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_2_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_2_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_2_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_2_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_2_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_2_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_2_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_2_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_2_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_2_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_2_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_2_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_2_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_2_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_2_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_2_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_2_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_2_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_2_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_2_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_2_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_2_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_2_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_2_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_2_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_2_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_2_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_2_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_2_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_2_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_2_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_2_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_2_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_2_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_2_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_2_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_2_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_2_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_2_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_2_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_2_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_2_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_2_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_2_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_2_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_1_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_1_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_1_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_1_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_1_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_1_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_1_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_1_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_1_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_1_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_1_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_1_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_1_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_1_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_1_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_1_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_1_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_1_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_1_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_1_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_1_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_1_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_1_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_1_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_1_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_1_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_1_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_1_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_1_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_1_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_1_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_1_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(wb_adr_i[0]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(wb_adr_i[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(wb_adr_i[2]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(wb_adr_i[3]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(wb_adr_i[4]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(wb_adr_i[5]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(wb_cyc_i),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input18 (.I(wb_dat_i[0]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(wb_dat_i[1]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(wb_dat_i[2]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input21 (.I(wb_dat_i[3]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input22 (.I(wb_dat_i[4]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input23 (.I(wb_dat_i[5]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input24 (.I(wb_dat_i[6]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(wb_dat_i[7]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input26 (.I(wb_rst_i),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input27 (.I(wb_stb_i),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(wb_we_i),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output29 (.I(net29),
    .Z(wb_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output30 (.I(net30),
    .Z(wb_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output31 (.I(net31),
    .Z(wb_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output32 (.I(net32),
    .Z(wb_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output33 (.I(net33),
    .Z(wb_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output34 (.I(net34),
    .Z(wb_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output35 (.I(net35),
    .Z(wb_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output36 (.I(net36),
    .Z(wb_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 output37 (.I(net37),
    .Z(wb_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap38 (.I(net39),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap39 (.I(_305_),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap40 (.I(net41),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 max_cap41 (.I(_224_),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap42 (.I(net43),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 wire43 (.I(_215_),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_12 max_cap44 (.I(net45),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 load_slew45 (.I(net26),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload0 (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload1 (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload2 (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload3 (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 clkload4 (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload5 (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 clkload6 (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_388 ();
endmodule
