VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_array_16x1
  CLASS BLOCK ;
  FOREIGN efuse_array_16x1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 44.480 BY 40.130 ;
  PIN COL_PROG_N[0]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 39.440 39.430 43.000 39.730 ;
    END
  END COL_PROG_N[0]
  PIN PRESET_N
    ANTENNAGATEAREA 1.220000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.010 19.885 1.290 40.130 ;
        RECT 1.010 19.505 1.370 19.885 ;
        RECT 1.010 0.000 1.290 19.505 ;
    END
  END PRESET_N
  PIN SENSE
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER Metal2 ;
        RECT 1.655 18.700 1.935 40.130 ;
        RECT 1.655 18.320 3.080 18.700 ;
        RECT 1.655 0.000 1.935 18.320 ;
    END
  END SENSE
  PIN OUT[0]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 2.300 11.030 2.680 11.410 ;
    END
  END OUT[0]
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 6.700 0.000 9.560 40.130 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3.710 0.000 4.710 40.130 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 0.070 0.000 1.070 40.130 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 39.990 0.000 44.240 40.130 ;
    END
  END VDD
  PIN BIT_SEL[0]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 37.740 24.225 38.020 39.505 ;
        RECT 37.700 23.845 38.080 24.225 ;
        RECT 37.740 0.000 38.020 23.845 ;
    END
  END BIT_SEL[0]
  PIN BIT_SEL[1]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 37.100 15.660 37.380 39.505 ;
        RECT 37.060 15.280 37.440 15.660 ;
        RECT 37.100 0.000 37.380 15.280 ;
    END
  END BIT_SEL[1]
  PIN BIT_SEL[2]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 36.460 26.065 36.740 39.505 ;
        RECT 36.420 25.685 36.800 26.065 ;
        RECT 36.460 0.000 36.740 25.685 ;
    END
  END BIT_SEL[2]
  PIN BIT_SEL[3]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 35.820 13.820 36.100 39.505 ;
        RECT 35.780 13.440 36.160 13.820 ;
        RECT 35.820 0.000 36.100 13.440 ;
    END
  END BIT_SEL[3]
  PIN BIT_SEL[4]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 35.180 27.905 35.460 39.505 ;
        RECT 35.140 27.525 35.520 27.905 ;
        RECT 35.180 0.000 35.460 27.525 ;
    END
  END BIT_SEL[4]
  PIN BIT_SEL[5]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 34.540 11.975 34.820 39.505 ;
        RECT 34.500 11.595 34.880 11.975 ;
        RECT 34.540 0.000 34.820 11.595 ;
    END
  END BIT_SEL[5]
  PIN BIT_SEL[6]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 33.900 30.550 34.180 39.505 ;
        RECT 33.860 30.170 34.240 30.550 ;
        RECT 33.900 0.000 34.180 30.170 ;
    END
  END BIT_SEL[6]
  PIN BIT_SEL[7]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 33.260 9.335 33.540 39.505 ;
        RECT 33.220 8.955 33.600 9.335 ;
        RECT 33.260 0.000 33.540 8.955 ;
    END
  END BIT_SEL[7]
  PIN BIT_SEL[8]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 32.620 32.390 32.900 39.505 ;
        RECT 32.580 32.010 32.960 32.390 ;
        RECT 32.620 0.000 32.900 32.010 ;
    END
  END BIT_SEL[8]
  PIN BIT_SEL[9]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 31.980 7.495 32.260 39.505 ;
        RECT 31.940 7.115 32.320 7.495 ;
        RECT 31.980 0.000 32.260 7.115 ;
    END
  END BIT_SEL[9]
  PIN BIT_SEL[10]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 31.340 34.230 31.620 39.505 ;
        RECT 31.300 33.850 31.680 34.230 ;
        RECT 31.340 0.000 31.620 33.850 ;
    END
  END BIT_SEL[10]
  PIN BIT_SEL[11]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 30.700 5.650 30.980 39.505 ;
        RECT 30.660 5.270 31.040 5.650 ;
        RECT 30.700 0.000 30.980 5.270 ;
    END
  END BIT_SEL[11]
  PIN BIT_SEL[12]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 30.060 36.875 30.340 39.505 ;
        RECT 30.020 36.495 30.400 36.875 ;
        RECT 30.060 0.000 30.340 36.495 ;
    END
  END BIT_SEL[12]
  PIN BIT_SEL[13]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 29.420 3.010 29.700 39.505 ;
        RECT 29.380 2.630 29.760 3.010 ;
        RECT 29.420 0.000 29.700 2.630 ;
    END
  END BIT_SEL[13]
  PIN BIT_SEL[14]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 28.780 38.715 29.060 39.505 ;
        RECT 28.740 38.335 29.120 38.715 ;
        RECT 28.780 0.000 29.060 38.335 ;
    END
  END BIT_SEL[14]
  PIN BIT_SEL[15]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 28.140 1.170 28.420 39.505 ;
        RECT 28.100 0.790 28.480 1.170 ;
        RECT 28.140 0.000 28.420 0.790 ;
    END
  END BIT_SEL[15]
  OBS
      LAYER Metal1 ;
        RECT 0.130 39.220 0.730 40.130 ;
        RECT 4.050 39.220 4.650 40.130 ;
        RECT 0.130 38.880 2.430 39.220 ;
        RECT 3.160 38.880 4.650 39.220 ;
        RECT 6.690 38.895 37.210 39.275 ;
        RECT 0.130 38.265 0.730 38.880 ;
        RECT 0.130 38.035 1.860 38.265 ;
        RECT 2.160 38.035 3.820 38.265 ;
        RECT 0.130 36.025 0.730 38.035 ;
        RECT 2.160 37.000 2.390 38.035 ;
        RECT 2.795 36.745 3.025 37.790 ;
        RECT 4.050 36.745 4.650 38.880 ;
        RECT 5.840 38.640 6.460 38.825 ;
        RECT 37.440 38.640 38.060 38.825 ;
        RECT 5.840 38.410 38.060 38.640 ;
        RECT 5.840 38.225 6.460 38.410 ;
        RECT 37.440 38.225 38.060 38.410 ;
        RECT 33.440 38.145 35.060 38.155 ;
        RECT 6.690 37.775 37.210 38.145 ;
        RECT 6.690 37.055 37.210 37.435 ;
        RECT 0.960 36.515 3.025 36.745 ;
        RECT 3.255 36.515 4.650 36.745 ;
        RECT 0.130 35.795 1.860 36.025 ;
        RECT 2.160 35.795 3.820 36.025 ;
        RECT 0.130 33.785 0.730 35.795 ;
        RECT 2.160 34.760 2.390 35.795 ;
        RECT 2.795 34.505 3.025 35.550 ;
        RECT 4.050 34.505 4.650 36.515 ;
        RECT 5.840 36.800 6.460 36.985 ;
        RECT 37.440 36.800 38.060 36.985 ;
        RECT 5.840 36.570 38.060 36.800 ;
        RECT 5.840 36.385 6.460 36.570 ;
        RECT 37.440 36.385 38.060 36.570 ;
        RECT 29.600 36.305 31.220 36.315 ;
        RECT 6.690 35.935 37.210 36.305 ;
        RECT 6.700 35.140 37.200 35.580 ;
        RECT 0.960 34.275 3.025 34.505 ;
        RECT 3.255 34.275 4.650 34.505 ;
        RECT 6.690 34.410 37.210 34.790 ;
        RECT 0.130 33.555 1.860 33.785 ;
        RECT 2.160 33.555 3.820 33.785 ;
        RECT 0.130 31.545 0.730 33.555 ;
        RECT 2.160 32.520 2.390 33.555 ;
        RECT 2.795 32.265 3.025 33.310 ;
        RECT 4.050 32.265 4.650 34.275 ;
        RECT 5.840 34.155 6.460 34.340 ;
        RECT 37.440 34.155 38.060 34.340 ;
        RECT 5.840 33.925 38.060 34.155 ;
        RECT 5.840 33.740 6.460 33.925 ;
        RECT 37.440 33.740 38.060 33.925 ;
        RECT 25.760 33.660 27.380 33.670 ;
        RECT 6.690 33.290 37.210 33.660 ;
        RECT 6.690 32.570 37.210 32.950 ;
        RECT 0.960 32.035 3.025 32.265 ;
        RECT 3.255 32.035 4.650 32.265 ;
        RECT 0.130 31.315 1.860 31.545 ;
        RECT 2.160 31.315 3.820 31.545 ;
        RECT 0.130 29.305 0.730 31.315 ;
        RECT 2.160 30.280 2.390 31.315 ;
        RECT 2.795 30.025 3.025 31.070 ;
        RECT 4.050 30.025 4.650 32.035 ;
        RECT 5.840 32.315 6.460 32.500 ;
        RECT 37.440 32.315 38.060 32.500 ;
        RECT 5.840 32.085 38.060 32.315 ;
        RECT 5.840 31.900 6.460 32.085 ;
        RECT 37.440 31.900 38.060 32.085 ;
        RECT 21.920 31.820 23.540 31.830 ;
        RECT 6.690 31.450 37.210 31.820 ;
        RECT 6.690 30.730 37.210 31.110 ;
        RECT 5.840 30.475 6.460 30.660 ;
        RECT 37.440 30.475 38.060 30.660 ;
        RECT 5.840 30.245 38.060 30.475 ;
        RECT 5.840 30.060 6.460 30.245 ;
        RECT 37.440 30.060 38.060 30.245 ;
        RECT 0.960 29.795 3.025 30.025 ;
        RECT 3.255 29.795 4.650 30.025 ;
        RECT 18.080 29.980 19.700 29.990 ;
        RECT 0.130 29.075 1.860 29.305 ;
        RECT 2.160 29.075 3.820 29.305 ;
        RECT 0.130 26.920 0.730 29.075 ;
        RECT 2.160 28.040 2.390 29.075 ;
        RECT 2.795 27.785 3.025 28.830 ;
        RECT 4.050 27.785 4.650 29.795 ;
        RECT 6.690 29.610 37.210 29.980 ;
        RECT 6.700 28.815 37.200 29.255 ;
        RECT 6.690 28.085 37.210 28.465 ;
        RECT 0.960 27.555 3.025 27.785 ;
        RECT 3.255 27.555 4.650 27.785 ;
        RECT 4.050 26.920 4.650 27.555 ;
        RECT 5.840 27.830 6.460 28.015 ;
        RECT 37.440 27.830 38.060 28.015 ;
        RECT 5.840 27.600 38.060 27.830 ;
        RECT 5.840 27.415 6.460 27.600 ;
        RECT 37.440 27.415 38.060 27.600 ;
        RECT 14.240 27.335 15.860 27.345 ;
        RECT 6.690 26.965 37.210 27.335 ;
        RECT 0.130 26.580 2.420 26.920 ;
        RECT 3.165 26.580 4.650 26.920 ;
        RECT 0.130 25.945 0.730 26.580 ;
        RECT 0.130 25.715 1.860 25.945 ;
        RECT 2.160 25.715 3.820 25.945 ;
        RECT 0.130 23.705 0.730 25.715 ;
        RECT 2.160 24.680 2.390 25.715 ;
        RECT 2.795 24.425 3.025 25.470 ;
        RECT 4.050 24.425 4.650 26.580 ;
        RECT 6.690 26.245 37.210 26.625 ;
        RECT 5.840 25.990 6.460 26.175 ;
        RECT 37.440 25.990 38.060 26.175 ;
        RECT 5.840 25.760 38.060 25.990 ;
        RECT 5.840 25.575 6.460 25.760 ;
        RECT 37.440 25.575 38.060 25.760 ;
        RECT 10.400 25.495 12.020 25.505 ;
        RECT 6.690 25.125 37.210 25.495 ;
        RECT 0.960 24.195 3.025 24.425 ;
        RECT 3.255 24.195 4.650 24.425 ;
        RECT 6.690 24.405 37.210 24.785 ;
        RECT 0.130 23.475 1.860 23.705 ;
        RECT 2.160 23.475 3.820 23.705 ;
        RECT 0.130 21.320 0.730 23.475 ;
        RECT 2.160 22.440 2.390 23.475 ;
        RECT 2.795 22.185 3.025 23.230 ;
        RECT 4.050 22.185 4.650 24.195 ;
        RECT 5.840 24.150 6.460 24.335 ;
        RECT 37.440 24.150 38.060 24.335 ;
        RECT 5.840 23.920 38.060 24.150 ;
        RECT 5.840 23.735 6.460 23.920 ;
        RECT 37.440 23.735 38.060 23.920 ;
        RECT 6.690 23.285 37.210 23.655 ;
        RECT 0.960 21.955 3.025 22.185 ;
        RECT 3.255 21.955 4.650 22.185 ;
        RECT 4.050 21.320 4.650 21.955 ;
        RECT 0.130 20.980 2.420 21.320 ;
        RECT 3.165 20.980 4.650 21.320 ;
        RECT 0.130 20.345 0.730 20.980 ;
        RECT 0.130 20.115 1.710 20.345 ;
        RECT 0.130 18.075 0.730 20.115 ;
        RECT 2.140 19.885 2.500 19.970 ;
        RECT 1.010 19.655 2.500 19.885 ;
        RECT 1.010 19.505 1.370 19.655 ;
        RECT 0.960 18.870 1.910 19.275 ;
        RECT 0.130 17.845 1.420 18.075 ;
        RECT 0.130 16.885 0.730 17.845 ;
        RECT 1.650 17.525 1.910 18.870 ;
        RECT 2.140 18.220 2.500 19.655 ;
        RECT 2.730 18.320 3.080 19.520 ;
        RECT 3.440 18.910 3.820 20.555 ;
        RECT 2.520 17.525 2.870 17.585 ;
        RECT 3.440 17.525 3.780 18.130 ;
        RECT 1.650 17.265 3.780 17.525 ;
        RECT 2.520 17.205 2.870 17.265 ;
        RECT 4.050 16.985 4.650 20.980 ;
        RECT 6.495 20.500 8.245 23.285 ;
        RECT 8.885 20.500 9.695 21.500 ;
        RECT 10.335 20.500 12.085 22.795 ;
        RECT 12.725 20.500 13.535 21.500 ;
        RECT 14.175 20.500 15.925 22.795 ;
        RECT 16.565 20.500 17.375 21.500 ;
        RECT 18.015 20.500 19.765 22.795 ;
        RECT 20.405 20.500 21.215 21.500 ;
        RECT 21.855 20.500 23.605 22.795 ;
        RECT 24.245 20.500 25.055 21.500 ;
        RECT 25.695 20.500 27.445 22.795 ;
        RECT 28.085 20.500 28.895 21.500 ;
        RECT 29.535 20.500 31.285 22.795 ;
        RECT 31.925 20.500 32.735 21.500 ;
        RECT 33.375 20.500 35.125 22.795 ;
        RECT 35.765 20.500 36.575 21.500 ;
        RECT 38.990 20.690 39.360 39.200 ;
        RECT 40.010 35.565 40.380 39.200 ;
        RECT 40.005 35.185 40.385 35.565 ;
        RECT 40.010 32.565 40.380 35.185 ;
        RECT 40.005 32.185 40.385 32.565 ;
        RECT 40.010 29.565 40.380 32.185 ;
        RECT 40.005 29.185 40.385 29.565 ;
        RECT 40.010 26.565 40.380 29.185 ;
        RECT 40.005 26.185 40.385 26.565 ;
        RECT 40.010 23.565 40.380 26.185 ;
        RECT 40.005 23.185 40.385 23.565 ;
        RECT 38.990 20.310 39.370 20.690 ;
        RECT 38.990 19.240 39.360 20.310 ;
        RECT 6.965 18.050 7.775 19.050 ;
        RECT 0.130 16.655 1.820 16.885 ;
        RECT 3.190 16.755 4.650 16.985 ;
        RECT 0.130 14.645 0.730 16.655 ;
        RECT 2.150 16.195 3.150 16.520 ;
        RECT 0.960 15.635 3.820 15.965 ;
        RECT 0.130 14.415 1.820 14.645 ;
        RECT 0.130 12.405 0.730 14.415 ;
        RECT 2.535 14.280 2.800 15.635 ;
        RECT 4.050 14.745 4.650 16.755 ;
        RECT 8.415 16.220 10.165 19.050 ;
        RECT 10.805 18.050 11.615 19.050 ;
        RECT 12.255 16.755 14.005 19.050 ;
        RECT 14.645 18.050 15.455 19.050 ;
        RECT 16.095 16.755 17.845 19.050 ;
        RECT 18.485 18.050 19.295 19.050 ;
        RECT 19.935 16.755 21.685 19.050 ;
        RECT 22.325 18.050 23.135 19.050 ;
        RECT 23.775 16.755 25.525 19.050 ;
        RECT 26.165 18.050 26.975 19.050 ;
        RECT 27.615 16.755 29.365 19.050 ;
        RECT 30.005 18.050 30.815 19.050 ;
        RECT 31.455 16.755 33.205 19.050 ;
        RECT 33.845 18.050 34.655 19.050 ;
        RECT 35.295 16.755 37.045 19.050 ;
        RECT 38.990 18.860 39.370 19.240 ;
        RECT 6.690 15.850 37.210 16.220 ;
        RECT 5.840 15.585 6.460 15.770 ;
        RECT 37.440 15.585 38.060 15.770 ;
        RECT 5.840 15.355 38.060 15.585 ;
        RECT 5.840 15.170 6.460 15.355 ;
        RECT 37.440 15.170 38.060 15.355 ;
        RECT 3.190 14.515 4.650 14.745 ;
        RECT 6.690 14.720 37.210 15.100 ;
        RECT 2.150 13.955 3.150 14.280 ;
        RECT 0.960 13.395 3.820 13.725 ;
        RECT 4.050 12.505 4.650 14.515 ;
        RECT 6.690 14.010 37.210 14.380 ;
        RECT 12.320 14.000 13.940 14.010 ;
        RECT 5.840 13.745 6.460 13.930 ;
        RECT 37.440 13.745 38.060 13.930 ;
        RECT 5.840 13.515 38.060 13.745 ;
        RECT 5.840 13.330 6.460 13.515 ;
        RECT 37.440 13.330 38.060 13.515 ;
        RECT 6.690 12.880 37.210 13.260 ;
        RECT 0.130 12.175 1.820 12.405 ;
        RECT 3.190 12.275 4.650 12.505 ;
        RECT 0.130 10.120 0.730 12.175 ;
        RECT 2.150 11.715 3.150 12.040 ;
        RECT 0.960 11.155 3.820 11.485 ;
        RECT 2.300 11.030 2.680 11.155 ;
        RECT 4.050 10.120 4.650 12.275 ;
        RECT 6.690 12.165 37.210 12.535 ;
        RECT 16.160 12.155 17.780 12.165 ;
        RECT 5.840 11.900 6.460 12.085 ;
        RECT 37.440 11.900 38.060 12.085 ;
        RECT 5.840 11.670 38.060 11.900 ;
        RECT 5.840 11.485 6.460 11.670 ;
        RECT 37.440 11.485 38.060 11.670 ;
        RECT 6.690 11.035 37.210 11.415 ;
        RECT 6.700 10.245 37.200 10.685 ;
        RECT 0.130 9.780 2.420 10.120 ;
        RECT 3.165 9.780 4.650 10.120 ;
        RECT 0.130 9.000 0.730 9.780 ;
        RECT 4.050 9.000 4.650 9.780 ;
        RECT 6.690 9.525 37.210 9.895 ;
        RECT 20.000 9.515 21.620 9.525 ;
        RECT 0.130 8.660 2.420 9.000 ;
        RECT 3.165 8.660 4.650 9.000 ;
        RECT 5.840 9.260 6.460 9.445 ;
        RECT 37.440 9.260 38.060 9.445 ;
        RECT 5.840 9.030 38.060 9.260 ;
        RECT 5.840 8.845 6.460 9.030 ;
        RECT 37.440 8.845 38.060 9.030 ;
        RECT 0.130 8.025 0.730 8.660 ;
        RECT 0.130 7.795 1.860 8.025 ;
        RECT 2.160 7.795 3.820 8.025 ;
        RECT 0.130 5.785 0.730 7.795 ;
        RECT 2.160 6.760 2.390 7.795 ;
        RECT 2.795 6.505 3.025 7.550 ;
        RECT 4.050 6.505 4.650 8.660 ;
        RECT 6.690 8.395 37.210 8.775 ;
        RECT 6.690 7.685 37.210 8.055 ;
        RECT 23.840 7.675 25.460 7.685 ;
        RECT 5.840 7.420 6.460 7.605 ;
        RECT 37.440 7.420 38.060 7.605 ;
        RECT 5.840 7.190 38.060 7.420 ;
        RECT 5.840 7.005 6.460 7.190 ;
        RECT 37.440 7.005 38.060 7.190 ;
        RECT 6.690 6.555 37.210 6.935 ;
        RECT 0.960 6.275 3.025 6.505 ;
        RECT 3.255 6.275 4.650 6.505 ;
        RECT 0.130 5.555 1.860 5.785 ;
        RECT 2.160 5.555 3.820 5.785 ;
        RECT 0.130 3.545 0.730 5.555 ;
        RECT 2.160 4.520 2.390 5.555 ;
        RECT 2.795 4.265 3.025 5.310 ;
        RECT 4.050 4.265 4.650 6.275 ;
        RECT 6.690 5.840 37.210 6.210 ;
        RECT 27.680 5.830 29.300 5.840 ;
        RECT 5.840 5.575 6.460 5.760 ;
        RECT 37.440 5.575 38.060 5.760 ;
        RECT 5.840 5.345 38.060 5.575 ;
        RECT 5.840 5.160 6.460 5.345 ;
        RECT 37.440 5.160 38.060 5.345 ;
        RECT 6.690 4.710 37.210 5.090 ;
        RECT 0.960 4.035 3.025 4.265 ;
        RECT 3.255 4.035 4.650 4.265 ;
        RECT 0.130 3.315 1.860 3.545 ;
        RECT 2.160 3.315 3.820 3.545 ;
        RECT 0.130 1.140 0.730 3.315 ;
        RECT 2.160 2.280 2.390 3.315 ;
        RECT 2.795 2.025 3.025 3.070 ;
        RECT 4.050 2.025 4.650 4.035 ;
        RECT 6.700 3.920 37.200 4.360 ;
        RECT 6.690 3.200 37.210 3.570 ;
        RECT 31.520 3.190 33.140 3.200 ;
        RECT 5.840 2.935 6.460 3.120 ;
        RECT 37.440 2.935 38.060 3.120 ;
        RECT 5.840 2.705 38.060 2.935 ;
        RECT 5.840 2.520 6.460 2.705 ;
        RECT 37.440 2.520 38.060 2.705 ;
        RECT 6.690 2.070 37.210 2.450 ;
        RECT 0.960 1.795 3.025 2.025 ;
        RECT 3.255 1.795 4.650 2.025 ;
        RECT 4.050 1.140 4.650 1.795 ;
        RECT 6.690 1.360 37.210 1.730 ;
        RECT 35.360 1.350 36.980 1.360 ;
        RECT 0.130 0.800 2.430 1.140 ;
        RECT 3.160 0.800 4.650 1.140 ;
        RECT 0.130 0.000 0.730 0.800 ;
        RECT 4.050 0.000 4.650 0.800 ;
        RECT 5.840 1.095 6.460 1.280 ;
        RECT 37.440 1.095 38.060 1.280 ;
        RECT 5.840 0.865 38.060 1.095 ;
        RECT 38.990 0.930 39.360 18.860 ;
        RECT 40.010 17.565 40.380 23.185 ;
        RECT 41.030 20.690 41.400 39.200 ;
        RECT 42.050 35.565 42.420 39.200 ;
        RECT 42.045 35.185 42.425 35.565 ;
        RECT 42.050 32.565 42.420 35.185 ;
        RECT 42.045 32.185 42.425 32.565 ;
        RECT 42.050 29.565 42.420 32.185 ;
        RECT 42.045 29.185 42.425 29.565 ;
        RECT 42.050 26.565 42.420 29.185 ;
        RECT 42.045 26.185 42.425 26.565 ;
        RECT 42.050 23.565 42.420 26.185 ;
        RECT 42.045 23.185 42.425 23.565 ;
        RECT 41.030 20.310 41.410 20.690 ;
        RECT 41.030 19.240 41.400 20.310 ;
        RECT 41.030 18.860 41.410 19.240 ;
        RECT 40.005 17.185 40.385 17.565 ;
        RECT 40.010 14.565 40.380 17.185 ;
        RECT 40.005 14.185 40.385 14.565 ;
        RECT 40.010 11.565 40.380 14.185 ;
        RECT 40.005 11.185 40.385 11.565 ;
        RECT 40.010 8.565 40.380 11.185 ;
        RECT 40.005 8.185 40.385 8.565 ;
        RECT 40.010 5.565 40.380 8.185 ;
        RECT 40.005 5.185 40.385 5.565 ;
        RECT 40.010 2.565 40.380 5.185 ;
        RECT 40.005 2.185 40.385 2.565 ;
        RECT 40.010 0.930 40.380 2.185 ;
        RECT 41.030 0.930 41.400 18.860 ;
        RECT 42.050 17.565 42.420 23.185 ;
        RECT 42.045 17.185 42.425 17.565 ;
        RECT 42.050 14.565 42.420 17.185 ;
        RECT 42.045 14.185 42.425 14.565 ;
        RECT 42.050 11.565 42.420 14.185 ;
        RECT 42.045 11.185 42.425 11.565 ;
        RECT 42.050 8.565 42.420 11.185 ;
        RECT 42.045 8.185 42.425 8.565 ;
        RECT 42.050 5.565 42.420 8.185 ;
        RECT 42.045 5.185 42.425 5.565 ;
        RECT 42.050 2.565 42.420 5.185 ;
        RECT 42.045 2.185 42.425 2.565 ;
        RECT 42.050 0.930 42.420 2.185 ;
        RECT 43.070 0.930 43.450 39.200 ;
        RECT 43.800 0.940 44.240 39.190 ;
        RECT 5.840 0.680 6.460 0.865 ;
        RECT 37.440 0.680 38.060 0.865 ;
        RECT 6.690 0.230 37.210 0.610 ;
      LAYER Metal2 ;
        RECT 6.700 38.895 9.560 39.275 ;
        RECT 37.560 38.335 37.940 38.715 ;
        RECT 0.240 36.685 0.620 37.065 ;
        RECT 4.160 36.685 4.540 37.065 ;
        RECT 6.700 37.055 9.560 37.435 ;
        RECT 6.700 35.170 9.560 35.550 ;
        RECT 6.700 34.410 9.560 34.790 ;
        RECT 0.240 33.685 0.620 34.065 ;
        RECT 4.160 33.685 4.540 34.065 ;
        RECT 6.700 32.570 9.560 32.950 ;
        RECT 0.240 30.685 0.620 31.065 ;
        RECT 4.160 30.685 4.540 31.065 ;
        RECT 6.700 30.730 9.560 31.110 ;
        RECT 6.700 28.845 9.560 29.225 ;
        RECT 6.700 28.085 9.560 28.465 ;
        RECT 0.240 27.685 0.620 28.065 ;
        RECT 4.160 27.685 4.540 28.065 ;
        RECT 6.700 26.245 9.560 26.625 ;
        RECT 0.240 24.685 0.620 25.065 ;
        RECT 4.160 24.685 4.540 25.065 ;
        RECT 6.700 24.405 9.560 24.785 ;
        RECT 0.240 21.685 0.620 22.065 ;
        RECT 4.160 21.685 4.540 22.065 ;
        RECT 10.335 21.695 12.085 25.505 ;
        RECT 14.175 21.695 15.925 27.345 ;
        RECT 18.015 21.695 19.765 29.990 ;
        RECT 21.855 21.695 23.605 31.830 ;
        RECT 25.695 21.695 27.445 33.670 ;
        RECT 29.535 21.695 31.285 36.315 ;
        RECT 33.375 21.695 35.125 38.155 ;
        RECT 37.560 36.495 37.940 36.875 ;
        RECT 40.005 35.185 40.385 35.565 ;
        RECT 42.045 35.185 42.425 35.565 ;
        RECT 43.830 35.185 44.210 35.565 ;
        RECT 37.560 33.850 37.940 34.230 ;
        RECT 37.560 32.010 37.940 32.390 ;
        RECT 40.005 32.185 40.385 32.565 ;
        RECT 42.045 32.185 42.425 32.565 ;
        RECT 43.830 32.185 44.210 32.565 ;
        RECT 37.560 30.170 37.940 30.550 ;
        RECT 40.005 29.185 40.385 29.565 ;
        RECT 42.045 29.185 42.425 29.565 ;
        RECT 43.830 29.185 44.210 29.565 ;
        RECT 37.560 27.525 37.940 27.905 ;
        RECT 40.005 26.185 40.385 26.565 ;
        RECT 42.045 26.185 42.425 26.565 ;
        RECT 43.830 26.185 44.210 26.565 ;
        RECT 37.560 25.685 37.940 26.065 ;
        RECT 37.560 23.845 37.940 24.225 ;
        RECT 40.005 23.185 40.385 23.565 ;
        RECT 42.045 23.185 42.425 23.565 ;
        RECT 43.830 23.185 44.210 23.565 ;
        RECT 9.100 21.310 9.480 21.500 ;
        RECT 12.940 21.310 13.320 21.500 ;
        RECT 16.780 21.310 17.160 21.500 ;
        RECT 20.620 21.310 21.000 21.500 ;
        RECT 24.460 21.310 24.840 21.500 ;
        RECT 28.300 21.310 28.680 21.500 ;
        RECT 32.140 21.310 32.520 21.500 ;
        RECT 35.980 21.310 36.360 21.500 ;
        RECT 3.430 20.500 44.480 21.310 ;
        RECT 0.240 18.685 0.620 19.065 ;
        RECT 3.430 19.050 4.240 20.500 ;
        RECT 38.990 20.310 39.370 20.500 ;
        RECT 41.030 20.310 41.410 20.500 ;
        RECT 43.070 20.310 43.450 20.500 ;
        RECT 38.990 19.050 39.370 19.240 ;
        RECT 41.030 19.050 41.410 19.240 ;
        RECT 43.070 19.050 43.450 19.240 ;
        RECT 3.430 18.240 44.480 19.050 ;
        RECT 7.180 18.050 7.560 18.240 ;
        RECT 11.020 18.050 11.400 18.240 ;
        RECT 14.860 18.050 15.240 18.240 ;
        RECT 18.700 18.050 19.080 18.240 ;
        RECT 22.540 18.050 22.920 18.240 ;
        RECT 26.380 18.050 26.760 18.240 ;
        RECT 30.220 18.050 30.600 18.240 ;
        RECT 34.060 18.050 34.440 18.240 ;
        RECT 0.240 15.685 0.620 16.065 ;
        RECT 2.520 13.395 2.870 17.585 ;
        RECT 0.240 12.685 0.620 13.065 ;
        RECT 3.150 12.040 3.500 15.955 ;
        RECT 4.160 15.685 4.540 16.065 ;
        RECT 6.700 14.720 9.560 15.100 ;
        RECT 12.255 14.000 14.005 17.855 ;
        RECT 4.160 12.685 4.540 13.065 ;
        RECT 6.700 12.880 9.560 13.260 ;
        RECT 16.095 12.155 17.845 17.855 ;
        RECT 2.745 11.715 3.500 12.040 ;
        RECT 2.300 11.030 2.680 11.410 ;
        RECT 6.700 11.035 9.560 11.415 ;
        RECT 6.700 10.275 9.560 10.655 ;
        RECT 0.240 9.685 0.620 10.065 ;
        RECT 4.160 9.685 4.540 10.065 ;
        RECT 19.935 9.515 21.685 17.855 ;
        RECT 6.700 8.395 9.560 8.775 ;
        RECT 23.775 7.675 25.525 17.855 ;
        RECT 0.240 6.685 0.620 7.065 ;
        RECT 4.160 6.685 4.540 7.065 ;
        RECT 6.700 6.555 9.560 6.935 ;
        RECT 27.615 5.830 29.365 17.855 ;
        RECT 6.700 4.710 9.560 5.090 ;
        RECT 0.240 3.685 0.620 4.065 ;
        RECT 4.160 3.685 4.540 4.065 ;
        RECT 6.700 3.950 9.560 4.330 ;
        RECT 31.455 3.190 33.205 17.855 ;
        RECT 6.700 2.070 9.560 2.450 ;
        RECT 35.295 1.350 37.045 17.855 ;
        RECT 40.005 17.185 40.385 17.565 ;
        RECT 42.045 17.185 42.425 17.565 ;
        RECT 43.830 17.185 44.210 17.565 ;
        RECT 37.560 15.280 37.940 15.660 ;
        RECT 40.005 14.185 40.385 14.565 ;
        RECT 42.045 14.185 42.425 14.565 ;
        RECT 43.830 14.185 44.210 14.565 ;
        RECT 37.560 13.440 37.940 13.820 ;
        RECT 37.560 11.595 37.940 11.975 ;
        RECT 40.005 11.185 40.385 11.565 ;
        RECT 42.045 11.185 42.425 11.565 ;
        RECT 43.830 11.185 44.210 11.565 ;
        RECT 37.560 8.955 37.940 9.335 ;
        RECT 40.005 8.185 40.385 8.565 ;
        RECT 42.045 8.185 42.425 8.565 ;
        RECT 43.830 8.185 44.210 8.565 ;
        RECT 37.560 7.115 37.940 7.495 ;
        RECT 37.560 5.270 37.940 5.650 ;
        RECT 40.005 5.185 40.385 5.565 ;
        RECT 42.045 5.185 42.425 5.565 ;
        RECT 43.830 5.185 44.210 5.565 ;
        RECT 37.560 2.630 37.940 3.010 ;
        RECT 40.005 2.185 40.385 2.565 ;
        RECT 42.045 2.185 42.425 2.565 ;
        RECT 43.830 2.185 44.210 2.565 ;
        RECT 0.240 0.685 0.620 1.065 ;
        RECT 4.160 0.685 4.540 1.065 ;
        RECT 37.560 0.790 37.940 1.170 ;
        RECT 6.700 0.230 9.560 0.610 ;
      LAYER Metal3 ;
        RECT 6.700 38.895 9.560 39.275 ;
        RECT 28.740 38.665 29.120 38.715 ;
        RECT 37.560 38.665 37.940 38.715 ;
        RECT 28.740 38.385 37.940 38.665 ;
        RECT 28.740 38.335 29.120 38.385 ;
        RECT 37.560 38.335 37.940 38.385 ;
        RECT 0.240 36.685 0.620 37.065 ;
        RECT 4.160 36.685 4.540 37.065 ;
        RECT 6.700 37.055 9.560 37.435 ;
        RECT 30.020 36.825 30.400 36.875 ;
        RECT 37.560 36.825 37.940 36.875 ;
        RECT 30.020 36.545 37.940 36.825 ;
        RECT 30.020 36.495 30.400 36.545 ;
        RECT 37.560 36.495 37.940 36.545 ;
        RECT 6.700 35.170 9.560 35.550 ;
        RECT 40.005 35.185 40.385 35.565 ;
        RECT 42.045 35.185 42.425 35.565 ;
        RECT 43.830 35.185 44.210 35.565 ;
        RECT 6.700 34.410 9.560 34.790 ;
        RECT 31.300 34.180 31.680 34.230 ;
        RECT 37.560 34.180 37.940 34.230 ;
        RECT 0.240 33.685 0.620 34.065 ;
        RECT 4.160 33.685 4.540 34.065 ;
        RECT 31.300 33.900 37.940 34.180 ;
        RECT 31.300 33.850 31.680 33.900 ;
        RECT 37.560 33.850 37.940 33.900 ;
        RECT 6.700 32.570 9.560 32.950 ;
        RECT 32.580 32.340 32.960 32.390 ;
        RECT 37.560 32.340 37.940 32.390 ;
        RECT 32.580 32.060 37.940 32.340 ;
        RECT 40.005 32.185 40.385 32.565 ;
        RECT 42.045 32.185 42.425 32.565 ;
        RECT 43.830 32.185 44.210 32.565 ;
        RECT 32.580 32.010 32.960 32.060 ;
        RECT 37.560 32.010 37.940 32.060 ;
        RECT 0.240 30.685 0.620 31.065 ;
        RECT 4.160 30.685 4.540 31.065 ;
        RECT 6.700 30.730 9.560 31.110 ;
        RECT 33.860 30.500 34.240 30.550 ;
        RECT 37.560 30.500 37.940 30.550 ;
        RECT 33.860 30.220 37.940 30.500 ;
        RECT 33.860 30.170 34.240 30.220 ;
        RECT 37.560 30.170 37.940 30.220 ;
        RECT 6.700 28.845 9.560 29.225 ;
        RECT 40.005 29.185 40.385 29.565 ;
        RECT 42.045 29.185 42.425 29.565 ;
        RECT 43.830 29.185 44.210 29.565 ;
        RECT 6.700 28.085 9.560 28.465 ;
        RECT 0.240 27.685 0.620 28.065 ;
        RECT 4.160 27.685 4.540 28.065 ;
        RECT 35.140 27.855 35.520 27.905 ;
        RECT 37.560 27.855 37.940 27.905 ;
        RECT 35.140 27.575 37.940 27.855 ;
        RECT 35.140 27.525 35.520 27.575 ;
        RECT 37.560 27.525 37.940 27.575 ;
        RECT 6.700 26.245 9.560 26.625 ;
        RECT 40.005 26.185 40.385 26.565 ;
        RECT 42.045 26.185 42.425 26.565 ;
        RECT 43.830 26.185 44.210 26.565 ;
        RECT 36.420 26.015 36.800 26.065 ;
        RECT 37.560 26.015 37.940 26.065 ;
        RECT 36.420 25.735 37.940 26.015 ;
        RECT 36.420 25.685 36.800 25.735 ;
        RECT 37.560 25.685 37.940 25.735 ;
        RECT 0.240 24.685 0.620 25.065 ;
        RECT 4.160 24.685 4.540 25.065 ;
        RECT 6.700 24.405 9.560 24.785 ;
        RECT 37.560 23.845 38.080 24.225 ;
        RECT 40.005 23.185 40.385 23.565 ;
        RECT 42.045 23.185 42.425 23.565 ;
        RECT 43.830 23.185 44.210 23.565 ;
        RECT 0.240 21.685 0.620 22.065 ;
        RECT 4.160 21.685 4.540 22.065 ;
        RECT 0.240 18.685 0.620 19.065 ;
        RECT 40.005 17.185 40.385 17.565 ;
        RECT 42.045 17.185 42.425 17.565 ;
        RECT 43.830 17.185 44.210 17.565 ;
        RECT 0.240 15.685 0.620 16.065 ;
        RECT 4.160 15.685 4.540 16.065 ;
        RECT 37.060 15.280 37.940 15.660 ;
        RECT 6.700 14.720 9.560 15.100 ;
        RECT 40.005 14.185 40.385 14.565 ;
        RECT 42.045 14.185 42.425 14.565 ;
        RECT 43.830 14.185 44.210 14.565 ;
        RECT 35.780 13.770 36.160 13.820 ;
        RECT 37.560 13.770 37.940 13.820 ;
        RECT 35.780 13.490 37.940 13.770 ;
        RECT 35.780 13.440 36.160 13.490 ;
        RECT 37.560 13.440 37.940 13.490 ;
        RECT 0.240 12.685 0.620 13.065 ;
        RECT 4.160 12.685 4.540 13.065 ;
        RECT 6.700 12.880 9.560 13.260 ;
        RECT 34.500 11.925 34.880 11.975 ;
        RECT 37.560 11.925 37.940 11.975 ;
        RECT 34.500 11.645 37.940 11.925 ;
        RECT 34.500 11.595 34.880 11.645 ;
        RECT 37.560 11.595 37.940 11.645 ;
        RECT 6.700 11.035 9.560 11.415 ;
        RECT 40.005 11.185 40.385 11.565 ;
        RECT 42.045 11.185 42.425 11.565 ;
        RECT 43.830 11.185 44.210 11.565 ;
        RECT 6.700 10.275 9.560 10.655 ;
        RECT 0.240 9.685 0.620 10.065 ;
        RECT 4.160 9.685 4.540 10.065 ;
        RECT 33.220 9.285 33.600 9.335 ;
        RECT 37.560 9.285 37.940 9.335 ;
        RECT 33.220 9.005 37.940 9.285 ;
        RECT 33.220 8.955 33.600 9.005 ;
        RECT 37.560 8.955 37.940 9.005 ;
        RECT 6.700 8.395 9.560 8.775 ;
        RECT 40.005 8.185 40.385 8.565 ;
        RECT 42.045 8.185 42.425 8.565 ;
        RECT 43.830 8.185 44.210 8.565 ;
        RECT 31.940 7.445 32.320 7.495 ;
        RECT 37.560 7.445 37.940 7.495 ;
        RECT 31.940 7.165 37.940 7.445 ;
        RECT 31.940 7.115 32.320 7.165 ;
        RECT 37.560 7.115 37.940 7.165 ;
        RECT 0.240 6.685 0.620 7.065 ;
        RECT 4.160 6.685 4.540 7.065 ;
        RECT 6.700 6.555 9.560 6.935 ;
        RECT 30.660 5.600 31.040 5.650 ;
        RECT 37.560 5.600 37.940 5.650 ;
        RECT 30.660 5.320 37.940 5.600 ;
        RECT 30.660 5.270 31.040 5.320 ;
        RECT 37.560 5.270 37.940 5.320 ;
        RECT 40.005 5.185 40.385 5.565 ;
        RECT 42.045 5.185 42.425 5.565 ;
        RECT 43.830 5.185 44.210 5.565 ;
        RECT 6.700 4.710 9.560 5.090 ;
        RECT 0.240 3.685 0.620 4.065 ;
        RECT 4.160 3.685 4.540 4.065 ;
        RECT 6.700 3.950 9.560 4.330 ;
        RECT 29.380 2.960 29.760 3.010 ;
        RECT 37.560 2.960 37.940 3.010 ;
        RECT 29.380 2.680 37.940 2.960 ;
        RECT 29.380 2.630 29.760 2.680 ;
        RECT 37.560 2.630 37.940 2.680 ;
        RECT 6.700 2.070 9.560 2.450 ;
        RECT 40.005 2.185 40.385 2.565 ;
        RECT 42.045 2.185 42.425 2.565 ;
        RECT 43.830 2.185 44.210 2.565 ;
        RECT 28.100 1.120 28.480 1.170 ;
        RECT 37.560 1.120 37.940 1.170 ;
        RECT 0.240 0.685 0.620 1.065 ;
        RECT 4.160 0.685 4.540 1.065 ;
        RECT 28.100 0.840 37.940 1.120 ;
        RECT 28.100 0.790 28.480 0.840 ;
        RECT 37.560 0.790 37.940 0.840 ;
        RECT 6.700 0.230 9.560 0.610 ;
  END
END efuse_array_16x1
END LIBRARY

