* eFuse array netlist with word_width=8, nwords=64
    
.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
X0 ZN I VSS VPW nfet_06v0 W=8.2e-07 L=6e-07  
X1 ZN I VDD VNW pfet_06v0 W=1.22e-06 L=5e-07
.ENDS

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
X00 ZN I VSS VPW nfet_06v0 W=8.2e-07 L=6e-07
X01 VSS I ZN VPW nfet_06v0 W=8.2e-07 L=6e-07
X10 ZN I VDD VNW pfet_06v0 W=1.22e-06 L=5e-07
X11 VDD I ZN VNW pfet_06v0 W=1.22e-06 L=5e-07
.ENDS

.subckt efuse_bitcell VSS SELECT ANODE
X0 ANODE CATHODE efuse
X1 CATHODE SELECT VSS VSS nfet_06v0 L=0.60u W=30.5u
.ends

.subckt efuse_senseamp  VDD PRESET_N OUT SENSE VSS FUSE
X2 net1 PRESET_N VDD VDD pfet_06v0 L=0.5u W=2.44u nf=2
x1 net2 OUT VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x2 net1 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
x3 net2 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X1 net1 SENSE FUSE VSS nfet_06v0 L=0.60u W=0.82u
.ends


.subckt efuse_bitline VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63] COL_PROG_N OUT
X0 VSS BIT_SEL[0] bitline efuse_bitcell
X1 VSS BIT_SEL[1] bitline efuse_bitcell
X2 VSS BIT_SEL[2] bitline efuse_bitcell
X3 VSS BIT_SEL[3] bitline efuse_bitcell
X4 VSS BIT_SEL[4] bitline efuse_bitcell
X5 VSS BIT_SEL[5] bitline efuse_bitcell
X6 VSS BIT_SEL[6] bitline efuse_bitcell
X7 VSS BIT_SEL[7] bitline efuse_bitcell
X8 VSS BIT_SEL[8] bitline efuse_bitcell
X9 VSS BIT_SEL[9] bitline efuse_bitcell
X10 VSS BIT_SEL[10] bitline efuse_bitcell
X11 VSS BIT_SEL[11] bitline efuse_bitcell
X12 VSS BIT_SEL[12] bitline efuse_bitcell
X13 VSS BIT_SEL[13] bitline efuse_bitcell
X14 VSS BIT_SEL[14] bitline efuse_bitcell
X15 VSS BIT_SEL[15] bitline efuse_bitcell
X16 VSS BIT_SEL[16] bitline efuse_bitcell
X17 VSS BIT_SEL[17] bitline efuse_bitcell
X18 VSS BIT_SEL[18] bitline efuse_bitcell
X19 VSS BIT_SEL[19] bitline efuse_bitcell
X20 VSS BIT_SEL[20] bitline efuse_bitcell
X21 VSS BIT_SEL[21] bitline efuse_bitcell
X22 VSS BIT_SEL[22] bitline efuse_bitcell
X23 VSS BIT_SEL[23] bitline efuse_bitcell
X24 VSS BIT_SEL[24] bitline efuse_bitcell
X25 VSS BIT_SEL[25] bitline efuse_bitcell
X26 VSS BIT_SEL[26] bitline efuse_bitcell
X27 VSS BIT_SEL[27] bitline efuse_bitcell
X28 VSS BIT_SEL[28] bitline efuse_bitcell
X29 VSS BIT_SEL[29] bitline efuse_bitcell
X30 VSS BIT_SEL[30] bitline efuse_bitcell
X31 VSS BIT_SEL[31] bitline efuse_bitcell
X32 VSS BIT_SEL[32] bitline efuse_bitcell
X33 VSS BIT_SEL[33] bitline efuse_bitcell
X34 VSS BIT_SEL[34] bitline efuse_bitcell
X35 VSS BIT_SEL[35] bitline efuse_bitcell
X36 VSS BIT_SEL[36] bitline efuse_bitcell
X37 VSS BIT_SEL[37] bitline efuse_bitcell
X38 VSS BIT_SEL[38] bitline efuse_bitcell
X39 VSS BIT_SEL[39] bitline efuse_bitcell
X40 VSS BIT_SEL[40] bitline efuse_bitcell
X41 VSS BIT_SEL[41] bitline efuse_bitcell
X42 VSS BIT_SEL[42] bitline efuse_bitcell
X43 VSS BIT_SEL[43] bitline efuse_bitcell
X44 VSS BIT_SEL[44] bitline efuse_bitcell
X45 VSS BIT_SEL[45] bitline efuse_bitcell
X46 VSS BIT_SEL[46] bitline efuse_bitcell
X47 VSS BIT_SEL[47] bitline efuse_bitcell
X48 VSS BIT_SEL[48] bitline efuse_bitcell
X49 VSS BIT_SEL[49] bitline efuse_bitcell
X50 VSS BIT_SEL[50] bitline efuse_bitcell
X51 VSS BIT_SEL[51] bitline efuse_bitcell
X52 VSS BIT_SEL[52] bitline efuse_bitcell
X53 VSS BIT_SEL[53] bitline efuse_bitcell
X54 VSS BIT_SEL[54] bitline efuse_bitcell
X55 VSS BIT_SEL[55] bitline efuse_bitcell
X56 VSS BIT_SEL[56] bitline efuse_bitcell
X57 VSS BIT_SEL[57] bitline efuse_bitcell
X58 VSS BIT_SEL[58] bitline efuse_bitcell
X59 VSS BIT_SEL[59] bitline efuse_bitcell
X60 VSS BIT_SEL[60] bitline efuse_bitcell
X61 VSS BIT_SEL[61] bitline efuse_bitcell
X62 VSS BIT_SEL[62] bitline efuse_bitcell
X63 VSS BIT_SEL[63] bitline efuse_bitcell
X0 bitline COL_PROG_N VDD VDD pfet_06v0 L=0.50u W=76.5u nf=2
X1 bitline COL_PROG_N VDD VDD pfet_06v0 L=0.50u W=76.5u nf=2
Xsense VDD PRESET_N OUT SENSE VSS bitline efuse_senseamp
.ends
    

.subckt efuse_array_64x8 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63] COL_PROG_N[0] OUT[0] COL_PROG_N[1] OUT[1] COL_PROG_N[2] OUT[2] COL_PROG_N[3] OUT[3] COL_PROG_N[4] OUT[4] COL_PROG_N[5] OUT[5] COL_PROG_N[6] OUT[6] COL_PROG_N[7] OUT[7] 
X0_0 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[0] OUT[0]  efuse_bitline
X0_1 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[1] OUT[1]  efuse_bitline
X0_2 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[2] OUT[2]  efuse_bitline
X0_3 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[3] OUT[3]  efuse_bitline
X0_4 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[4] OUT[4]  efuse_bitline
X0_5 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[5] OUT[5]  efuse_bitline
X0_6 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[6] OUT[6]  efuse_bitline
X0_7 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[7] OUT[7]  efuse_bitline

.ends
    
.end
    