VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_array_32x8
  CLASS BLOCK ;
  FOREIGN efuse_array_32x8 ;
  ORIGIN -24.960 -66.885 ;
  SIZE 76.930 BY 315.825 ;
  PIN COL_PROG_N[0]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 96.850 106.315 100.410 106.615 ;
    END
  END COL_PROG_N[0]
  PIN OUT[0]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 77.995 28.780 78.325 ;
    END
  END OUT[0]
  PIN COL_PROG_N[1]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 96.850 145.700 100.410 146.000 ;
    END
  END COL_PROG_N[1]
  PIN OUT[1]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 117.380 28.780 117.710 ;
    END
  END OUT[1]
  PIN COL_PROG_N[2]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 96.850 185.085 100.410 185.385 ;
    END
  END COL_PROG_N[2]
  PIN OUT[2]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 156.765 28.780 157.095 ;
    END
  END OUT[2]
  PIN COL_PROG_N[3]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 96.850 224.470 100.410 224.770 ;
    END
  END COL_PROG_N[3]
  PIN OUT[3]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 196.150 28.780 196.480 ;
    END
  END OUT[3]
  PIN COL_PROG_N[4]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 96.850 263.855 100.410 264.155 ;
    END
  END COL_PROG_N[4]
  PIN OUT[4]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 235.535 28.780 235.865 ;
    END
  END OUT[4]
  PIN COL_PROG_N[5]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 96.850 303.240 100.410 303.540 ;
    END
  END COL_PROG_N[5]
  PIN OUT[5]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 274.920 28.780 275.250 ;
    END
  END OUT[5]
  PIN COL_PROG_N[6]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 96.850 342.625 100.410 342.925 ;
    END
  END COL_PROG_N[6]
  PIN OUT[6]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 314.305 28.780 314.635 ;
    END
  END OUT[6]
  PIN COL_PROG_N[7]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 96.850 382.010 100.410 382.310 ;
    END
  END COL_PROG_N[7]
  PIN OUT[7]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 353.690 28.780 354.020 ;
    END
  END OUT[7]
  PIN PRESET_N
    ANTENNAGATEAREA 9.760000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.970 362.420 26.250 382.710 ;
        RECT 25.970 362.040 26.330 362.420 ;
        RECT 25.970 323.035 26.250 362.040 ;
        RECT 25.970 322.655 26.330 323.035 ;
        RECT 25.970 283.650 26.250 322.655 ;
        RECT 25.970 283.270 26.330 283.650 ;
        RECT 25.970 244.265 26.250 283.270 ;
        RECT 25.970 243.885 26.330 244.265 ;
        RECT 25.970 204.880 26.250 243.885 ;
        RECT 25.970 204.500 26.330 204.880 ;
        RECT 25.970 165.495 26.250 204.500 ;
        RECT 25.970 165.115 26.330 165.495 ;
        RECT 25.970 126.110 26.250 165.115 ;
        RECT 25.970 125.730 26.330 126.110 ;
        RECT 25.970 86.725 26.250 125.730 ;
        RECT 25.970 86.345 26.330 86.725 ;
        RECT 25.970 66.885 26.250 86.345 ;
    END
  END PRESET_N
  PIN SENSE
    ANTENNAGATEAREA 3.936000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.615 361.235 26.895 382.710 ;
        RECT 26.615 360.855 28.040 361.235 ;
        RECT 26.615 321.850 26.895 360.855 ;
        RECT 26.615 321.470 28.040 321.850 ;
        RECT 26.615 282.465 26.895 321.470 ;
        RECT 26.615 282.085 28.040 282.465 ;
        RECT 26.615 243.080 26.895 282.085 ;
        RECT 26.615 242.700 28.040 243.080 ;
        RECT 26.615 203.695 26.895 242.700 ;
        RECT 26.615 203.315 28.040 203.695 ;
        RECT 26.615 164.310 26.895 203.315 ;
        RECT 26.615 163.930 28.040 164.310 ;
        RECT 26.615 124.925 26.895 163.930 ;
        RECT 26.615 124.545 28.040 124.925 ;
        RECT 26.615 85.540 26.895 124.545 ;
        RECT 26.615 85.160 28.040 85.540 ;
        RECT 26.615 66.885 26.895 85.160 ;
    END
  END SENSE
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 63.880 66.885 66.880 382.710 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 28.670 66.885 29.670 382.710 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 31.430 66.885 34.430 382.710 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 97.400 66.885 101.650 382.710 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 25.030 66.885 26.030 382.710 ;
    END
  END VDD
  PIN BIT_SEL[0]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 62.700 366.805 62.980 382.085 ;
        RECT 62.660 366.425 63.040 366.805 ;
        RECT 62.700 327.420 62.980 366.425 ;
        RECT 62.660 327.040 63.040 327.420 ;
        RECT 62.700 288.035 62.980 327.040 ;
        RECT 62.660 287.655 63.040 288.035 ;
        RECT 62.700 248.650 62.980 287.655 ;
        RECT 62.660 248.270 63.040 248.650 ;
        RECT 62.700 209.265 62.980 248.270 ;
        RECT 62.660 208.885 63.040 209.265 ;
        RECT 62.700 169.880 62.980 208.885 ;
        RECT 62.660 169.500 63.040 169.880 ;
        RECT 62.700 130.495 62.980 169.500 ;
        RECT 62.660 130.115 63.040 130.495 ;
        RECT 62.700 91.110 62.980 130.115 ;
        RECT 62.660 90.730 63.040 91.110 ;
        RECT 62.700 66.885 62.980 90.730 ;
    END
  END BIT_SEL[0]
  PIN BIT_SEL[16]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 95.150 366.805 95.430 382.085 ;
        RECT 95.110 366.425 95.490 366.805 ;
        RECT 95.150 327.420 95.430 366.425 ;
        RECT 95.110 327.040 95.490 327.420 ;
        RECT 95.150 288.035 95.430 327.040 ;
        RECT 95.110 287.655 95.490 288.035 ;
        RECT 95.150 248.650 95.430 287.655 ;
        RECT 95.110 248.270 95.490 248.650 ;
        RECT 95.150 209.265 95.430 248.270 ;
        RECT 95.110 208.885 95.490 209.265 ;
        RECT 95.150 169.880 95.430 208.885 ;
        RECT 95.110 169.500 95.490 169.880 ;
        RECT 95.150 130.495 95.430 169.500 ;
        RECT 95.110 130.115 95.490 130.495 ;
        RECT 95.150 91.110 95.430 130.115 ;
        RECT 95.110 90.730 95.490 91.110 ;
        RECT 95.150 66.885 95.430 90.730 ;
    END
  END BIT_SEL[16]
  PIN BIT_SEL[17]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 94.510 358.240 94.790 382.085 ;
        RECT 94.470 357.860 94.850 358.240 ;
        RECT 94.510 318.855 94.790 357.860 ;
        RECT 94.470 318.475 94.850 318.855 ;
        RECT 94.510 279.470 94.790 318.475 ;
        RECT 94.470 279.090 94.850 279.470 ;
        RECT 94.510 240.085 94.790 279.090 ;
        RECT 94.470 239.705 94.850 240.085 ;
        RECT 94.510 200.700 94.790 239.705 ;
        RECT 94.470 200.320 94.850 200.700 ;
        RECT 94.510 161.315 94.790 200.320 ;
        RECT 94.470 160.935 94.850 161.315 ;
        RECT 94.510 121.930 94.790 160.935 ;
        RECT 94.470 121.550 94.850 121.930 ;
        RECT 94.510 82.545 94.790 121.550 ;
        RECT 94.470 82.165 94.850 82.545 ;
        RECT 94.510 66.885 94.790 82.165 ;
    END
  END BIT_SEL[17]
  PIN BIT_SEL[18]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 93.870 368.645 94.150 382.085 ;
        RECT 93.830 368.265 94.210 368.645 ;
        RECT 93.870 329.260 94.150 368.265 ;
        RECT 93.830 328.880 94.210 329.260 ;
        RECT 93.870 289.875 94.150 328.880 ;
        RECT 93.830 289.495 94.210 289.875 ;
        RECT 93.870 250.490 94.150 289.495 ;
        RECT 93.830 250.110 94.210 250.490 ;
        RECT 93.870 211.105 94.150 250.110 ;
        RECT 93.830 210.725 94.210 211.105 ;
        RECT 93.870 171.720 94.150 210.725 ;
        RECT 93.830 171.340 94.210 171.720 ;
        RECT 93.870 132.335 94.150 171.340 ;
        RECT 93.830 131.955 94.210 132.335 ;
        RECT 93.870 92.950 94.150 131.955 ;
        RECT 93.830 92.570 94.210 92.950 ;
        RECT 93.870 66.885 94.150 92.570 ;
    END
  END BIT_SEL[18]
  PIN BIT_SEL[19]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 93.230 356.400 93.510 382.085 ;
        RECT 93.190 356.020 93.570 356.400 ;
        RECT 93.230 317.015 93.510 356.020 ;
        RECT 93.190 316.635 93.570 317.015 ;
        RECT 93.230 277.630 93.510 316.635 ;
        RECT 93.190 277.250 93.570 277.630 ;
        RECT 93.230 238.245 93.510 277.250 ;
        RECT 93.190 237.865 93.570 238.245 ;
        RECT 93.230 198.860 93.510 237.865 ;
        RECT 93.190 198.480 93.570 198.860 ;
        RECT 93.230 159.475 93.510 198.480 ;
        RECT 93.190 159.095 93.570 159.475 ;
        RECT 93.230 120.090 93.510 159.095 ;
        RECT 93.190 119.710 93.570 120.090 ;
        RECT 93.230 80.705 93.510 119.710 ;
        RECT 93.190 80.325 93.570 80.705 ;
        RECT 93.230 66.885 93.510 80.325 ;
    END
  END BIT_SEL[19]
  PIN BIT_SEL[20]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 92.590 370.485 92.870 382.085 ;
        RECT 92.550 370.105 92.930 370.485 ;
        RECT 92.590 331.100 92.870 370.105 ;
        RECT 92.550 330.720 92.930 331.100 ;
        RECT 92.590 291.715 92.870 330.720 ;
        RECT 92.550 291.335 92.930 291.715 ;
        RECT 92.590 252.330 92.870 291.335 ;
        RECT 92.550 251.950 92.930 252.330 ;
        RECT 92.590 212.945 92.870 251.950 ;
        RECT 92.550 212.565 92.930 212.945 ;
        RECT 92.590 173.560 92.870 212.565 ;
        RECT 92.550 173.180 92.930 173.560 ;
        RECT 92.590 134.175 92.870 173.180 ;
        RECT 92.550 133.795 92.930 134.175 ;
        RECT 92.590 94.790 92.870 133.795 ;
        RECT 92.550 94.410 92.930 94.790 ;
        RECT 92.590 66.885 92.870 94.410 ;
    END
  END BIT_SEL[20]
  PIN BIT_SEL[21]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 91.950 354.555 92.230 382.085 ;
        RECT 91.910 354.175 92.290 354.555 ;
        RECT 91.950 315.170 92.230 354.175 ;
        RECT 91.910 314.790 92.290 315.170 ;
        RECT 91.950 275.785 92.230 314.790 ;
        RECT 91.910 275.405 92.290 275.785 ;
        RECT 91.950 236.400 92.230 275.405 ;
        RECT 91.910 236.020 92.290 236.400 ;
        RECT 91.950 197.015 92.230 236.020 ;
        RECT 91.910 196.635 92.290 197.015 ;
        RECT 91.950 157.630 92.230 196.635 ;
        RECT 91.910 157.250 92.290 157.630 ;
        RECT 91.950 118.245 92.230 157.250 ;
        RECT 91.910 117.865 92.290 118.245 ;
        RECT 91.950 78.860 92.230 117.865 ;
        RECT 91.910 78.480 92.290 78.860 ;
        RECT 91.950 66.885 92.230 78.480 ;
    END
  END BIT_SEL[21]
  PIN BIT_SEL[22]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 91.310 373.130 91.590 382.085 ;
        RECT 91.270 372.750 91.650 373.130 ;
        RECT 91.310 333.745 91.590 372.750 ;
        RECT 91.270 333.365 91.650 333.745 ;
        RECT 91.310 294.360 91.590 333.365 ;
        RECT 91.270 293.980 91.650 294.360 ;
        RECT 91.310 254.975 91.590 293.980 ;
        RECT 91.270 254.595 91.650 254.975 ;
        RECT 91.310 215.590 91.590 254.595 ;
        RECT 91.270 215.210 91.650 215.590 ;
        RECT 91.310 176.205 91.590 215.210 ;
        RECT 91.270 175.825 91.650 176.205 ;
        RECT 91.310 136.820 91.590 175.825 ;
        RECT 91.270 136.440 91.650 136.820 ;
        RECT 91.310 97.435 91.590 136.440 ;
        RECT 91.270 97.055 91.650 97.435 ;
        RECT 91.310 66.885 91.590 97.055 ;
    END
  END BIT_SEL[22]
  PIN BIT_SEL[23]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 90.670 351.915 90.950 382.085 ;
        RECT 90.630 351.535 91.010 351.915 ;
        RECT 90.670 312.530 90.950 351.535 ;
        RECT 90.630 312.150 91.010 312.530 ;
        RECT 90.670 273.145 90.950 312.150 ;
        RECT 90.630 272.765 91.010 273.145 ;
        RECT 90.670 233.760 90.950 272.765 ;
        RECT 90.630 233.380 91.010 233.760 ;
        RECT 90.670 194.375 90.950 233.380 ;
        RECT 90.630 193.995 91.010 194.375 ;
        RECT 90.670 154.990 90.950 193.995 ;
        RECT 90.630 154.610 91.010 154.990 ;
        RECT 90.670 115.605 90.950 154.610 ;
        RECT 90.630 115.225 91.010 115.605 ;
        RECT 90.670 76.220 90.950 115.225 ;
        RECT 90.630 75.840 91.010 76.220 ;
        RECT 90.670 66.885 90.950 75.840 ;
    END
  END BIT_SEL[23]
  PIN BIT_SEL[24]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 90.030 374.970 90.310 382.085 ;
        RECT 89.990 374.590 90.370 374.970 ;
        RECT 90.030 335.585 90.310 374.590 ;
        RECT 89.990 335.205 90.370 335.585 ;
        RECT 90.030 296.200 90.310 335.205 ;
        RECT 89.990 295.820 90.370 296.200 ;
        RECT 90.030 256.815 90.310 295.820 ;
        RECT 89.990 256.435 90.370 256.815 ;
        RECT 90.030 217.430 90.310 256.435 ;
        RECT 89.990 217.050 90.370 217.430 ;
        RECT 90.030 178.045 90.310 217.050 ;
        RECT 89.990 177.665 90.370 178.045 ;
        RECT 90.030 138.660 90.310 177.665 ;
        RECT 89.990 138.280 90.370 138.660 ;
        RECT 90.030 99.275 90.310 138.280 ;
        RECT 89.990 98.895 90.370 99.275 ;
        RECT 90.030 66.885 90.310 98.895 ;
    END
  END BIT_SEL[24]
  PIN BIT_SEL[25]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 89.390 350.075 89.670 382.085 ;
        RECT 89.350 349.695 89.730 350.075 ;
        RECT 89.390 310.690 89.670 349.695 ;
        RECT 89.350 310.310 89.730 310.690 ;
        RECT 89.390 271.305 89.670 310.310 ;
        RECT 89.350 270.925 89.730 271.305 ;
        RECT 89.390 231.920 89.670 270.925 ;
        RECT 89.350 231.540 89.730 231.920 ;
        RECT 89.390 192.535 89.670 231.540 ;
        RECT 89.350 192.155 89.730 192.535 ;
        RECT 89.390 153.150 89.670 192.155 ;
        RECT 89.350 152.770 89.730 153.150 ;
        RECT 89.390 113.765 89.670 152.770 ;
        RECT 89.350 113.385 89.730 113.765 ;
        RECT 89.390 74.380 89.670 113.385 ;
        RECT 89.350 74.000 89.730 74.380 ;
        RECT 89.390 66.885 89.670 74.000 ;
    END
  END BIT_SEL[25]
  PIN BIT_SEL[26]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 88.750 376.810 89.030 382.085 ;
        RECT 88.710 376.430 89.090 376.810 ;
        RECT 88.750 337.425 89.030 376.430 ;
        RECT 88.710 337.045 89.090 337.425 ;
        RECT 88.750 298.040 89.030 337.045 ;
        RECT 88.710 297.660 89.090 298.040 ;
        RECT 88.750 258.655 89.030 297.660 ;
        RECT 88.710 258.275 89.090 258.655 ;
        RECT 88.750 219.270 89.030 258.275 ;
        RECT 88.710 218.890 89.090 219.270 ;
        RECT 88.750 179.885 89.030 218.890 ;
        RECT 88.710 179.505 89.090 179.885 ;
        RECT 88.750 140.500 89.030 179.505 ;
        RECT 88.710 140.120 89.090 140.500 ;
        RECT 88.750 101.115 89.030 140.120 ;
        RECT 88.710 100.735 89.090 101.115 ;
        RECT 88.750 66.885 89.030 100.735 ;
    END
  END BIT_SEL[26]
  PIN BIT_SEL[27]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 88.110 348.230 88.390 382.085 ;
        RECT 88.070 347.850 88.450 348.230 ;
        RECT 88.110 308.845 88.390 347.850 ;
        RECT 88.070 308.465 88.450 308.845 ;
        RECT 88.110 269.460 88.390 308.465 ;
        RECT 88.070 269.080 88.450 269.460 ;
        RECT 88.110 230.075 88.390 269.080 ;
        RECT 88.070 229.695 88.450 230.075 ;
        RECT 88.110 190.690 88.390 229.695 ;
        RECT 88.070 190.310 88.450 190.690 ;
        RECT 88.110 151.305 88.390 190.310 ;
        RECT 88.070 150.925 88.450 151.305 ;
        RECT 88.110 111.920 88.390 150.925 ;
        RECT 88.070 111.540 88.450 111.920 ;
        RECT 88.110 72.535 88.390 111.540 ;
        RECT 88.070 72.155 88.450 72.535 ;
        RECT 88.110 66.885 88.390 72.155 ;
    END
  END BIT_SEL[27]
  PIN BIT_SEL[28]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 87.470 379.455 87.750 382.085 ;
        RECT 87.430 379.075 87.810 379.455 ;
        RECT 87.470 340.070 87.750 379.075 ;
        RECT 87.430 339.690 87.810 340.070 ;
        RECT 87.470 300.685 87.750 339.690 ;
        RECT 87.430 300.305 87.810 300.685 ;
        RECT 87.470 261.300 87.750 300.305 ;
        RECT 87.430 260.920 87.810 261.300 ;
        RECT 87.470 221.915 87.750 260.920 ;
        RECT 87.430 221.535 87.810 221.915 ;
        RECT 87.470 182.530 87.750 221.535 ;
        RECT 87.430 182.150 87.810 182.530 ;
        RECT 87.470 143.145 87.750 182.150 ;
        RECT 87.430 142.765 87.810 143.145 ;
        RECT 87.470 103.760 87.750 142.765 ;
        RECT 87.430 103.380 87.810 103.760 ;
        RECT 87.470 66.885 87.750 103.380 ;
    END
  END BIT_SEL[28]
  PIN BIT_SEL[29]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 86.830 345.590 87.110 382.085 ;
        RECT 86.790 345.210 87.170 345.590 ;
        RECT 86.830 306.205 87.110 345.210 ;
        RECT 86.790 305.825 87.170 306.205 ;
        RECT 86.830 266.820 87.110 305.825 ;
        RECT 86.790 266.440 87.170 266.820 ;
        RECT 86.830 227.435 87.110 266.440 ;
        RECT 86.790 227.055 87.170 227.435 ;
        RECT 86.830 188.050 87.110 227.055 ;
        RECT 86.790 187.670 87.170 188.050 ;
        RECT 86.830 148.665 87.110 187.670 ;
        RECT 86.790 148.285 87.170 148.665 ;
        RECT 86.830 109.280 87.110 148.285 ;
        RECT 86.790 108.900 87.170 109.280 ;
        RECT 86.830 69.895 87.110 108.900 ;
        RECT 86.790 69.515 87.170 69.895 ;
        RECT 86.830 66.885 87.110 69.515 ;
    END
  END BIT_SEL[29]
  PIN BIT_SEL[30]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 86.190 381.295 86.470 382.085 ;
        RECT 86.150 380.915 86.530 381.295 ;
        RECT 86.190 341.910 86.470 380.915 ;
        RECT 86.150 341.530 86.530 341.910 ;
        RECT 86.190 302.525 86.470 341.530 ;
        RECT 86.150 302.145 86.530 302.525 ;
        RECT 86.190 263.140 86.470 302.145 ;
        RECT 86.150 262.760 86.530 263.140 ;
        RECT 86.190 223.755 86.470 262.760 ;
        RECT 86.150 223.375 86.530 223.755 ;
        RECT 86.190 184.370 86.470 223.375 ;
        RECT 86.150 183.990 86.530 184.370 ;
        RECT 86.190 144.985 86.470 183.990 ;
        RECT 86.150 144.605 86.530 144.985 ;
        RECT 86.190 105.600 86.470 144.605 ;
        RECT 86.150 105.220 86.530 105.600 ;
        RECT 86.190 66.885 86.470 105.220 ;
    END
  END BIT_SEL[30]
  PIN BIT_SEL[31]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 85.550 343.750 85.830 382.085 ;
        RECT 85.510 343.370 85.890 343.750 ;
        RECT 85.550 304.365 85.830 343.370 ;
        RECT 85.510 303.985 85.890 304.365 ;
        RECT 85.550 264.980 85.830 303.985 ;
        RECT 85.510 264.600 85.890 264.980 ;
        RECT 85.550 225.595 85.830 264.600 ;
        RECT 85.510 225.215 85.890 225.595 ;
        RECT 85.550 186.210 85.830 225.215 ;
        RECT 85.510 185.830 85.890 186.210 ;
        RECT 85.550 146.825 85.830 185.830 ;
        RECT 85.510 146.445 85.890 146.825 ;
        RECT 85.550 107.440 85.830 146.445 ;
        RECT 85.510 107.060 85.890 107.440 ;
        RECT 85.550 68.055 85.830 107.060 ;
        RECT 85.510 67.675 85.890 68.055 ;
        RECT 85.550 66.885 85.830 67.675 ;
    END
  END BIT_SEL[31]
  PIN BIT_SEL[1]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 62.060 358.240 62.340 382.085 ;
        RECT 62.020 357.860 62.400 358.240 ;
        RECT 62.060 318.855 62.340 357.860 ;
        RECT 62.020 318.475 62.400 318.855 ;
        RECT 62.060 279.470 62.340 318.475 ;
        RECT 62.020 279.090 62.400 279.470 ;
        RECT 62.060 240.085 62.340 279.090 ;
        RECT 62.020 239.705 62.400 240.085 ;
        RECT 62.060 200.700 62.340 239.705 ;
        RECT 62.020 200.320 62.400 200.700 ;
        RECT 62.060 161.315 62.340 200.320 ;
        RECT 62.020 160.935 62.400 161.315 ;
        RECT 62.060 121.930 62.340 160.935 ;
        RECT 62.020 121.550 62.400 121.930 ;
        RECT 62.060 82.545 62.340 121.550 ;
        RECT 62.020 82.165 62.400 82.545 ;
        RECT 62.060 66.885 62.340 82.165 ;
    END
  END BIT_SEL[1]
  PIN BIT_SEL[2]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 61.420 368.645 61.700 382.085 ;
        RECT 61.380 368.265 61.760 368.645 ;
        RECT 61.420 329.260 61.700 368.265 ;
        RECT 61.380 328.880 61.760 329.260 ;
        RECT 61.420 289.875 61.700 328.880 ;
        RECT 61.380 289.495 61.760 289.875 ;
        RECT 61.420 250.490 61.700 289.495 ;
        RECT 61.380 250.110 61.760 250.490 ;
        RECT 61.420 211.105 61.700 250.110 ;
        RECT 61.380 210.725 61.760 211.105 ;
        RECT 61.420 171.720 61.700 210.725 ;
        RECT 61.380 171.340 61.760 171.720 ;
        RECT 61.420 132.335 61.700 171.340 ;
        RECT 61.380 131.955 61.760 132.335 ;
        RECT 61.420 92.950 61.700 131.955 ;
        RECT 61.380 92.570 61.760 92.950 ;
        RECT 61.420 66.885 61.700 92.570 ;
    END
  END BIT_SEL[2]
  PIN BIT_SEL[3]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 60.780 356.400 61.060 382.085 ;
        RECT 60.740 356.020 61.120 356.400 ;
        RECT 60.780 317.015 61.060 356.020 ;
        RECT 60.740 316.635 61.120 317.015 ;
        RECT 60.780 277.630 61.060 316.635 ;
        RECT 60.740 277.250 61.120 277.630 ;
        RECT 60.780 238.245 61.060 277.250 ;
        RECT 60.740 237.865 61.120 238.245 ;
        RECT 60.780 198.860 61.060 237.865 ;
        RECT 60.740 198.480 61.120 198.860 ;
        RECT 60.780 159.475 61.060 198.480 ;
        RECT 60.740 159.095 61.120 159.475 ;
        RECT 60.780 120.090 61.060 159.095 ;
        RECT 60.740 119.710 61.120 120.090 ;
        RECT 60.780 80.705 61.060 119.710 ;
        RECT 60.740 80.325 61.120 80.705 ;
        RECT 60.780 66.885 61.060 80.325 ;
    END
  END BIT_SEL[3]
  PIN BIT_SEL[4]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 60.140 370.485 60.420 382.085 ;
        RECT 60.100 370.105 60.480 370.485 ;
        RECT 60.140 331.100 60.420 370.105 ;
        RECT 60.100 330.720 60.480 331.100 ;
        RECT 60.140 291.715 60.420 330.720 ;
        RECT 60.100 291.335 60.480 291.715 ;
        RECT 60.140 252.330 60.420 291.335 ;
        RECT 60.100 251.950 60.480 252.330 ;
        RECT 60.140 212.945 60.420 251.950 ;
        RECT 60.100 212.565 60.480 212.945 ;
        RECT 60.140 173.560 60.420 212.565 ;
        RECT 60.100 173.180 60.480 173.560 ;
        RECT 60.140 134.175 60.420 173.180 ;
        RECT 60.100 133.795 60.480 134.175 ;
        RECT 60.140 94.790 60.420 133.795 ;
        RECT 60.100 94.410 60.480 94.790 ;
        RECT 60.140 66.885 60.420 94.410 ;
    END
  END BIT_SEL[4]
  PIN BIT_SEL[5]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 59.500 354.555 59.780 382.085 ;
        RECT 59.460 354.175 59.840 354.555 ;
        RECT 59.500 315.170 59.780 354.175 ;
        RECT 59.460 314.790 59.840 315.170 ;
        RECT 59.500 275.785 59.780 314.790 ;
        RECT 59.460 275.405 59.840 275.785 ;
        RECT 59.500 236.400 59.780 275.405 ;
        RECT 59.460 236.020 59.840 236.400 ;
        RECT 59.500 197.015 59.780 236.020 ;
        RECT 59.460 196.635 59.840 197.015 ;
        RECT 59.500 157.630 59.780 196.635 ;
        RECT 59.460 157.250 59.840 157.630 ;
        RECT 59.500 118.245 59.780 157.250 ;
        RECT 59.460 117.865 59.840 118.245 ;
        RECT 59.500 78.860 59.780 117.865 ;
        RECT 59.460 78.480 59.840 78.860 ;
        RECT 59.500 66.885 59.780 78.480 ;
    END
  END BIT_SEL[5]
  PIN BIT_SEL[6]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 58.860 373.130 59.140 382.085 ;
        RECT 58.820 372.750 59.200 373.130 ;
        RECT 58.860 333.745 59.140 372.750 ;
        RECT 58.820 333.365 59.200 333.745 ;
        RECT 58.860 294.360 59.140 333.365 ;
        RECT 58.820 293.980 59.200 294.360 ;
        RECT 58.860 254.975 59.140 293.980 ;
        RECT 58.820 254.595 59.200 254.975 ;
        RECT 58.860 215.590 59.140 254.595 ;
        RECT 58.820 215.210 59.200 215.590 ;
        RECT 58.860 176.205 59.140 215.210 ;
        RECT 58.820 175.825 59.200 176.205 ;
        RECT 58.860 136.820 59.140 175.825 ;
        RECT 58.820 136.440 59.200 136.820 ;
        RECT 58.860 97.435 59.140 136.440 ;
        RECT 58.820 97.055 59.200 97.435 ;
        RECT 58.860 66.885 59.140 97.055 ;
    END
  END BIT_SEL[6]
  PIN BIT_SEL[7]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 58.220 351.915 58.500 382.085 ;
        RECT 58.180 351.535 58.560 351.915 ;
        RECT 58.220 312.530 58.500 351.535 ;
        RECT 58.180 312.150 58.560 312.530 ;
        RECT 58.220 273.145 58.500 312.150 ;
        RECT 58.180 272.765 58.560 273.145 ;
        RECT 58.220 233.760 58.500 272.765 ;
        RECT 58.180 233.380 58.560 233.760 ;
        RECT 58.220 194.375 58.500 233.380 ;
        RECT 58.180 193.995 58.560 194.375 ;
        RECT 58.220 154.990 58.500 193.995 ;
        RECT 58.180 154.610 58.560 154.990 ;
        RECT 58.220 115.605 58.500 154.610 ;
        RECT 58.180 115.225 58.560 115.605 ;
        RECT 58.220 76.220 58.500 115.225 ;
        RECT 58.180 75.840 58.560 76.220 ;
        RECT 58.220 66.885 58.500 75.840 ;
    END
  END BIT_SEL[7]
  PIN BIT_SEL[8]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 57.580 374.970 57.860 382.085 ;
        RECT 57.540 374.590 57.920 374.970 ;
        RECT 57.580 335.585 57.860 374.590 ;
        RECT 57.540 335.205 57.920 335.585 ;
        RECT 57.580 296.200 57.860 335.205 ;
        RECT 57.540 295.820 57.920 296.200 ;
        RECT 57.580 256.815 57.860 295.820 ;
        RECT 57.540 256.435 57.920 256.815 ;
        RECT 57.580 217.430 57.860 256.435 ;
        RECT 57.540 217.050 57.920 217.430 ;
        RECT 57.580 178.045 57.860 217.050 ;
        RECT 57.540 177.665 57.920 178.045 ;
        RECT 57.580 138.660 57.860 177.665 ;
        RECT 57.540 138.280 57.920 138.660 ;
        RECT 57.580 99.275 57.860 138.280 ;
        RECT 57.540 98.895 57.920 99.275 ;
        RECT 57.580 66.885 57.860 98.895 ;
    END
  END BIT_SEL[8]
  PIN BIT_SEL[9]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 56.940 350.075 57.220 382.085 ;
        RECT 56.900 349.695 57.280 350.075 ;
        RECT 56.940 310.690 57.220 349.695 ;
        RECT 56.900 310.310 57.280 310.690 ;
        RECT 56.940 271.305 57.220 310.310 ;
        RECT 56.900 270.925 57.280 271.305 ;
        RECT 56.940 231.920 57.220 270.925 ;
        RECT 56.900 231.540 57.280 231.920 ;
        RECT 56.940 192.535 57.220 231.540 ;
        RECT 56.900 192.155 57.280 192.535 ;
        RECT 56.940 153.150 57.220 192.155 ;
        RECT 56.900 152.770 57.280 153.150 ;
        RECT 56.940 113.765 57.220 152.770 ;
        RECT 56.900 113.385 57.280 113.765 ;
        RECT 56.940 74.380 57.220 113.385 ;
        RECT 56.900 74.000 57.280 74.380 ;
        RECT 56.940 66.885 57.220 74.000 ;
    END
  END BIT_SEL[9]
  PIN BIT_SEL[10]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 56.300 376.810 56.580 382.085 ;
        RECT 56.260 376.430 56.640 376.810 ;
        RECT 56.300 337.425 56.580 376.430 ;
        RECT 56.260 337.045 56.640 337.425 ;
        RECT 56.300 298.040 56.580 337.045 ;
        RECT 56.260 297.660 56.640 298.040 ;
        RECT 56.300 258.655 56.580 297.660 ;
        RECT 56.260 258.275 56.640 258.655 ;
        RECT 56.300 219.270 56.580 258.275 ;
        RECT 56.260 218.890 56.640 219.270 ;
        RECT 56.300 179.885 56.580 218.890 ;
        RECT 56.260 179.505 56.640 179.885 ;
        RECT 56.300 140.500 56.580 179.505 ;
        RECT 56.260 140.120 56.640 140.500 ;
        RECT 56.300 101.115 56.580 140.120 ;
        RECT 56.260 100.735 56.640 101.115 ;
        RECT 56.300 66.885 56.580 100.735 ;
    END
  END BIT_SEL[10]
  PIN BIT_SEL[11]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 55.660 348.230 55.940 382.085 ;
        RECT 55.620 347.850 56.000 348.230 ;
        RECT 55.660 308.845 55.940 347.850 ;
        RECT 55.620 308.465 56.000 308.845 ;
        RECT 55.660 269.460 55.940 308.465 ;
        RECT 55.620 269.080 56.000 269.460 ;
        RECT 55.660 230.075 55.940 269.080 ;
        RECT 55.620 229.695 56.000 230.075 ;
        RECT 55.660 190.690 55.940 229.695 ;
        RECT 55.620 190.310 56.000 190.690 ;
        RECT 55.660 151.305 55.940 190.310 ;
        RECT 55.620 150.925 56.000 151.305 ;
        RECT 55.660 111.920 55.940 150.925 ;
        RECT 55.620 111.540 56.000 111.920 ;
        RECT 55.660 72.535 55.940 111.540 ;
        RECT 55.620 72.155 56.000 72.535 ;
        RECT 55.660 66.885 55.940 72.155 ;
    END
  END BIT_SEL[11]
  PIN BIT_SEL[12]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 55.020 379.455 55.300 382.085 ;
        RECT 54.980 379.075 55.360 379.455 ;
        RECT 55.020 340.070 55.300 379.075 ;
        RECT 54.980 339.690 55.360 340.070 ;
        RECT 55.020 300.685 55.300 339.690 ;
        RECT 54.980 300.305 55.360 300.685 ;
        RECT 55.020 261.300 55.300 300.305 ;
        RECT 54.980 260.920 55.360 261.300 ;
        RECT 55.020 221.915 55.300 260.920 ;
        RECT 54.980 221.535 55.360 221.915 ;
        RECT 55.020 182.530 55.300 221.535 ;
        RECT 54.980 182.150 55.360 182.530 ;
        RECT 55.020 143.145 55.300 182.150 ;
        RECT 54.980 142.765 55.360 143.145 ;
        RECT 55.020 103.760 55.300 142.765 ;
        RECT 54.980 103.380 55.360 103.760 ;
        RECT 55.020 66.885 55.300 103.380 ;
    END
  END BIT_SEL[12]
  PIN BIT_SEL[13]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 54.380 345.590 54.660 382.085 ;
        RECT 54.340 345.210 54.720 345.590 ;
        RECT 54.380 306.205 54.660 345.210 ;
        RECT 54.340 305.825 54.720 306.205 ;
        RECT 54.380 266.820 54.660 305.825 ;
        RECT 54.340 266.440 54.720 266.820 ;
        RECT 54.380 227.435 54.660 266.440 ;
        RECT 54.340 227.055 54.720 227.435 ;
        RECT 54.380 188.050 54.660 227.055 ;
        RECT 54.340 187.670 54.720 188.050 ;
        RECT 54.380 148.665 54.660 187.670 ;
        RECT 54.340 148.285 54.720 148.665 ;
        RECT 54.380 109.280 54.660 148.285 ;
        RECT 54.340 108.900 54.720 109.280 ;
        RECT 54.380 69.895 54.660 108.900 ;
        RECT 54.340 69.515 54.720 69.895 ;
        RECT 54.380 66.885 54.660 69.515 ;
    END
  END BIT_SEL[13]
  PIN BIT_SEL[14]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 53.740 381.295 54.020 382.085 ;
        RECT 53.700 380.915 54.080 381.295 ;
        RECT 53.740 341.910 54.020 380.915 ;
        RECT 53.700 341.530 54.080 341.910 ;
        RECT 53.740 302.525 54.020 341.530 ;
        RECT 53.700 302.145 54.080 302.525 ;
        RECT 53.740 263.140 54.020 302.145 ;
        RECT 53.700 262.760 54.080 263.140 ;
        RECT 53.740 223.755 54.020 262.760 ;
        RECT 53.700 223.375 54.080 223.755 ;
        RECT 53.740 184.370 54.020 223.375 ;
        RECT 53.700 183.990 54.080 184.370 ;
        RECT 53.740 144.985 54.020 183.990 ;
        RECT 53.700 144.605 54.080 144.985 ;
        RECT 53.740 105.600 54.020 144.605 ;
        RECT 53.700 105.220 54.080 105.600 ;
        RECT 53.740 66.885 54.020 105.220 ;
    END
  END BIT_SEL[14]
  PIN BIT_SEL[15]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 53.100 343.750 53.380 382.085 ;
        RECT 53.060 343.370 53.440 343.750 ;
        RECT 53.100 304.365 53.380 343.370 ;
        RECT 53.060 303.985 53.440 304.365 ;
        RECT 53.100 264.980 53.380 303.985 ;
        RECT 53.060 264.600 53.440 264.980 ;
        RECT 53.100 225.595 53.380 264.600 ;
        RECT 53.060 225.215 53.440 225.595 ;
        RECT 53.100 186.210 53.380 225.215 ;
        RECT 53.060 185.830 53.440 186.210 ;
        RECT 53.100 146.825 53.380 185.830 ;
        RECT 53.060 146.445 53.440 146.825 ;
        RECT 53.100 107.440 53.380 146.445 ;
        RECT 53.060 107.060 53.440 107.440 ;
        RECT 53.100 68.055 53.380 107.060 ;
        RECT 53.060 67.675 53.440 68.055 ;
        RECT 53.100 66.885 53.380 67.675 ;
    END
  END BIT_SEL[15]
  OBS
      LAYER Metal1 ;
        RECT 25.090 363.855 25.690 382.710 ;
        RECT 29.010 363.855 29.610 382.710 ;
        RECT 31.650 381.475 62.170 381.855 ;
        RECT 64.100 381.475 94.620 381.855 ;
        RECT 30.800 381.220 31.420 381.405 ;
        RECT 62.400 381.220 63.020 381.405 ;
        RECT 30.800 380.990 63.020 381.220 ;
        RECT 30.800 380.805 31.420 380.990 ;
        RECT 62.400 380.805 63.020 380.990 ;
        RECT 63.250 381.220 63.870 381.405 ;
        RECT 94.850 381.220 95.470 381.405 ;
        RECT 63.250 380.990 95.470 381.220 ;
        RECT 63.250 380.805 63.870 380.990 ;
        RECT 94.850 380.805 95.470 380.990 ;
        RECT 58.400 380.725 60.020 380.735 ;
        RECT 90.850 380.725 92.470 380.735 ;
        RECT 31.650 380.355 62.170 380.725 ;
        RECT 64.100 380.355 94.620 380.725 ;
        RECT 31.650 379.635 62.170 380.015 ;
        RECT 64.100 379.635 94.620 380.015 ;
        RECT 30.800 379.380 31.420 379.565 ;
        RECT 62.400 379.380 63.020 379.565 ;
        RECT 30.800 379.150 63.020 379.380 ;
        RECT 30.800 378.965 31.420 379.150 ;
        RECT 62.400 378.965 63.020 379.150 ;
        RECT 63.250 379.380 63.870 379.565 ;
        RECT 94.850 379.380 95.470 379.565 ;
        RECT 63.250 379.150 95.470 379.380 ;
        RECT 63.250 378.965 63.870 379.150 ;
        RECT 94.850 378.965 95.470 379.150 ;
        RECT 54.560 378.885 56.180 378.895 ;
        RECT 87.010 378.885 88.630 378.895 ;
        RECT 31.650 378.515 62.170 378.885 ;
        RECT 64.100 378.515 94.620 378.885 ;
        RECT 31.660 377.720 62.160 378.160 ;
        RECT 64.110 377.720 94.610 378.160 ;
        RECT 31.650 376.990 62.170 377.370 ;
        RECT 64.100 376.990 94.620 377.370 ;
        RECT 30.800 376.735 31.420 376.920 ;
        RECT 62.400 376.735 63.020 376.920 ;
        RECT 30.800 376.505 63.020 376.735 ;
        RECT 30.800 376.320 31.420 376.505 ;
        RECT 62.400 376.320 63.020 376.505 ;
        RECT 63.250 376.735 63.870 376.920 ;
        RECT 94.850 376.735 95.470 376.920 ;
        RECT 63.250 376.505 95.470 376.735 ;
        RECT 63.250 376.320 63.870 376.505 ;
        RECT 94.850 376.320 95.470 376.505 ;
        RECT 50.720 376.240 52.340 376.250 ;
        RECT 83.170 376.240 84.790 376.250 ;
        RECT 31.650 375.870 62.170 376.240 ;
        RECT 64.100 375.870 94.620 376.240 ;
        RECT 31.650 375.150 62.170 375.530 ;
        RECT 64.100 375.150 94.620 375.530 ;
        RECT 30.800 374.895 31.420 375.080 ;
        RECT 62.400 374.895 63.020 375.080 ;
        RECT 30.800 374.665 63.020 374.895 ;
        RECT 30.800 374.480 31.420 374.665 ;
        RECT 62.400 374.480 63.020 374.665 ;
        RECT 63.250 374.895 63.870 375.080 ;
        RECT 94.850 374.895 95.470 375.080 ;
        RECT 63.250 374.665 95.470 374.895 ;
        RECT 63.250 374.480 63.870 374.665 ;
        RECT 94.850 374.480 95.470 374.665 ;
        RECT 46.880 374.400 48.500 374.410 ;
        RECT 79.330 374.400 80.950 374.410 ;
        RECT 31.650 374.030 62.170 374.400 ;
        RECT 64.100 374.030 94.620 374.400 ;
        RECT 31.650 373.310 62.170 373.690 ;
        RECT 64.100 373.310 94.620 373.690 ;
        RECT 30.800 373.055 31.420 373.240 ;
        RECT 62.400 373.055 63.020 373.240 ;
        RECT 30.800 372.825 63.020 373.055 ;
        RECT 30.800 372.640 31.420 372.825 ;
        RECT 62.400 372.640 63.020 372.825 ;
        RECT 63.250 373.055 63.870 373.240 ;
        RECT 94.850 373.055 95.470 373.240 ;
        RECT 63.250 372.825 95.470 373.055 ;
        RECT 63.250 372.640 63.870 372.825 ;
        RECT 94.850 372.640 95.470 372.825 ;
        RECT 43.040 372.560 44.660 372.570 ;
        RECT 75.490 372.560 77.110 372.570 ;
        RECT 31.650 372.190 62.170 372.560 ;
        RECT 64.100 372.190 94.620 372.560 ;
        RECT 31.660 371.395 62.160 371.835 ;
        RECT 64.110 371.395 94.610 371.835 ;
        RECT 31.650 370.665 62.170 371.045 ;
        RECT 64.100 370.665 94.620 371.045 ;
        RECT 30.800 370.410 31.420 370.595 ;
        RECT 62.400 370.410 63.020 370.595 ;
        RECT 30.800 370.180 63.020 370.410 ;
        RECT 30.800 369.995 31.420 370.180 ;
        RECT 62.400 369.995 63.020 370.180 ;
        RECT 63.250 370.410 63.870 370.595 ;
        RECT 94.850 370.410 95.470 370.595 ;
        RECT 63.250 370.180 95.470 370.410 ;
        RECT 63.250 369.995 63.870 370.180 ;
        RECT 94.850 369.995 95.470 370.180 ;
        RECT 39.200 369.915 40.820 369.925 ;
        RECT 71.650 369.915 73.270 369.925 ;
        RECT 31.650 369.545 62.170 369.915 ;
        RECT 64.100 369.545 94.620 369.915 ;
        RECT 31.650 368.825 62.170 369.205 ;
        RECT 64.100 368.825 94.620 369.205 ;
        RECT 30.800 368.570 31.420 368.755 ;
        RECT 62.400 368.570 63.020 368.755 ;
        RECT 30.800 368.340 63.020 368.570 ;
        RECT 30.800 368.155 31.420 368.340 ;
        RECT 62.400 368.155 63.020 368.340 ;
        RECT 63.250 368.570 63.870 368.755 ;
        RECT 94.850 368.570 95.470 368.755 ;
        RECT 63.250 368.340 95.470 368.570 ;
        RECT 63.250 368.155 63.870 368.340 ;
        RECT 94.850 368.155 95.470 368.340 ;
        RECT 35.360 368.075 36.980 368.085 ;
        RECT 67.810 368.075 69.430 368.085 ;
        RECT 31.650 367.705 62.170 368.075 ;
        RECT 64.100 367.705 94.620 368.075 ;
        RECT 31.650 366.985 62.170 367.365 ;
        RECT 64.100 366.985 94.620 367.365 ;
        RECT 30.800 366.730 31.420 366.915 ;
        RECT 62.400 366.730 63.020 366.915 ;
        RECT 30.800 366.500 63.020 366.730 ;
        RECT 30.800 366.315 31.420 366.500 ;
        RECT 62.400 366.315 63.020 366.500 ;
        RECT 63.250 366.730 63.870 366.915 ;
        RECT 94.850 366.730 95.470 366.915 ;
        RECT 63.250 366.500 95.470 366.730 ;
        RECT 63.250 366.315 63.870 366.500 ;
        RECT 94.850 366.315 95.470 366.500 ;
        RECT 31.650 365.865 62.170 366.235 ;
        RECT 64.100 365.865 94.620 366.235 ;
        RECT 25.090 363.515 27.380 363.855 ;
        RECT 28.125 363.515 29.610 363.855 ;
        RECT 25.090 362.880 25.690 363.515 ;
        RECT 25.090 362.650 26.670 362.880 ;
        RECT 25.090 360.610 25.690 362.650 ;
        RECT 27.100 362.420 27.460 362.505 ;
        RECT 25.970 362.190 27.460 362.420 ;
        RECT 25.970 362.040 26.330 362.190 ;
        RECT 25.920 361.405 26.870 361.810 ;
        RECT 25.090 360.380 26.380 360.610 ;
        RECT 25.090 359.420 25.690 360.380 ;
        RECT 26.610 360.060 26.870 361.405 ;
        RECT 27.100 360.755 27.460 362.190 ;
        RECT 27.690 360.855 28.040 362.055 ;
        RECT 28.400 361.445 28.780 363.090 ;
        RECT 27.480 360.060 27.830 360.120 ;
        RECT 28.400 360.060 28.740 360.665 ;
        RECT 26.610 359.800 28.740 360.060 ;
        RECT 27.480 359.740 27.830 359.800 ;
        RECT 29.010 359.520 29.610 363.515 ;
        RECT 31.455 363.080 33.205 365.865 ;
        RECT 33.845 363.080 34.655 364.080 ;
        RECT 35.295 363.080 37.045 365.375 ;
        RECT 37.685 363.080 38.495 364.080 ;
        RECT 39.135 363.080 40.885 365.375 ;
        RECT 41.525 363.080 42.335 364.080 ;
        RECT 42.975 363.080 44.725 365.375 ;
        RECT 45.365 363.080 46.175 364.080 ;
        RECT 46.815 363.080 48.565 365.375 ;
        RECT 49.205 363.080 50.015 364.080 ;
        RECT 50.655 363.080 52.405 365.375 ;
        RECT 53.045 363.080 53.855 364.080 ;
        RECT 54.495 363.080 56.245 365.375 ;
        RECT 56.885 363.080 57.695 364.080 ;
        RECT 58.335 363.080 60.085 365.375 ;
        RECT 60.725 363.080 61.535 364.080 ;
        RECT 63.905 363.080 65.655 365.865 ;
        RECT 66.295 363.080 67.105 364.080 ;
        RECT 67.745 363.080 69.495 365.375 ;
        RECT 70.135 363.080 70.945 364.080 ;
        RECT 71.585 363.080 73.335 365.375 ;
        RECT 73.975 363.080 74.785 364.080 ;
        RECT 75.425 363.080 77.175 365.375 ;
        RECT 77.815 363.080 78.625 364.080 ;
        RECT 79.265 363.080 81.015 365.375 ;
        RECT 81.655 363.080 82.465 364.080 ;
        RECT 83.105 363.080 84.855 365.375 ;
        RECT 85.495 363.080 86.305 364.080 ;
        RECT 86.945 363.080 88.695 365.375 ;
        RECT 89.335 363.080 90.145 364.080 ;
        RECT 90.785 363.080 92.535 365.375 ;
        RECT 93.175 363.080 93.985 364.080 ;
        RECT 96.400 363.270 96.770 381.780 ;
        RECT 97.420 378.145 97.790 381.780 ;
        RECT 97.415 377.765 97.795 378.145 ;
        RECT 97.420 375.145 97.790 377.765 ;
        RECT 97.415 374.765 97.795 375.145 ;
        RECT 97.420 372.145 97.790 374.765 ;
        RECT 97.415 371.765 97.795 372.145 ;
        RECT 97.420 369.145 97.790 371.765 ;
        RECT 97.415 368.765 97.795 369.145 ;
        RECT 97.420 366.145 97.790 368.765 ;
        RECT 97.415 365.765 97.795 366.145 ;
        RECT 96.400 362.890 96.780 363.270 ;
        RECT 96.400 361.820 96.770 362.890 ;
        RECT 31.925 360.630 32.735 361.630 ;
        RECT 25.090 359.190 26.780 359.420 ;
        RECT 28.150 359.290 29.610 359.520 ;
        RECT 25.090 357.180 25.690 359.190 ;
        RECT 27.110 358.730 28.110 359.055 ;
        RECT 25.920 358.170 28.780 358.500 ;
        RECT 25.090 356.950 26.780 357.180 ;
        RECT 25.090 354.940 25.690 356.950 ;
        RECT 27.495 356.815 27.760 358.170 ;
        RECT 29.010 357.280 29.610 359.290 ;
        RECT 33.375 358.800 35.125 361.630 ;
        RECT 35.765 360.630 36.575 361.630 ;
        RECT 37.215 359.335 38.965 361.630 ;
        RECT 39.605 360.630 40.415 361.630 ;
        RECT 41.055 359.335 42.805 361.630 ;
        RECT 43.445 360.630 44.255 361.630 ;
        RECT 44.895 359.335 46.645 361.630 ;
        RECT 47.285 360.630 48.095 361.630 ;
        RECT 48.735 359.335 50.485 361.630 ;
        RECT 51.125 360.630 51.935 361.630 ;
        RECT 52.575 359.335 54.325 361.630 ;
        RECT 54.965 360.630 55.775 361.630 ;
        RECT 56.415 359.335 58.165 361.630 ;
        RECT 58.805 360.630 59.615 361.630 ;
        RECT 60.255 359.335 62.005 361.630 ;
        RECT 64.375 360.630 65.185 361.630 ;
        RECT 65.825 358.800 67.575 361.630 ;
        RECT 68.215 360.630 69.025 361.630 ;
        RECT 69.665 359.335 71.415 361.630 ;
        RECT 72.055 360.630 72.865 361.630 ;
        RECT 73.505 359.335 75.255 361.630 ;
        RECT 75.895 360.630 76.705 361.630 ;
        RECT 77.345 359.335 79.095 361.630 ;
        RECT 79.735 360.630 80.545 361.630 ;
        RECT 81.185 359.335 82.935 361.630 ;
        RECT 83.575 360.630 84.385 361.630 ;
        RECT 85.025 359.335 86.775 361.630 ;
        RECT 87.415 360.630 88.225 361.630 ;
        RECT 88.865 359.335 90.615 361.630 ;
        RECT 91.255 360.630 92.065 361.630 ;
        RECT 92.705 359.335 94.455 361.630 ;
        RECT 96.400 361.440 96.780 361.820 ;
        RECT 31.650 358.430 62.170 358.800 ;
        RECT 64.100 358.430 94.620 358.800 ;
        RECT 30.800 358.165 31.420 358.350 ;
        RECT 62.400 358.165 63.020 358.350 ;
        RECT 30.800 357.935 63.020 358.165 ;
        RECT 30.800 357.750 31.420 357.935 ;
        RECT 62.400 357.750 63.020 357.935 ;
        RECT 63.250 358.165 63.870 358.350 ;
        RECT 94.850 358.165 95.470 358.350 ;
        RECT 63.250 357.935 95.470 358.165 ;
        RECT 63.250 357.750 63.870 357.935 ;
        RECT 94.850 357.750 95.470 357.935 ;
        RECT 31.650 357.300 62.170 357.680 ;
        RECT 64.100 357.300 94.620 357.680 ;
        RECT 28.150 357.050 29.610 357.280 ;
        RECT 27.110 356.490 28.110 356.815 ;
        RECT 25.920 355.930 28.780 356.260 ;
        RECT 29.010 355.040 29.610 357.050 ;
        RECT 31.650 356.590 62.170 356.960 ;
        RECT 64.100 356.590 94.620 356.960 ;
        RECT 37.280 356.580 38.900 356.590 ;
        RECT 69.730 356.580 71.350 356.590 ;
        RECT 30.800 356.325 31.420 356.510 ;
        RECT 62.400 356.325 63.020 356.510 ;
        RECT 30.800 356.095 63.020 356.325 ;
        RECT 30.800 355.910 31.420 356.095 ;
        RECT 62.400 355.910 63.020 356.095 ;
        RECT 63.250 356.325 63.870 356.510 ;
        RECT 94.850 356.325 95.470 356.510 ;
        RECT 63.250 356.095 95.470 356.325 ;
        RECT 63.250 355.910 63.870 356.095 ;
        RECT 94.850 355.910 95.470 356.095 ;
        RECT 31.650 355.460 62.170 355.840 ;
        RECT 64.100 355.460 94.620 355.840 ;
        RECT 25.090 354.710 26.780 354.940 ;
        RECT 28.150 354.810 29.610 355.040 ;
        RECT 25.090 352.655 25.690 354.710 ;
        RECT 27.110 354.250 28.110 354.575 ;
        RECT 29.010 352.655 29.610 354.810 ;
        RECT 31.650 354.745 62.170 355.115 ;
        RECT 64.100 354.745 94.620 355.115 ;
        RECT 41.120 354.735 42.740 354.745 ;
        RECT 73.570 354.735 75.190 354.745 ;
        RECT 30.800 354.480 31.420 354.665 ;
        RECT 62.400 354.480 63.020 354.665 ;
        RECT 30.800 354.250 63.020 354.480 ;
        RECT 30.800 354.065 31.420 354.250 ;
        RECT 62.400 354.065 63.020 354.250 ;
        RECT 63.250 354.480 63.870 354.665 ;
        RECT 94.850 354.480 95.470 354.665 ;
        RECT 63.250 354.250 95.470 354.480 ;
        RECT 63.250 354.065 63.870 354.250 ;
        RECT 94.850 354.065 95.470 354.250 ;
        RECT 31.650 353.615 62.170 353.995 ;
        RECT 64.100 353.615 94.620 353.995 ;
        RECT 31.660 352.825 62.160 353.265 ;
        RECT 64.110 352.825 94.610 353.265 ;
        RECT 25.090 352.315 27.380 352.655 ;
        RECT 28.125 352.315 29.610 352.655 ;
        RECT 25.090 324.470 25.690 352.315 ;
        RECT 29.010 324.470 29.610 352.315 ;
        RECT 31.650 352.105 62.170 352.475 ;
        RECT 64.100 352.105 94.620 352.475 ;
        RECT 44.960 352.095 46.580 352.105 ;
        RECT 77.410 352.095 79.030 352.105 ;
        RECT 30.800 351.840 31.420 352.025 ;
        RECT 62.400 351.840 63.020 352.025 ;
        RECT 30.800 351.610 63.020 351.840 ;
        RECT 30.800 351.425 31.420 351.610 ;
        RECT 62.400 351.425 63.020 351.610 ;
        RECT 63.250 351.840 63.870 352.025 ;
        RECT 94.850 351.840 95.470 352.025 ;
        RECT 63.250 351.610 95.470 351.840 ;
        RECT 63.250 351.425 63.870 351.610 ;
        RECT 94.850 351.425 95.470 351.610 ;
        RECT 31.650 350.975 62.170 351.355 ;
        RECT 64.100 350.975 94.620 351.355 ;
        RECT 31.650 350.265 62.170 350.635 ;
        RECT 64.100 350.265 94.620 350.635 ;
        RECT 48.800 350.255 50.420 350.265 ;
        RECT 81.250 350.255 82.870 350.265 ;
        RECT 30.800 350.000 31.420 350.185 ;
        RECT 62.400 350.000 63.020 350.185 ;
        RECT 30.800 349.770 63.020 350.000 ;
        RECT 30.800 349.585 31.420 349.770 ;
        RECT 62.400 349.585 63.020 349.770 ;
        RECT 63.250 350.000 63.870 350.185 ;
        RECT 94.850 350.000 95.470 350.185 ;
        RECT 63.250 349.770 95.470 350.000 ;
        RECT 63.250 349.585 63.870 349.770 ;
        RECT 94.850 349.585 95.470 349.770 ;
        RECT 31.650 349.135 62.170 349.515 ;
        RECT 64.100 349.135 94.620 349.515 ;
        RECT 31.650 348.420 62.170 348.790 ;
        RECT 64.100 348.420 94.620 348.790 ;
        RECT 52.640 348.410 54.260 348.420 ;
        RECT 85.090 348.410 86.710 348.420 ;
        RECT 30.800 348.155 31.420 348.340 ;
        RECT 62.400 348.155 63.020 348.340 ;
        RECT 30.800 347.925 63.020 348.155 ;
        RECT 30.800 347.740 31.420 347.925 ;
        RECT 62.400 347.740 63.020 347.925 ;
        RECT 63.250 348.155 63.870 348.340 ;
        RECT 94.850 348.155 95.470 348.340 ;
        RECT 63.250 347.925 95.470 348.155 ;
        RECT 63.250 347.740 63.870 347.925 ;
        RECT 94.850 347.740 95.470 347.925 ;
        RECT 31.650 347.290 62.170 347.670 ;
        RECT 64.100 347.290 94.620 347.670 ;
        RECT 31.660 346.500 62.160 346.940 ;
        RECT 64.110 346.500 94.610 346.940 ;
        RECT 31.650 345.780 62.170 346.150 ;
        RECT 64.100 345.780 94.620 346.150 ;
        RECT 56.480 345.770 58.100 345.780 ;
        RECT 88.930 345.770 90.550 345.780 ;
        RECT 30.800 345.515 31.420 345.700 ;
        RECT 62.400 345.515 63.020 345.700 ;
        RECT 30.800 345.285 63.020 345.515 ;
        RECT 30.800 345.100 31.420 345.285 ;
        RECT 62.400 345.100 63.020 345.285 ;
        RECT 63.250 345.515 63.870 345.700 ;
        RECT 94.850 345.515 95.470 345.700 ;
        RECT 63.250 345.285 95.470 345.515 ;
        RECT 63.250 345.100 63.870 345.285 ;
        RECT 94.850 345.100 95.470 345.285 ;
        RECT 31.650 344.650 62.170 345.030 ;
        RECT 64.100 344.650 94.620 345.030 ;
        RECT 31.650 343.940 62.170 344.310 ;
        RECT 64.100 343.940 94.620 344.310 ;
        RECT 60.320 343.930 61.940 343.940 ;
        RECT 92.770 343.930 94.390 343.940 ;
        RECT 30.800 343.675 31.420 343.860 ;
        RECT 62.400 343.675 63.020 343.860 ;
        RECT 30.800 343.445 63.020 343.675 ;
        RECT 30.800 343.260 31.420 343.445 ;
        RECT 62.400 343.260 63.020 343.445 ;
        RECT 63.250 343.675 63.870 343.860 ;
        RECT 94.850 343.675 95.470 343.860 ;
        RECT 63.250 343.445 95.470 343.675 ;
        RECT 96.400 343.510 96.770 361.440 ;
        RECT 97.420 360.145 97.790 365.765 ;
        RECT 98.440 363.270 98.810 381.780 ;
        RECT 99.460 378.145 99.830 381.780 ;
        RECT 99.455 377.765 99.835 378.145 ;
        RECT 99.460 375.145 99.830 377.765 ;
        RECT 99.455 374.765 99.835 375.145 ;
        RECT 99.460 372.145 99.830 374.765 ;
        RECT 99.455 371.765 99.835 372.145 ;
        RECT 99.460 369.145 99.830 371.765 ;
        RECT 99.455 368.765 99.835 369.145 ;
        RECT 99.460 366.145 99.830 368.765 ;
        RECT 99.455 365.765 99.835 366.145 ;
        RECT 98.440 362.890 98.820 363.270 ;
        RECT 98.440 361.820 98.810 362.890 ;
        RECT 98.440 361.440 98.820 361.820 ;
        RECT 97.415 359.765 97.795 360.145 ;
        RECT 97.420 357.145 97.790 359.765 ;
        RECT 97.415 356.765 97.795 357.145 ;
        RECT 97.420 354.145 97.790 356.765 ;
        RECT 97.415 353.765 97.795 354.145 ;
        RECT 97.420 351.145 97.790 353.765 ;
        RECT 97.415 350.765 97.795 351.145 ;
        RECT 97.420 348.145 97.790 350.765 ;
        RECT 97.415 347.765 97.795 348.145 ;
        RECT 97.420 345.145 97.790 347.765 ;
        RECT 97.415 344.765 97.795 345.145 ;
        RECT 97.420 343.510 97.790 344.765 ;
        RECT 98.440 343.510 98.810 361.440 ;
        RECT 99.460 360.145 99.830 365.765 ;
        RECT 99.455 359.765 99.835 360.145 ;
        RECT 99.460 357.145 99.830 359.765 ;
        RECT 99.455 356.765 99.835 357.145 ;
        RECT 99.460 354.145 99.830 356.765 ;
        RECT 99.455 353.765 99.835 354.145 ;
        RECT 99.460 351.145 99.830 353.765 ;
        RECT 99.455 350.765 99.835 351.145 ;
        RECT 99.460 348.145 99.830 350.765 ;
        RECT 99.455 347.765 99.835 348.145 ;
        RECT 99.460 345.145 99.830 347.765 ;
        RECT 99.455 344.765 99.835 345.145 ;
        RECT 99.460 343.510 99.830 344.765 ;
        RECT 100.480 343.510 100.860 381.780 ;
        RECT 101.210 343.520 101.650 381.770 ;
        RECT 63.250 343.260 63.870 343.445 ;
        RECT 94.850 343.260 95.470 343.445 ;
        RECT 31.650 342.810 62.170 343.190 ;
        RECT 64.100 342.810 94.620 343.190 ;
        RECT 31.650 342.090 62.170 342.470 ;
        RECT 64.100 342.090 94.620 342.470 ;
        RECT 30.800 341.835 31.420 342.020 ;
        RECT 62.400 341.835 63.020 342.020 ;
        RECT 30.800 341.605 63.020 341.835 ;
        RECT 30.800 341.420 31.420 341.605 ;
        RECT 62.400 341.420 63.020 341.605 ;
        RECT 63.250 341.835 63.870 342.020 ;
        RECT 94.850 341.835 95.470 342.020 ;
        RECT 63.250 341.605 95.470 341.835 ;
        RECT 63.250 341.420 63.870 341.605 ;
        RECT 94.850 341.420 95.470 341.605 ;
        RECT 58.400 341.340 60.020 341.350 ;
        RECT 90.850 341.340 92.470 341.350 ;
        RECT 31.650 340.970 62.170 341.340 ;
        RECT 64.100 340.970 94.620 341.340 ;
        RECT 31.650 340.250 62.170 340.630 ;
        RECT 64.100 340.250 94.620 340.630 ;
        RECT 30.800 339.995 31.420 340.180 ;
        RECT 62.400 339.995 63.020 340.180 ;
        RECT 30.800 339.765 63.020 339.995 ;
        RECT 30.800 339.580 31.420 339.765 ;
        RECT 62.400 339.580 63.020 339.765 ;
        RECT 63.250 339.995 63.870 340.180 ;
        RECT 94.850 339.995 95.470 340.180 ;
        RECT 63.250 339.765 95.470 339.995 ;
        RECT 63.250 339.580 63.870 339.765 ;
        RECT 94.850 339.580 95.470 339.765 ;
        RECT 54.560 339.500 56.180 339.510 ;
        RECT 87.010 339.500 88.630 339.510 ;
        RECT 31.650 339.130 62.170 339.500 ;
        RECT 64.100 339.130 94.620 339.500 ;
        RECT 31.660 338.335 62.160 338.775 ;
        RECT 64.110 338.335 94.610 338.775 ;
        RECT 31.650 337.605 62.170 337.985 ;
        RECT 64.100 337.605 94.620 337.985 ;
        RECT 30.800 337.350 31.420 337.535 ;
        RECT 62.400 337.350 63.020 337.535 ;
        RECT 30.800 337.120 63.020 337.350 ;
        RECT 30.800 336.935 31.420 337.120 ;
        RECT 62.400 336.935 63.020 337.120 ;
        RECT 63.250 337.350 63.870 337.535 ;
        RECT 94.850 337.350 95.470 337.535 ;
        RECT 63.250 337.120 95.470 337.350 ;
        RECT 63.250 336.935 63.870 337.120 ;
        RECT 94.850 336.935 95.470 337.120 ;
        RECT 50.720 336.855 52.340 336.865 ;
        RECT 83.170 336.855 84.790 336.865 ;
        RECT 31.650 336.485 62.170 336.855 ;
        RECT 64.100 336.485 94.620 336.855 ;
        RECT 31.650 335.765 62.170 336.145 ;
        RECT 64.100 335.765 94.620 336.145 ;
        RECT 30.800 335.510 31.420 335.695 ;
        RECT 62.400 335.510 63.020 335.695 ;
        RECT 30.800 335.280 63.020 335.510 ;
        RECT 30.800 335.095 31.420 335.280 ;
        RECT 62.400 335.095 63.020 335.280 ;
        RECT 63.250 335.510 63.870 335.695 ;
        RECT 94.850 335.510 95.470 335.695 ;
        RECT 63.250 335.280 95.470 335.510 ;
        RECT 63.250 335.095 63.870 335.280 ;
        RECT 94.850 335.095 95.470 335.280 ;
        RECT 46.880 335.015 48.500 335.025 ;
        RECT 79.330 335.015 80.950 335.025 ;
        RECT 31.650 334.645 62.170 335.015 ;
        RECT 64.100 334.645 94.620 335.015 ;
        RECT 31.650 333.925 62.170 334.305 ;
        RECT 64.100 333.925 94.620 334.305 ;
        RECT 30.800 333.670 31.420 333.855 ;
        RECT 62.400 333.670 63.020 333.855 ;
        RECT 30.800 333.440 63.020 333.670 ;
        RECT 30.800 333.255 31.420 333.440 ;
        RECT 62.400 333.255 63.020 333.440 ;
        RECT 63.250 333.670 63.870 333.855 ;
        RECT 94.850 333.670 95.470 333.855 ;
        RECT 63.250 333.440 95.470 333.670 ;
        RECT 63.250 333.255 63.870 333.440 ;
        RECT 94.850 333.255 95.470 333.440 ;
        RECT 43.040 333.175 44.660 333.185 ;
        RECT 75.490 333.175 77.110 333.185 ;
        RECT 31.650 332.805 62.170 333.175 ;
        RECT 64.100 332.805 94.620 333.175 ;
        RECT 31.660 332.010 62.160 332.450 ;
        RECT 64.110 332.010 94.610 332.450 ;
        RECT 31.650 331.280 62.170 331.660 ;
        RECT 64.100 331.280 94.620 331.660 ;
        RECT 30.800 331.025 31.420 331.210 ;
        RECT 62.400 331.025 63.020 331.210 ;
        RECT 30.800 330.795 63.020 331.025 ;
        RECT 30.800 330.610 31.420 330.795 ;
        RECT 62.400 330.610 63.020 330.795 ;
        RECT 63.250 331.025 63.870 331.210 ;
        RECT 94.850 331.025 95.470 331.210 ;
        RECT 63.250 330.795 95.470 331.025 ;
        RECT 63.250 330.610 63.870 330.795 ;
        RECT 94.850 330.610 95.470 330.795 ;
        RECT 39.200 330.530 40.820 330.540 ;
        RECT 71.650 330.530 73.270 330.540 ;
        RECT 31.650 330.160 62.170 330.530 ;
        RECT 64.100 330.160 94.620 330.530 ;
        RECT 31.650 329.440 62.170 329.820 ;
        RECT 64.100 329.440 94.620 329.820 ;
        RECT 30.800 329.185 31.420 329.370 ;
        RECT 62.400 329.185 63.020 329.370 ;
        RECT 30.800 328.955 63.020 329.185 ;
        RECT 30.800 328.770 31.420 328.955 ;
        RECT 62.400 328.770 63.020 328.955 ;
        RECT 63.250 329.185 63.870 329.370 ;
        RECT 94.850 329.185 95.470 329.370 ;
        RECT 63.250 328.955 95.470 329.185 ;
        RECT 63.250 328.770 63.870 328.955 ;
        RECT 94.850 328.770 95.470 328.955 ;
        RECT 35.360 328.690 36.980 328.700 ;
        RECT 67.810 328.690 69.430 328.700 ;
        RECT 31.650 328.320 62.170 328.690 ;
        RECT 64.100 328.320 94.620 328.690 ;
        RECT 31.650 327.600 62.170 327.980 ;
        RECT 64.100 327.600 94.620 327.980 ;
        RECT 30.800 327.345 31.420 327.530 ;
        RECT 62.400 327.345 63.020 327.530 ;
        RECT 30.800 327.115 63.020 327.345 ;
        RECT 30.800 326.930 31.420 327.115 ;
        RECT 62.400 326.930 63.020 327.115 ;
        RECT 63.250 327.345 63.870 327.530 ;
        RECT 94.850 327.345 95.470 327.530 ;
        RECT 63.250 327.115 95.470 327.345 ;
        RECT 63.250 326.930 63.870 327.115 ;
        RECT 94.850 326.930 95.470 327.115 ;
        RECT 31.650 326.480 62.170 326.850 ;
        RECT 64.100 326.480 94.620 326.850 ;
        RECT 25.090 324.130 27.380 324.470 ;
        RECT 28.125 324.130 29.610 324.470 ;
        RECT 25.090 323.495 25.690 324.130 ;
        RECT 25.090 323.265 26.670 323.495 ;
        RECT 25.090 321.225 25.690 323.265 ;
        RECT 27.100 323.035 27.460 323.120 ;
        RECT 25.970 322.805 27.460 323.035 ;
        RECT 25.970 322.655 26.330 322.805 ;
        RECT 25.920 322.020 26.870 322.425 ;
        RECT 25.090 320.995 26.380 321.225 ;
        RECT 25.090 320.035 25.690 320.995 ;
        RECT 26.610 320.675 26.870 322.020 ;
        RECT 27.100 321.370 27.460 322.805 ;
        RECT 27.690 321.470 28.040 322.670 ;
        RECT 28.400 322.060 28.780 323.705 ;
        RECT 27.480 320.675 27.830 320.735 ;
        RECT 28.400 320.675 28.740 321.280 ;
        RECT 26.610 320.415 28.740 320.675 ;
        RECT 27.480 320.355 27.830 320.415 ;
        RECT 29.010 320.135 29.610 324.130 ;
        RECT 31.455 323.695 33.205 326.480 ;
        RECT 33.845 323.695 34.655 324.695 ;
        RECT 35.295 323.695 37.045 325.990 ;
        RECT 37.685 323.695 38.495 324.695 ;
        RECT 39.135 323.695 40.885 325.990 ;
        RECT 41.525 323.695 42.335 324.695 ;
        RECT 42.975 323.695 44.725 325.990 ;
        RECT 45.365 323.695 46.175 324.695 ;
        RECT 46.815 323.695 48.565 325.990 ;
        RECT 49.205 323.695 50.015 324.695 ;
        RECT 50.655 323.695 52.405 325.990 ;
        RECT 53.045 323.695 53.855 324.695 ;
        RECT 54.495 323.695 56.245 325.990 ;
        RECT 56.885 323.695 57.695 324.695 ;
        RECT 58.335 323.695 60.085 325.990 ;
        RECT 60.725 323.695 61.535 324.695 ;
        RECT 63.905 323.695 65.655 326.480 ;
        RECT 66.295 323.695 67.105 324.695 ;
        RECT 67.745 323.695 69.495 325.990 ;
        RECT 70.135 323.695 70.945 324.695 ;
        RECT 71.585 323.695 73.335 325.990 ;
        RECT 73.975 323.695 74.785 324.695 ;
        RECT 75.425 323.695 77.175 325.990 ;
        RECT 77.815 323.695 78.625 324.695 ;
        RECT 79.265 323.695 81.015 325.990 ;
        RECT 81.655 323.695 82.465 324.695 ;
        RECT 83.105 323.695 84.855 325.990 ;
        RECT 85.495 323.695 86.305 324.695 ;
        RECT 86.945 323.695 88.695 325.990 ;
        RECT 89.335 323.695 90.145 324.695 ;
        RECT 90.785 323.695 92.535 325.990 ;
        RECT 93.175 323.695 93.985 324.695 ;
        RECT 96.400 323.885 96.770 342.395 ;
        RECT 97.420 338.760 97.790 342.395 ;
        RECT 97.415 338.380 97.795 338.760 ;
        RECT 97.420 335.760 97.790 338.380 ;
        RECT 97.415 335.380 97.795 335.760 ;
        RECT 97.420 332.760 97.790 335.380 ;
        RECT 97.415 332.380 97.795 332.760 ;
        RECT 97.420 329.760 97.790 332.380 ;
        RECT 97.415 329.380 97.795 329.760 ;
        RECT 97.420 326.760 97.790 329.380 ;
        RECT 97.415 326.380 97.795 326.760 ;
        RECT 96.400 323.505 96.780 323.885 ;
        RECT 96.400 322.435 96.770 323.505 ;
        RECT 31.925 321.245 32.735 322.245 ;
        RECT 25.090 319.805 26.780 320.035 ;
        RECT 28.150 319.905 29.610 320.135 ;
        RECT 25.090 317.795 25.690 319.805 ;
        RECT 27.110 319.345 28.110 319.670 ;
        RECT 25.920 318.785 28.780 319.115 ;
        RECT 25.090 317.565 26.780 317.795 ;
        RECT 25.090 315.555 25.690 317.565 ;
        RECT 27.495 317.430 27.760 318.785 ;
        RECT 29.010 317.895 29.610 319.905 ;
        RECT 33.375 319.415 35.125 322.245 ;
        RECT 35.765 321.245 36.575 322.245 ;
        RECT 37.215 319.950 38.965 322.245 ;
        RECT 39.605 321.245 40.415 322.245 ;
        RECT 41.055 319.950 42.805 322.245 ;
        RECT 43.445 321.245 44.255 322.245 ;
        RECT 44.895 319.950 46.645 322.245 ;
        RECT 47.285 321.245 48.095 322.245 ;
        RECT 48.735 319.950 50.485 322.245 ;
        RECT 51.125 321.245 51.935 322.245 ;
        RECT 52.575 319.950 54.325 322.245 ;
        RECT 54.965 321.245 55.775 322.245 ;
        RECT 56.415 319.950 58.165 322.245 ;
        RECT 58.805 321.245 59.615 322.245 ;
        RECT 60.255 319.950 62.005 322.245 ;
        RECT 64.375 321.245 65.185 322.245 ;
        RECT 65.825 319.415 67.575 322.245 ;
        RECT 68.215 321.245 69.025 322.245 ;
        RECT 69.665 319.950 71.415 322.245 ;
        RECT 72.055 321.245 72.865 322.245 ;
        RECT 73.505 319.950 75.255 322.245 ;
        RECT 75.895 321.245 76.705 322.245 ;
        RECT 77.345 319.950 79.095 322.245 ;
        RECT 79.735 321.245 80.545 322.245 ;
        RECT 81.185 319.950 82.935 322.245 ;
        RECT 83.575 321.245 84.385 322.245 ;
        RECT 85.025 319.950 86.775 322.245 ;
        RECT 87.415 321.245 88.225 322.245 ;
        RECT 88.865 319.950 90.615 322.245 ;
        RECT 91.255 321.245 92.065 322.245 ;
        RECT 92.705 319.950 94.455 322.245 ;
        RECT 96.400 322.055 96.780 322.435 ;
        RECT 31.650 319.045 62.170 319.415 ;
        RECT 64.100 319.045 94.620 319.415 ;
        RECT 30.800 318.780 31.420 318.965 ;
        RECT 62.400 318.780 63.020 318.965 ;
        RECT 30.800 318.550 63.020 318.780 ;
        RECT 30.800 318.365 31.420 318.550 ;
        RECT 62.400 318.365 63.020 318.550 ;
        RECT 63.250 318.780 63.870 318.965 ;
        RECT 94.850 318.780 95.470 318.965 ;
        RECT 63.250 318.550 95.470 318.780 ;
        RECT 63.250 318.365 63.870 318.550 ;
        RECT 94.850 318.365 95.470 318.550 ;
        RECT 31.650 317.915 62.170 318.295 ;
        RECT 64.100 317.915 94.620 318.295 ;
        RECT 28.150 317.665 29.610 317.895 ;
        RECT 27.110 317.105 28.110 317.430 ;
        RECT 25.920 316.545 28.780 316.875 ;
        RECT 29.010 315.655 29.610 317.665 ;
        RECT 31.650 317.205 62.170 317.575 ;
        RECT 64.100 317.205 94.620 317.575 ;
        RECT 37.280 317.195 38.900 317.205 ;
        RECT 69.730 317.195 71.350 317.205 ;
        RECT 30.800 316.940 31.420 317.125 ;
        RECT 62.400 316.940 63.020 317.125 ;
        RECT 30.800 316.710 63.020 316.940 ;
        RECT 30.800 316.525 31.420 316.710 ;
        RECT 62.400 316.525 63.020 316.710 ;
        RECT 63.250 316.940 63.870 317.125 ;
        RECT 94.850 316.940 95.470 317.125 ;
        RECT 63.250 316.710 95.470 316.940 ;
        RECT 63.250 316.525 63.870 316.710 ;
        RECT 94.850 316.525 95.470 316.710 ;
        RECT 31.650 316.075 62.170 316.455 ;
        RECT 64.100 316.075 94.620 316.455 ;
        RECT 25.090 315.325 26.780 315.555 ;
        RECT 28.150 315.425 29.610 315.655 ;
        RECT 25.090 313.270 25.690 315.325 ;
        RECT 27.110 314.865 28.110 315.190 ;
        RECT 29.010 313.270 29.610 315.425 ;
        RECT 31.650 315.360 62.170 315.730 ;
        RECT 64.100 315.360 94.620 315.730 ;
        RECT 41.120 315.350 42.740 315.360 ;
        RECT 73.570 315.350 75.190 315.360 ;
        RECT 30.800 315.095 31.420 315.280 ;
        RECT 62.400 315.095 63.020 315.280 ;
        RECT 30.800 314.865 63.020 315.095 ;
        RECT 30.800 314.680 31.420 314.865 ;
        RECT 62.400 314.680 63.020 314.865 ;
        RECT 63.250 315.095 63.870 315.280 ;
        RECT 94.850 315.095 95.470 315.280 ;
        RECT 63.250 314.865 95.470 315.095 ;
        RECT 63.250 314.680 63.870 314.865 ;
        RECT 94.850 314.680 95.470 314.865 ;
        RECT 31.650 314.230 62.170 314.610 ;
        RECT 64.100 314.230 94.620 314.610 ;
        RECT 31.660 313.440 62.160 313.880 ;
        RECT 64.110 313.440 94.610 313.880 ;
        RECT 25.090 312.930 27.380 313.270 ;
        RECT 28.125 312.930 29.610 313.270 ;
        RECT 25.090 285.085 25.690 312.930 ;
        RECT 29.010 285.085 29.610 312.930 ;
        RECT 31.650 312.720 62.170 313.090 ;
        RECT 64.100 312.720 94.620 313.090 ;
        RECT 44.960 312.710 46.580 312.720 ;
        RECT 77.410 312.710 79.030 312.720 ;
        RECT 30.800 312.455 31.420 312.640 ;
        RECT 62.400 312.455 63.020 312.640 ;
        RECT 30.800 312.225 63.020 312.455 ;
        RECT 30.800 312.040 31.420 312.225 ;
        RECT 62.400 312.040 63.020 312.225 ;
        RECT 63.250 312.455 63.870 312.640 ;
        RECT 94.850 312.455 95.470 312.640 ;
        RECT 63.250 312.225 95.470 312.455 ;
        RECT 63.250 312.040 63.870 312.225 ;
        RECT 94.850 312.040 95.470 312.225 ;
        RECT 31.650 311.590 62.170 311.970 ;
        RECT 64.100 311.590 94.620 311.970 ;
        RECT 31.650 310.880 62.170 311.250 ;
        RECT 64.100 310.880 94.620 311.250 ;
        RECT 48.800 310.870 50.420 310.880 ;
        RECT 81.250 310.870 82.870 310.880 ;
        RECT 30.800 310.615 31.420 310.800 ;
        RECT 62.400 310.615 63.020 310.800 ;
        RECT 30.800 310.385 63.020 310.615 ;
        RECT 30.800 310.200 31.420 310.385 ;
        RECT 62.400 310.200 63.020 310.385 ;
        RECT 63.250 310.615 63.870 310.800 ;
        RECT 94.850 310.615 95.470 310.800 ;
        RECT 63.250 310.385 95.470 310.615 ;
        RECT 63.250 310.200 63.870 310.385 ;
        RECT 94.850 310.200 95.470 310.385 ;
        RECT 31.650 309.750 62.170 310.130 ;
        RECT 64.100 309.750 94.620 310.130 ;
        RECT 31.650 309.035 62.170 309.405 ;
        RECT 64.100 309.035 94.620 309.405 ;
        RECT 52.640 309.025 54.260 309.035 ;
        RECT 85.090 309.025 86.710 309.035 ;
        RECT 30.800 308.770 31.420 308.955 ;
        RECT 62.400 308.770 63.020 308.955 ;
        RECT 30.800 308.540 63.020 308.770 ;
        RECT 30.800 308.355 31.420 308.540 ;
        RECT 62.400 308.355 63.020 308.540 ;
        RECT 63.250 308.770 63.870 308.955 ;
        RECT 94.850 308.770 95.470 308.955 ;
        RECT 63.250 308.540 95.470 308.770 ;
        RECT 63.250 308.355 63.870 308.540 ;
        RECT 94.850 308.355 95.470 308.540 ;
        RECT 31.650 307.905 62.170 308.285 ;
        RECT 64.100 307.905 94.620 308.285 ;
        RECT 31.660 307.115 62.160 307.555 ;
        RECT 64.110 307.115 94.610 307.555 ;
        RECT 31.650 306.395 62.170 306.765 ;
        RECT 64.100 306.395 94.620 306.765 ;
        RECT 56.480 306.385 58.100 306.395 ;
        RECT 88.930 306.385 90.550 306.395 ;
        RECT 30.800 306.130 31.420 306.315 ;
        RECT 62.400 306.130 63.020 306.315 ;
        RECT 30.800 305.900 63.020 306.130 ;
        RECT 30.800 305.715 31.420 305.900 ;
        RECT 62.400 305.715 63.020 305.900 ;
        RECT 63.250 306.130 63.870 306.315 ;
        RECT 94.850 306.130 95.470 306.315 ;
        RECT 63.250 305.900 95.470 306.130 ;
        RECT 63.250 305.715 63.870 305.900 ;
        RECT 94.850 305.715 95.470 305.900 ;
        RECT 31.650 305.265 62.170 305.645 ;
        RECT 64.100 305.265 94.620 305.645 ;
        RECT 31.650 304.555 62.170 304.925 ;
        RECT 64.100 304.555 94.620 304.925 ;
        RECT 60.320 304.545 61.940 304.555 ;
        RECT 92.770 304.545 94.390 304.555 ;
        RECT 30.800 304.290 31.420 304.475 ;
        RECT 62.400 304.290 63.020 304.475 ;
        RECT 30.800 304.060 63.020 304.290 ;
        RECT 30.800 303.875 31.420 304.060 ;
        RECT 62.400 303.875 63.020 304.060 ;
        RECT 63.250 304.290 63.870 304.475 ;
        RECT 94.850 304.290 95.470 304.475 ;
        RECT 63.250 304.060 95.470 304.290 ;
        RECT 96.400 304.125 96.770 322.055 ;
        RECT 97.420 320.760 97.790 326.380 ;
        RECT 98.440 323.885 98.810 342.395 ;
        RECT 99.460 338.760 99.830 342.395 ;
        RECT 99.455 338.380 99.835 338.760 ;
        RECT 99.460 335.760 99.830 338.380 ;
        RECT 99.455 335.380 99.835 335.760 ;
        RECT 99.460 332.760 99.830 335.380 ;
        RECT 99.455 332.380 99.835 332.760 ;
        RECT 99.460 329.760 99.830 332.380 ;
        RECT 99.455 329.380 99.835 329.760 ;
        RECT 99.460 326.760 99.830 329.380 ;
        RECT 99.455 326.380 99.835 326.760 ;
        RECT 98.440 323.505 98.820 323.885 ;
        RECT 98.440 322.435 98.810 323.505 ;
        RECT 98.440 322.055 98.820 322.435 ;
        RECT 97.415 320.380 97.795 320.760 ;
        RECT 97.420 317.760 97.790 320.380 ;
        RECT 97.415 317.380 97.795 317.760 ;
        RECT 97.420 314.760 97.790 317.380 ;
        RECT 97.415 314.380 97.795 314.760 ;
        RECT 97.420 311.760 97.790 314.380 ;
        RECT 97.415 311.380 97.795 311.760 ;
        RECT 97.420 308.760 97.790 311.380 ;
        RECT 97.415 308.380 97.795 308.760 ;
        RECT 97.420 305.760 97.790 308.380 ;
        RECT 97.415 305.380 97.795 305.760 ;
        RECT 97.420 304.125 97.790 305.380 ;
        RECT 98.440 304.125 98.810 322.055 ;
        RECT 99.460 320.760 99.830 326.380 ;
        RECT 99.455 320.380 99.835 320.760 ;
        RECT 99.460 317.760 99.830 320.380 ;
        RECT 99.455 317.380 99.835 317.760 ;
        RECT 99.460 314.760 99.830 317.380 ;
        RECT 99.455 314.380 99.835 314.760 ;
        RECT 99.460 311.760 99.830 314.380 ;
        RECT 99.455 311.380 99.835 311.760 ;
        RECT 99.460 308.760 99.830 311.380 ;
        RECT 99.455 308.380 99.835 308.760 ;
        RECT 99.460 305.760 99.830 308.380 ;
        RECT 99.455 305.380 99.835 305.760 ;
        RECT 99.460 304.125 99.830 305.380 ;
        RECT 100.480 304.125 100.860 342.395 ;
        RECT 101.210 304.135 101.650 342.385 ;
        RECT 63.250 303.875 63.870 304.060 ;
        RECT 94.850 303.875 95.470 304.060 ;
        RECT 31.650 303.425 62.170 303.805 ;
        RECT 64.100 303.425 94.620 303.805 ;
        RECT 31.650 302.705 62.170 303.085 ;
        RECT 64.100 302.705 94.620 303.085 ;
        RECT 30.800 302.450 31.420 302.635 ;
        RECT 62.400 302.450 63.020 302.635 ;
        RECT 30.800 302.220 63.020 302.450 ;
        RECT 30.800 302.035 31.420 302.220 ;
        RECT 62.400 302.035 63.020 302.220 ;
        RECT 63.250 302.450 63.870 302.635 ;
        RECT 94.850 302.450 95.470 302.635 ;
        RECT 63.250 302.220 95.470 302.450 ;
        RECT 63.250 302.035 63.870 302.220 ;
        RECT 94.850 302.035 95.470 302.220 ;
        RECT 58.400 301.955 60.020 301.965 ;
        RECT 90.850 301.955 92.470 301.965 ;
        RECT 31.650 301.585 62.170 301.955 ;
        RECT 64.100 301.585 94.620 301.955 ;
        RECT 31.650 300.865 62.170 301.245 ;
        RECT 64.100 300.865 94.620 301.245 ;
        RECT 30.800 300.610 31.420 300.795 ;
        RECT 62.400 300.610 63.020 300.795 ;
        RECT 30.800 300.380 63.020 300.610 ;
        RECT 30.800 300.195 31.420 300.380 ;
        RECT 62.400 300.195 63.020 300.380 ;
        RECT 63.250 300.610 63.870 300.795 ;
        RECT 94.850 300.610 95.470 300.795 ;
        RECT 63.250 300.380 95.470 300.610 ;
        RECT 63.250 300.195 63.870 300.380 ;
        RECT 94.850 300.195 95.470 300.380 ;
        RECT 54.560 300.115 56.180 300.125 ;
        RECT 87.010 300.115 88.630 300.125 ;
        RECT 31.650 299.745 62.170 300.115 ;
        RECT 64.100 299.745 94.620 300.115 ;
        RECT 31.660 298.950 62.160 299.390 ;
        RECT 64.110 298.950 94.610 299.390 ;
        RECT 31.650 298.220 62.170 298.600 ;
        RECT 64.100 298.220 94.620 298.600 ;
        RECT 30.800 297.965 31.420 298.150 ;
        RECT 62.400 297.965 63.020 298.150 ;
        RECT 30.800 297.735 63.020 297.965 ;
        RECT 30.800 297.550 31.420 297.735 ;
        RECT 62.400 297.550 63.020 297.735 ;
        RECT 63.250 297.965 63.870 298.150 ;
        RECT 94.850 297.965 95.470 298.150 ;
        RECT 63.250 297.735 95.470 297.965 ;
        RECT 63.250 297.550 63.870 297.735 ;
        RECT 94.850 297.550 95.470 297.735 ;
        RECT 50.720 297.470 52.340 297.480 ;
        RECT 83.170 297.470 84.790 297.480 ;
        RECT 31.650 297.100 62.170 297.470 ;
        RECT 64.100 297.100 94.620 297.470 ;
        RECT 31.650 296.380 62.170 296.760 ;
        RECT 64.100 296.380 94.620 296.760 ;
        RECT 30.800 296.125 31.420 296.310 ;
        RECT 62.400 296.125 63.020 296.310 ;
        RECT 30.800 295.895 63.020 296.125 ;
        RECT 30.800 295.710 31.420 295.895 ;
        RECT 62.400 295.710 63.020 295.895 ;
        RECT 63.250 296.125 63.870 296.310 ;
        RECT 94.850 296.125 95.470 296.310 ;
        RECT 63.250 295.895 95.470 296.125 ;
        RECT 63.250 295.710 63.870 295.895 ;
        RECT 94.850 295.710 95.470 295.895 ;
        RECT 46.880 295.630 48.500 295.640 ;
        RECT 79.330 295.630 80.950 295.640 ;
        RECT 31.650 295.260 62.170 295.630 ;
        RECT 64.100 295.260 94.620 295.630 ;
        RECT 31.650 294.540 62.170 294.920 ;
        RECT 64.100 294.540 94.620 294.920 ;
        RECT 30.800 294.285 31.420 294.470 ;
        RECT 62.400 294.285 63.020 294.470 ;
        RECT 30.800 294.055 63.020 294.285 ;
        RECT 30.800 293.870 31.420 294.055 ;
        RECT 62.400 293.870 63.020 294.055 ;
        RECT 63.250 294.285 63.870 294.470 ;
        RECT 94.850 294.285 95.470 294.470 ;
        RECT 63.250 294.055 95.470 294.285 ;
        RECT 63.250 293.870 63.870 294.055 ;
        RECT 94.850 293.870 95.470 294.055 ;
        RECT 43.040 293.790 44.660 293.800 ;
        RECT 75.490 293.790 77.110 293.800 ;
        RECT 31.650 293.420 62.170 293.790 ;
        RECT 64.100 293.420 94.620 293.790 ;
        RECT 31.660 292.625 62.160 293.065 ;
        RECT 64.110 292.625 94.610 293.065 ;
        RECT 31.650 291.895 62.170 292.275 ;
        RECT 64.100 291.895 94.620 292.275 ;
        RECT 30.800 291.640 31.420 291.825 ;
        RECT 62.400 291.640 63.020 291.825 ;
        RECT 30.800 291.410 63.020 291.640 ;
        RECT 30.800 291.225 31.420 291.410 ;
        RECT 62.400 291.225 63.020 291.410 ;
        RECT 63.250 291.640 63.870 291.825 ;
        RECT 94.850 291.640 95.470 291.825 ;
        RECT 63.250 291.410 95.470 291.640 ;
        RECT 63.250 291.225 63.870 291.410 ;
        RECT 94.850 291.225 95.470 291.410 ;
        RECT 39.200 291.145 40.820 291.155 ;
        RECT 71.650 291.145 73.270 291.155 ;
        RECT 31.650 290.775 62.170 291.145 ;
        RECT 64.100 290.775 94.620 291.145 ;
        RECT 31.650 290.055 62.170 290.435 ;
        RECT 64.100 290.055 94.620 290.435 ;
        RECT 30.800 289.800 31.420 289.985 ;
        RECT 62.400 289.800 63.020 289.985 ;
        RECT 30.800 289.570 63.020 289.800 ;
        RECT 30.800 289.385 31.420 289.570 ;
        RECT 62.400 289.385 63.020 289.570 ;
        RECT 63.250 289.800 63.870 289.985 ;
        RECT 94.850 289.800 95.470 289.985 ;
        RECT 63.250 289.570 95.470 289.800 ;
        RECT 63.250 289.385 63.870 289.570 ;
        RECT 94.850 289.385 95.470 289.570 ;
        RECT 35.360 289.305 36.980 289.315 ;
        RECT 67.810 289.305 69.430 289.315 ;
        RECT 31.650 288.935 62.170 289.305 ;
        RECT 64.100 288.935 94.620 289.305 ;
        RECT 31.650 288.215 62.170 288.595 ;
        RECT 64.100 288.215 94.620 288.595 ;
        RECT 30.800 287.960 31.420 288.145 ;
        RECT 62.400 287.960 63.020 288.145 ;
        RECT 30.800 287.730 63.020 287.960 ;
        RECT 30.800 287.545 31.420 287.730 ;
        RECT 62.400 287.545 63.020 287.730 ;
        RECT 63.250 287.960 63.870 288.145 ;
        RECT 94.850 287.960 95.470 288.145 ;
        RECT 63.250 287.730 95.470 287.960 ;
        RECT 63.250 287.545 63.870 287.730 ;
        RECT 94.850 287.545 95.470 287.730 ;
        RECT 31.650 287.095 62.170 287.465 ;
        RECT 64.100 287.095 94.620 287.465 ;
        RECT 25.090 284.745 27.380 285.085 ;
        RECT 28.125 284.745 29.610 285.085 ;
        RECT 25.090 284.110 25.690 284.745 ;
        RECT 25.090 283.880 26.670 284.110 ;
        RECT 25.090 281.840 25.690 283.880 ;
        RECT 27.100 283.650 27.460 283.735 ;
        RECT 25.970 283.420 27.460 283.650 ;
        RECT 25.970 283.270 26.330 283.420 ;
        RECT 25.920 282.635 26.870 283.040 ;
        RECT 25.090 281.610 26.380 281.840 ;
        RECT 25.090 280.650 25.690 281.610 ;
        RECT 26.610 281.290 26.870 282.635 ;
        RECT 27.100 281.985 27.460 283.420 ;
        RECT 27.690 282.085 28.040 283.285 ;
        RECT 28.400 282.675 28.780 284.320 ;
        RECT 27.480 281.290 27.830 281.350 ;
        RECT 28.400 281.290 28.740 281.895 ;
        RECT 26.610 281.030 28.740 281.290 ;
        RECT 27.480 280.970 27.830 281.030 ;
        RECT 29.010 280.750 29.610 284.745 ;
        RECT 31.455 284.310 33.205 287.095 ;
        RECT 33.845 284.310 34.655 285.310 ;
        RECT 35.295 284.310 37.045 286.605 ;
        RECT 37.685 284.310 38.495 285.310 ;
        RECT 39.135 284.310 40.885 286.605 ;
        RECT 41.525 284.310 42.335 285.310 ;
        RECT 42.975 284.310 44.725 286.605 ;
        RECT 45.365 284.310 46.175 285.310 ;
        RECT 46.815 284.310 48.565 286.605 ;
        RECT 49.205 284.310 50.015 285.310 ;
        RECT 50.655 284.310 52.405 286.605 ;
        RECT 53.045 284.310 53.855 285.310 ;
        RECT 54.495 284.310 56.245 286.605 ;
        RECT 56.885 284.310 57.695 285.310 ;
        RECT 58.335 284.310 60.085 286.605 ;
        RECT 60.725 284.310 61.535 285.310 ;
        RECT 63.905 284.310 65.655 287.095 ;
        RECT 66.295 284.310 67.105 285.310 ;
        RECT 67.745 284.310 69.495 286.605 ;
        RECT 70.135 284.310 70.945 285.310 ;
        RECT 71.585 284.310 73.335 286.605 ;
        RECT 73.975 284.310 74.785 285.310 ;
        RECT 75.425 284.310 77.175 286.605 ;
        RECT 77.815 284.310 78.625 285.310 ;
        RECT 79.265 284.310 81.015 286.605 ;
        RECT 81.655 284.310 82.465 285.310 ;
        RECT 83.105 284.310 84.855 286.605 ;
        RECT 85.495 284.310 86.305 285.310 ;
        RECT 86.945 284.310 88.695 286.605 ;
        RECT 89.335 284.310 90.145 285.310 ;
        RECT 90.785 284.310 92.535 286.605 ;
        RECT 93.175 284.310 93.985 285.310 ;
        RECT 96.400 284.500 96.770 303.010 ;
        RECT 97.420 299.375 97.790 303.010 ;
        RECT 97.415 298.995 97.795 299.375 ;
        RECT 97.420 296.375 97.790 298.995 ;
        RECT 97.415 295.995 97.795 296.375 ;
        RECT 97.420 293.375 97.790 295.995 ;
        RECT 97.415 292.995 97.795 293.375 ;
        RECT 97.420 290.375 97.790 292.995 ;
        RECT 97.415 289.995 97.795 290.375 ;
        RECT 97.420 287.375 97.790 289.995 ;
        RECT 97.415 286.995 97.795 287.375 ;
        RECT 96.400 284.120 96.780 284.500 ;
        RECT 96.400 283.050 96.770 284.120 ;
        RECT 31.925 281.860 32.735 282.860 ;
        RECT 25.090 280.420 26.780 280.650 ;
        RECT 28.150 280.520 29.610 280.750 ;
        RECT 25.090 278.410 25.690 280.420 ;
        RECT 27.110 279.960 28.110 280.285 ;
        RECT 25.920 279.400 28.780 279.730 ;
        RECT 25.090 278.180 26.780 278.410 ;
        RECT 25.090 276.170 25.690 278.180 ;
        RECT 27.495 278.045 27.760 279.400 ;
        RECT 29.010 278.510 29.610 280.520 ;
        RECT 33.375 280.030 35.125 282.860 ;
        RECT 35.765 281.860 36.575 282.860 ;
        RECT 37.215 280.565 38.965 282.860 ;
        RECT 39.605 281.860 40.415 282.860 ;
        RECT 41.055 280.565 42.805 282.860 ;
        RECT 43.445 281.860 44.255 282.860 ;
        RECT 44.895 280.565 46.645 282.860 ;
        RECT 47.285 281.860 48.095 282.860 ;
        RECT 48.735 280.565 50.485 282.860 ;
        RECT 51.125 281.860 51.935 282.860 ;
        RECT 52.575 280.565 54.325 282.860 ;
        RECT 54.965 281.860 55.775 282.860 ;
        RECT 56.415 280.565 58.165 282.860 ;
        RECT 58.805 281.860 59.615 282.860 ;
        RECT 60.255 280.565 62.005 282.860 ;
        RECT 64.375 281.860 65.185 282.860 ;
        RECT 65.825 280.030 67.575 282.860 ;
        RECT 68.215 281.860 69.025 282.860 ;
        RECT 69.665 280.565 71.415 282.860 ;
        RECT 72.055 281.860 72.865 282.860 ;
        RECT 73.505 280.565 75.255 282.860 ;
        RECT 75.895 281.860 76.705 282.860 ;
        RECT 77.345 280.565 79.095 282.860 ;
        RECT 79.735 281.860 80.545 282.860 ;
        RECT 81.185 280.565 82.935 282.860 ;
        RECT 83.575 281.860 84.385 282.860 ;
        RECT 85.025 280.565 86.775 282.860 ;
        RECT 87.415 281.860 88.225 282.860 ;
        RECT 88.865 280.565 90.615 282.860 ;
        RECT 91.255 281.860 92.065 282.860 ;
        RECT 92.705 280.565 94.455 282.860 ;
        RECT 96.400 282.670 96.780 283.050 ;
        RECT 31.650 279.660 62.170 280.030 ;
        RECT 64.100 279.660 94.620 280.030 ;
        RECT 30.800 279.395 31.420 279.580 ;
        RECT 62.400 279.395 63.020 279.580 ;
        RECT 30.800 279.165 63.020 279.395 ;
        RECT 30.800 278.980 31.420 279.165 ;
        RECT 62.400 278.980 63.020 279.165 ;
        RECT 63.250 279.395 63.870 279.580 ;
        RECT 94.850 279.395 95.470 279.580 ;
        RECT 63.250 279.165 95.470 279.395 ;
        RECT 63.250 278.980 63.870 279.165 ;
        RECT 94.850 278.980 95.470 279.165 ;
        RECT 31.650 278.530 62.170 278.910 ;
        RECT 64.100 278.530 94.620 278.910 ;
        RECT 28.150 278.280 29.610 278.510 ;
        RECT 27.110 277.720 28.110 278.045 ;
        RECT 25.920 277.160 28.780 277.490 ;
        RECT 29.010 276.270 29.610 278.280 ;
        RECT 31.650 277.820 62.170 278.190 ;
        RECT 64.100 277.820 94.620 278.190 ;
        RECT 37.280 277.810 38.900 277.820 ;
        RECT 69.730 277.810 71.350 277.820 ;
        RECT 30.800 277.555 31.420 277.740 ;
        RECT 62.400 277.555 63.020 277.740 ;
        RECT 30.800 277.325 63.020 277.555 ;
        RECT 30.800 277.140 31.420 277.325 ;
        RECT 62.400 277.140 63.020 277.325 ;
        RECT 63.250 277.555 63.870 277.740 ;
        RECT 94.850 277.555 95.470 277.740 ;
        RECT 63.250 277.325 95.470 277.555 ;
        RECT 63.250 277.140 63.870 277.325 ;
        RECT 94.850 277.140 95.470 277.325 ;
        RECT 31.650 276.690 62.170 277.070 ;
        RECT 64.100 276.690 94.620 277.070 ;
        RECT 25.090 275.940 26.780 276.170 ;
        RECT 28.150 276.040 29.610 276.270 ;
        RECT 25.090 273.885 25.690 275.940 ;
        RECT 27.110 275.480 28.110 275.805 ;
        RECT 29.010 273.885 29.610 276.040 ;
        RECT 31.650 275.975 62.170 276.345 ;
        RECT 64.100 275.975 94.620 276.345 ;
        RECT 41.120 275.965 42.740 275.975 ;
        RECT 73.570 275.965 75.190 275.975 ;
        RECT 30.800 275.710 31.420 275.895 ;
        RECT 62.400 275.710 63.020 275.895 ;
        RECT 30.800 275.480 63.020 275.710 ;
        RECT 30.800 275.295 31.420 275.480 ;
        RECT 62.400 275.295 63.020 275.480 ;
        RECT 63.250 275.710 63.870 275.895 ;
        RECT 94.850 275.710 95.470 275.895 ;
        RECT 63.250 275.480 95.470 275.710 ;
        RECT 63.250 275.295 63.870 275.480 ;
        RECT 94.850 275.295 95.470 275.480 ;
        RECT 31.650 274.845 62.170 275.225 ;
        RECT 64.100 274.845 94.620 275.225 ;
        RECT 31.660 274.055 62.160 274.495 ;
        RECT 64.110 274.055 94.610 274.495 ;
        RECT 25.090 273.545 27.380 273.885 ;
        RECT 28.125 273.545 29.610 273.885 ;
        RECT 25.090 245.700 25.690 273.545 ;
        RECT 29.010 245.700 29.610 273.545 ;
        RECT 31.650 273.335 62.170 273.705 ;
        RECT 64.100 273.335 94.620 273.705 ;
        RECT 44.960 273.325 46.580 273.335 ;
        RECT 77.410 273.325 79.030 273.335 ;
        RECT 30.800 273.070 31.420 273.255 ;
        RECT 62.400 273.070 63.020 273.255 ;
        RECT 30.800 272.840 63.020 273.070 ;
        RECT 30.800 272.655 31.420 272.840 ;
        RECT 62.400 272.655 63.020 272.840 ;
        RECT 63.250 273.070 63.870 273.255 ;
        RECT 94.850 273.070 95.470 273.255 ;
        RECT 63.250 272.840 95.470 273.070 ;
        RECT 63.250 272.655 63.870 272.840 ;
        RECT 94.850 272.655 95.470 272.840 ;
        RECT 31.650 272.205 62.170 272.585 ;
        RECT 64.100 272.205 94.620 272.585 ;
        RECT 31.650 271.495 62.170 271.865 ;
        RECT 64.100 271.495 94.620 271.865 ;
        RECT 48.800 271.485 50.420 271.495 ;
        RECT 81.250 271.485 82.870 271.495 ;
        RECT 30.800 271.230 31.420 271.415 ;
        RECT 62.400 271.230 63.020 271.415 ;
        RECT 30.800 271.000 63.020 271.230 ;
        RECT 30.800 270.815 31.420 271.000 ;
        RECT 62.400 270.815 63.020 271.000 ;
        RECT 63.250 271.230 63.870 271.415 ;
        RECT 94.850 271.230 95.470 271.415 ;
        RECT 63.250 271.000 95.470 271.230 ;
        RECT 63.250 270.815 63.870 271.000 ;
        RECT 94.850 270.815 95.470 271.000 ;
        RECT 31.650 270.365 62.170 270.745 ;
        RECT 64.100 270.365 94.620 270.745 ;
        RECT 31.650 269.650 62.170 270.020 ;
        RECT 64.100 269.650 94.620 270.020 ;
        RECT 52.640 269.640 54.260 269.650 ;
        RECT 85.090 269.640 86.710 269.650 ;
        RECT 30.800 269.385 31.420 269.570 ;
        RECT 62.400 269.385 63.020 269.570 ;
        RECT 30.800 269.155 63.020 269.385 ;
        RECT 30.800 268.970 31.420 269.155 ;
        RECT 62.400 268.970 63.020 269.155 ;
        RECT 63.250 269.385 63.870 269.570 ;
        RECT 94.850 269.385 95.470 269.570 ;
        RECT 63.250 269.155 95.470 269.385 ;
        RECT 63.250 268.970 63.870 269.155 ;
        RECT 94.850 268.970 95.470 269.155 ;
        RECT 31.650 268.520 62.170 268.900 ;
        RECT 64.100 268.520 94.620 268.900 ;
        RECT 31.660 267.730 62.160 268.170 ;
        RECT 64.110 267.730 94.610 268.170 ;
        RECT 31.650 267.010 62.170 267.380 ;
        RECT 64.100 267.010 94.620 267.380 ;
        RECT 56.480 267.000 58.100 267.010 ;
        RECT 88.930 267.000 90.550 267.010 ;
        RECT 30.800 266.745 31.420 266.930 ;
        RECT 62.400 266.745 63.020 266.930 ;
        RECT 30.800 266.515 63.020 266.745 ;
        RECT 30.800 266.330 31.420 266.515 ;
        RECT 62.400 266.330 63.020 266.515 ;
        RECT 63.250 266.745 63.870 266.930 ;
        RECT 94.850 266.745 95.470 266.930 ;
        RECT 63.250 266.515 95.470 266.745 ;
        RECT 63.250 266.330 63.870 266.515 ;
        RECT 94.850 266.330 95.470 266.515 ;
        RECT 31.650 265.880 62.170 266.260 ;
        RECT 64.100 265.880 94.620 266.260 ;
        RECT 31.650 265.170 62.170 265.540 ;
        RECT 64.100 265.170 94.620 265.540 ;
        RECT 60.320 265.160 61.940 265.170 ;
        RECT 92.770 265.160 94.390 265.170 ;
        RECT 30.800 264.905 31.420 265.090 ;
        RECT 62.400 264.905 63.020 265.090 ;
        RECT 30.800 264.675 63.020 264.905 ;
        RECT 30.800 264.490 31.420 264.675 ;
        RECT 62.400 264.490 63.020 264.675 ;
        RECT 63.250 264.905 63.870 265.090 ;
        RECT 94.850 264.905 95.470 265.090 ;
        RECT 63.250 264.675 95.470 264.905 ;
        RECT 96.400 264.740 96.770 282.670 ;
        RECT 97.420 281.375 97.790 286.995 ;
        RECT 98.440 284.500 98.810 303.010 ;
        RECT 99.460 299.375 99.830 303.010 ;
        RECT 99.455 298.995 99.835 299.375 ;
        RECT 99.460 296.375 99.830 298.995 ;
        RECT 99.455 295.995 99.835 296.375 ;
        RECT 99.460 293.375 99.830 295.995 ;
        RECT 99.455 292.995 99.835 293.375 ;
        RECT 99.460 290.375 99.830 292.995 ;
        RECT 99.455 289.995 99.835 290.375 ;
        RECT 99.460 287.375 99.830 289.995 ;
        RECT 99.455 286.995 99.835 287.375 ;
        RECT 98.440 284.120 98.820 284.500 ;
        RECT 98.440 283.050 98.810 284.120 ;
        RECT 98.440 282.670 98.820 283.050 ;
        RECT 97.415 280.995 97.795 281.375 ;
        RECT 97.420 278.375 97.790 280.995 ;
        RECT 97.415 277.995 97.795 278.375 ;
        RECT 97.420 275.375 97.790 277.995 ;
        RECT 97.415 274.995 97.795 275.375 ;
        RECT 97.420 272.375 97.790 274.995 ;
        RECT 97.415 271.995 97.795 272.375 ;
        RECT 97.420 269.375 97.790 271.995 ;
        RECT 97.415 268.995 97.795 269.375 ;
        RECT 97.420 266.375 97.790 268.995 ;
        RECT 97.415 265.995 97.795 266.375 ;
        RECT 97.420 264.740 97.790 265.995 ;
        RECT 98.440 264.740 98.810 282.670 ;
        RECT 99.460 281.375 99.830 286.995 ;
        RECT 99.455 280.995 99.835 281.375 ;
        RECT 99.460 278.375 99.830 280.995 ;
        RECT 99.455 277.995 99.835 278.375 ;
        RECT 99.460 275.375 99.830 277.995 ;
        RECT 99.455 274.995 99.835 275.375 ;
        RECT 99.460 272.375 99.830 274.995 ;
        RECT 99.455 271.995 99.835 272.375 ;
        RECT 99.460 269.375 99.830 271.995 ;
        RECT 99.455 268.995 99.835 269.375 ;
        RECT 99.460 266.375 99.830 268.995 ;
        RECT 99.455 265.995 99.835 266.375 ;
        RECT 99.460 264.740 99.830 265.995 ;
        RECT 100.480 264.740 100.860 303.010 ;
        RECT 101.210 264.750 101.650 303.000 ;
        RECT 63.250 264.490 63.870 264.675 ;
        RECT 94.850 264.490 95.470 264.675 ;
        RECT 31.650 264.040 62.170 264.420 ;
        RECT 64.100 264.040 94.620 264.420 ;
        RECT 31.650 263.320 62.170 263.700 ;
        RECT 64.100 263.320 94.620 263.700 ;
        RECT 30.800 263.065 31.420 263.250 ;
        RECT 62.400 263.065 63.020 263.250 ;
        RECT 30.800 262.835 63.020 263.065 ;
        RECT 30.800 262.650 31.420 262.835 ;
        RECT 62.400 262.650 63.020 262.835 ;
        RECT 63.250 263.065 63.870 263.250 ;
        RECT 94.850 263.065 95.470 263.250 ;
        RECT 63.250 262.835 95.470 263.065 ;
        RECT 63.250 262.650 63.870 262.835 ;
        RECT 94.850 262.650 95.470 262.835 ;
        RECT 58.400 262.570 60.020 262.580 ;
        RECT 90.850 262.570 92.470 262.580 ;
        RECT 31.650 262.200 62.170 262.570 ;
        RECT 64.100 262.200 94.620 262.570 ;
        RECT 31.650 261.480 62.170 261.860 ;
        RECT 64.100 261.480 94.620 261.860 ;
        RECT 30.800 261.225 31.420 261.410 ;
        RECT 62.400 261.225 63.020 261.410 ;
        RECT 30.800 260.995 63.020 261.225 ;
        RECT 30.800 260.810 31.420 260.995 ;
        RECT 62.400 260.810 63.020 260.995 ;
        RECT 63.250 261.225 63.870 261.410 ;
        RECT 94.850 261.225 95.470 261.410 ;
        RECT 63.250 260.995 95.470 261.225 ;
        RECT 63.250 260.810 63.870 260.995 ;
        RECT 94.850 260.810 95.470 260.995 ;
        RECT 54.560 260.730 56.180 260.740 ;
        RECT 87.010 260.730 88.630 260.740 ;
        RECT 31.650 260.360 62.170 260.730 ;
        RECT 64.100 260.360 94.620 260.730 ;
        RECT 31.660 259.565 62.160 260.005 ;
        RECT 64.110 259.565 94.610 260.005 ;
        RECT 31.650 258.835 62.170 259.215 ;
        RECT 64.100 258.835 94.620 259.215 ;
        RECT 30.800 258.580 31.420 258.765 ;
        RECT 62.400 258.580 63.020 258.765 ;
        RECT 30.800 258.350 63.020 258.580 ;
        RECT 30.800 258.165 31.420 258.350 ;
        RECT 62.400 258.165 63.020 258.350 ;
        RECT 63.250 258.580 63.870 258.765 ;
        RECT 94.850 258.580 95.470 258.765 ;
        RECT 63.250 258.350 95.470 258.580 ;
        RECT 63.250 258.165 63.870 258.350 ;
        RECT 94.850 258.165 95.470 258.350 ;
        RECT 50.720 258.085 52.340 258.095 ;
        RECT 83.170 258.085 84.790 258.095 ;
        RECT 31.650 257.715 62.170 258.085 ;
        RECT 64.100 257.715 94.620 258.085 ;
        RECT 31.650 256.995 62.170 257.375 ;
        RECT 64.100 256.995 94.620 257.375 ;
        RECT 30.800 256.740 31.420 256.925 ;
        RECT 62.400 256.740 63.020 256.925 ;
        RECT 30.800 256.510 63.020 256.740 ;
        RECT 30.800 256.325 31.420 256.510 ;
        RECT 62.400 256.325 63.020 256.510 ;
        RECT 63.250 256.740 63.870 256.925 ;
        RECT 94.850 256.740 95.470 256.925 ;
        RECT 63.250 256.510 95.470 256.740 ;
        RECT 63.250 256.325 63.870 256.510 ;
        RECT 94.850 256.325 95.470 256.510 ;
        RECT 46.880 256.245 48.500 256.255 ;
        RECT 79.330 256.245 80.950 256.255 ;
        RECT 31.650 255.875 62.170 256.245 ;
        RECT 64.100 255.875 94.620 256.245 ;
        RECT 31.650 255.155 62.170 255.535 ;
        RECT 64.100 255.155 94.620 255.535 ;
        RECT 30.800 254.900 31.420 255.085 ;
        RECT 62.400 254.900 63.020 255.085 ;
        RECT 30.800 254.670 63.020 254.900 ;
        RECT 30.800 254.485 31.420 254.670 ;
        RECT 62.400 254.485 63.020 254.670 ;
        RECT 63.250 254.900 63.870 255.085 ;
        RECT 94.850 254.900 95.470 255.085 ;
        RECT 63.250 254.670 95.470 254.900 ;
        RECT 63.250 254.485 63.870 254.670 ;
        RECT 94.850 254.485 95.470 254.670 ;
        RECT 43.040 254.405 44.660 254.415 ;
        RECT 75.490 254.405 77.110 254.415 ;
        RECT 31.650 254.035 62.170 254.405 ;
        RECT 64.100 254.035 94.620 254.405 ;
        RECT 31.660 253.240 62.160 253.680 ;
        RECT 64.110 253.240 94.610 253.680 ;
        RECT 31.650 252.510 62.170 252.890 ;
        RECT 64.100 252.510 94.620 252.890 ;
        RECT 30.800 252.255 31.420 252.440 ;
        RECT 62.400 252.255 63.020 252.440 ;
        RECT 30.800 252.025 63.020 252.255 ;
        RECT 30.800 251.840 31.420 252.025 ;
        RECT 62.400 251.840 63.020 252.025 ;
        RECT 63.250 252.255 63.870 252.440 ;
        RECT 94.850 252.255 95.470 252.440 ;
        RECT 63.250 252.025 95.470 252.255 ;
        RECT 63.250 251.840 63.870 252.025 ;
        RECT 94.850 251.840 95.470 252.025 ;
        RECT 39.200 251.760 40.820 251.770 ;
        RECT 71.650 251.760 73.270 251.770 ;
        RECT 31.650 251.390 62.170 251.760 ;
        RECT 64.100 251.390 94.620 251.760 ;
        RECT 31.650 250.670 62.170 251.050 ;
        RECT 64.100 250.670 94.620 251.050 ;
        RECT 30.800 250.415 31.420 250.600 ;
        RECT 62.400 250.415 63.020 250.600 ;
        RECT 30.800 250.185 63.020 250.415 ;
        RECT 30.800 250.000 31.420 250.185 ;
        RECT 62.400 250.000 63.020 250.185 ;
        RECT 63.250 250.415 63.870 250.600 ;
        RECT 94.850 250.415 95.470 250.600 ;
        RECT 63.250 250.185 95.470 250.415 ;
        RECT 63.250 250.000 63.870 250.185 ;
        RECT 94.850 250.000 95.470 250.185 ;
        RECT 35.360 249.920 36.980 249.930 ;
        RECT 67.810 249.920 69.430 249.930 ;
        RECT 31.650 249.550 62.170 249.920 ;
        RECT 64.100 249.550 94.620 249.920 ;
        RECT 31.650 248.830 62.170 249.210 ;
        RECT 64.100 248.830 94.620 249.210 ;
        RECT 30.800 248.575 31.420 248.760 ;
        RECT 62.400 248.575 63.020 248.760 ;
        RECT 30.800 248.345 63.020 248.575 ;
        RECT 30.800 248.160 31.420 248.345 ;
        RECT 62.400 248.160 63.020 248.345 ;
        RECT 63.250 248.575 63.870 248.760 ;
        RECT 94.850 248.575 95.470 248.760 ;
        RECT 63.250 248.345 95.470 248.575 ;
        RECT 63.250 248.160 63.870 248.345 ;
        RECT 94.850 248.160 95.470 248.345 ;
        RECT 31.650 247.710 62.170 248.080 ;
        RECT 64.100 247.710 94.620 248.080 ;
        RECT 25.090 245.360 27.380 245.700 ;
        RECT 28.125 245.360 29.610 245.700 ;
        RECT 25.090 244.725 25.690 245.360 ;
        RECT 25.090 244.495 26.670 244.725 ;
        RECT 25.090 242.455 25.690 244.495 ;
        RECT 27.100 244.265 27.460 244.350 ;
        RECT 25.970 244.035 27.460 244.265 ;
        RECT 25.970 243.885 26.330 244.035 ;
        RECT 25.920 243.250 26.870 243.655 ;
        RECT 25.090 242.225 26.380 242.455 ;
        RECT 25.090 241.265 25.690 242.225 ;
        RECT 26.610 241.905 26.870 243.250 ;
        RECT 27.100 242.600 27.460 244.035 ;
        RECT 27.690 242.700 28.040 243.900 ;
        RECT 28.400 243.290 28.780 244.935 ;
        RECT 27.480 241.905 27.830 241.965 ;
        RECT 28.400 241.905 28.740 242.510 ;
        RECT 26.610 241.645 28.740 241.905 ;
        RECT 27.480 241.585 27.830 241.645 ;
        RECT 29.010 241.365 29.610 245.360 ;
        RECT 31.455 244.925 33.205 247.710 ;
        RECT 33.845 244.925 34.655 245.925 ;
        RECT 35.295 244.925 37.045 247.220 ;
        RECT 37.685 244.925 38.495 245.925 ;
        RECT 39.135 244.925 40.885 247.220 ;
        RECT 41.525 244.925 42.335 245.925 ;
        RECT 42.975 244.925 44.725 247.220 ;
        RECT 45.365 244.925 46.175 245.925 ;
        RECT 46.815 244.925 48.565 247.220 ;
        RECT 49.205 244.925 50.015 245.925 ;
        RECT 50.655 244.925 52.405 247.220 ;
        RECT 53.045 244.925 53.855 245.925 ;
        RECT 54.495 244.925 56.245 247.220 ;
        RECT 56.885 244.925 57.695 245.925 ;
        RECT 58.335 244.925 60.085 247.220 ;
        RECT 60.725 244.925 61.535 245.925 ;
        RECT 63.905 244.925 65.655 247.710 ;
        RECT 66.295 244.925 67.105 245.925 ;
        RECT 67.745 244.925 69.495 247.220 ;
        RECT 70.135 244.925 70.945 245.925 ;
        RECT 71.585 244.925 73.335 247.220 ;
        RECT 73.975 244.925 74.785 245.925 ;
        RECT 75.425 244.925 77.175 247.220 ;
        RECT 77.815 244.925 78.625 245.925 ;
        RECT 79.265 244.925 81.015 247.220 ;
        RECT 81.655 244.925 82.465 245.925 ;
        RECT 83.105 244.925 84.855 247.220 ;
        RECT 85.495 244.925 86.305 245.925 ;
        RECT 86.945 244.925 88.695 247.220 ;
        RECT 89.335 244.925 90.145 245.925 ;
        RECT 90.785 244.925 92.535 247.220 ;
        RECT 93.175 244.925 93.985 245.925 ;
        RECT 96.400 245.115 96.770 263.625 ;
        RECT 97.420 259.990 97.790 263.625 ;
        RECT 97.415 259.610 97.795 259.990 ;
        RECT 97.420 256.990 97.790 259.610 ;
        RECT 97.415 256.610 97.795 256.990 ;
        RECT 97.420 253.990 97.790 256.610 ;
        RECT 97.415 253.610 97.795 253.990 ;
        RECT 97.420 250.990 97.790 253.610 ;
        RECT 97.415 250.610 97.795 250.990 ;
        RECT 97.420 247.990 97.790 250.610 ;
        RECT 97.415 247.610 97.795 247.990 ;
        RECT 96.400 244.735 96.780 245.115 ;
        RECT 96.400 243.665 96.770 244.735 ;
        RECT 31.925 242.475 32.735 243.475 ;
        RECT 25.090 241.035 26.780 241.265 ;
        RECT 28.150 241.135 29.610 241.365 ;
        RECT 25.090 239.025 25.690 241.035 ;
        RECT 27.110 240.575 28.110 240.900 ;
        RECT 25.920 240.015 28.780 240.345 ;
        RECT 25.090 238.795 26.780 239.025 ;
        RECT 25.090 236.785 25.690 238.795 ;
        RECT 27.495 238.660 27.760 240.015 ;
        RECT 29.010 239.125 29.610 241.135 ;
        RECT 33.375 240.645 35.125 243.475 ;
        RECT 35.765 242.475 36.575 243.475 ;
        RECT 37.215 241.180 38.965 243.475 ;
        RECT 39.605 242.475 40.415 243.475 ;
        RECT 41.055 241.180 42.805 243.475 ;
        RECT 43.445 242.475 44.255 243.475 ;
        RECT 44.895 241.180 46.645 243.475 ;
        RECT 47.285 242.475 48.095 243.475 ;
        RECT 48.735 241.180 50.485 243.475 ;
        RECT 51.125 242.475 51.935 243.475 ;
        RECT 52.575 241.180 54.325 243.475 ;
        RECT 54.965 242.475 55.775 243.475 ;
        RECT 56.415 241.180 58.165 243.475 ;
        RECT 58.805 242.475 59.615 243.475 ;
        RECT 60.255 241.180 62.005 243.475 ;
        RECT 64.375 242.475 65.185 243.475 ;
        RECT 65.825 240.645 67.575 243.475 ;
        RECT 68.215 242.475 69.025 243.475 ;
        RECT 69.665 241.180 71.415 243.475 ;
        RECT 72.055 242.475 72.865 243.475 ;
        RECT 73.505 241.180 75.255 243.475 ;
        RECT 75.895 242.475 76.705 243.475 ;
        RECT 77.345 241.180 79.095 243.475 ;
        RECT 79.735 242.475 80.545 243.475 ;
        RECT 81.185 241.180 82.935 243.475 ;
        RECT 83.575 242.475 84.385 243.475 ;
        RECT 85.025 241.180 86.775 243.475 ;
        RECT 87.415 242.475 88.225 243.475 ;
        RECT 88.865 241.180 90.615 243.475 ;
        RECT 91.255 242.475 92.065 243.475 ;
        RECT 92.705 241.180 94.455 243.475 ;
        RECT 96.400 243.285 96.780 243.665 ;
        RECT 31.650 240.275 62.170 240.645 ;
        RECT 64.100 240.275 94.620 240.645 ;
        RECT 30.800 240.010 31.420 240.195 ;
        RECT 62.400 240.010 63.020 240.195 ;
        RECT 30.800 239.780 63.020 240.010 ;
        RECT 30.800 239.595 31.420 239.780 ;
        RECT 62.400 239.595 63.020 239.780 ;
        RECT 63.250 240.010 63.870 240.195 ;
        RECT 94.850 240.010 95.470 240.195 ;
        RECT 63.250 239.780 95.470 240.010 ;
        RECT 63.250 239.595 63.870 239.780 ;
        RECT 94.850 239.595 95.470 239.780 ;
        RECT 31.650 239.145 62.170 239.525 ;
        RECT 64.100 239.145 94.620 239.525 ;
        RECT 28.150 238.895 29.610 239.125 ;
        RECT 27.110 238.335 28.110 238.660 ;
        RECT 25.920 237.775 28.780 238.105 ;
        RECT 29.010 236.885 29.610 238.895 ;
        RECT 31.650 238.435 62.170 238.805 ;
        RECT 64.100 238.435 94.620 238.805 ;
        RECT 37.280 238.425 38.900 238.435 ;
        RECT 69.730 238.425 71.350 238.435 ;
        RECT 30.800 238.170 31.420 238.355 ;
        RECT 62.400 238.170 63.020 238.355 ;
        RECT 30.800 237.940 63.020 238.170 ;
        RECT 30.800 237.755 31.420 237.940 ;
        RECT 62.400 237.755 63.020 237.940 ;
        RECT 63.250 238.170 63.870 238.355 ;
        RECT 94.850 238.170 95.470 238.355 ;
        RECT 63.250 237.940 95.470 238.170 ;
        RECT 63.250 237.755 63.870 237.940 ;
        RECT 94.850 237.755 95.470 237.940 ;
        RECT 31.650 237.305 62.170 237.685 ;
        RECT 64.100 237.305 94.620 237.685 ;
        RECT 25.090 236.555 26.780 236.785 ;
        RECT 28.150 236.655 29.610 236.885 ;
        RECT 25.090 234.500 25.690 236.555 ;
        RECT 27.110 236.095 28.110 236.420 ;
        RECT 29.010 234.500 29.610 236.655 ;
        RECT 31.650 236.590 62.170 236.960 ;
        RECT 64.100 236.590 94.620 236.960 ;
        RECT 41.120 236.580 42.740 236.590 ;
        RECT 73.570 236.580 75.190 236.590 ;
        RECT 30.800 236.325 31.420 236.510 ;
        RECT 62.400 236.325 63.020 236.510 ;
        RECT 30.800 236.095 63.020 236.325 ;
        RECT 30.800 235.910 31.420 236.095 ;
        RECT 62.400 235.910 63.020 236.095 ;
        RECT 63.250 236.325 63.870 236.510 ;
        RECT 94.850 236.325 95.470 236.510 ;
        RECT 63.250 236.095 95.470 236.325 ;
        RECT 63.250 235.910 63.870 236.095 ;
        RECT 94.850 235.910 95.470 236.095 ;
        RECT 31.650 235.460 62.170 235.840 ;
        RECT 64.100 235.460 94.620 235.840 ;
        RECT 31.660 234.670 62.160 235.110 ;
        RECT 64.110 234.670 94.610 235.110 ;
        RECT 25.090 234.160 27.380 234.500 ;
        RECT 28.125 234.160 29.610 234.500 ;
        RECT 25.090 206.315 25.690 234.160 ;
        RECT 29.010 206.315 29.610 234.160 ;
        RECT 31.650 233.950 62.170 234.320 ;
        RECT 64.100 233.950 94.620 234.320 ;
        RECT 44.960 233.940 46.580 233.950 ;
        RECT 77.410 233.940 79.030 233.950 ;
        RECT 30.800 233.685 31.420 233.870 ;
        RECT 62.400 233.685 63.020 233.870 ;
        RECT 30.800 233.455 63.020 233.685 ;
        RECT 30.800 233.270 31.420 233.455 ;
        RECT 62.400 233.270 63.020 233.455 ;
        RECT 63.250 233.685 63.870 233.870 ;
        RECT 94.850 233.685 95.470 233.870 ;
        RECT 63.250 233.455 95.470 233.685 ;
        RECT 63.250 233.270 63.870 233.455 ;
        RECT 94.850 233.270 95.470 233.455 ;
        RECT 31.650 232.820 62.170 233.200 ;
        RECT 64.100 232.820 94.620 233.200 ;
        RECT 31.650 232.110 62.170 232.480 ;
        RECT 64.100 232.110 94.620 232.480 ;
        RECT 48.800 232.100 50.420 232.110 ;
        RECT 81.250 232.100 82.870 232.110 ;
        RECT 30.800 231.845 31.420 232.030 ;
        RECT 62.400 231.845 63.020 232.030 ;
        RECT 30.800 231.615 63.020 231.845 ;
        RECT 30.800 231.430 31.420 231.615 ;
        RECT 62.400 231.430 63.020 231.615 ;
        RECT 63.250 231.845 63.870 232.030 ;
        RECT 94.850 231.845 95.470 232.030 ;
        RECT 63.250 231.615 95.470 231.845 ;
        RECT 63.250 231.430 63.870 231.615 ;
        RECT 94.850 231.430 95.470 231.615 ;
        RECT 31.650 230.980 62.170 231.360 ;
        RECT 64.100 230.980 94.620 231.360 ;
        RECT 31.650 230.265 62.170 230.635 ;
        RECT 64.100 230.265 94.620 230.635 ;
        RECT 52.640 230.255 54.260 230.265 ;
        RECT 85.090 230.255 86.710 230.265 ;
        RECT 30.800 230.000 31.420 230.185 ;
        RECT 62.400 230.000 63.020 230.185 ;
        RECT 30.800 229.770 63.020 230.000 ;
        RECT 30.800 229.585 31.420 229.770 ;
        RECT 62.400 229.585 63.020 229.770 ;
        RECT 63.250 230.000 63.870 230.185 ;
        RECT 94.850 230.000 95.470 230.185 ;
        RECT 63.250 229.770 95.470 230.000 ;
        RECT 63.250 229.585 63.870 229.770 ;
        RECT 94.850 229.585 95.470 229.770 ;
        RECT 31.650 229.135 62.170 229.515 ;
        RECT 64.100 229.135 94.620 229.515 ;
        RECT 31.660 228.345 62.160 228.785 ;
        RECT 64.110 228.345 94.610 228.785 ;
        RECT 31.650 227.625 62.170 227.995 ;
        RECT 64.100 227.625 94.620 227.995 ;
        RECT 56.480 227.615 58.100 227.625 ;
        RECT 88.930 227.615 90.550 227.625 ;
        RECT 30.800 227.360 31.420 227.545 ;
        RECT 62.400 227.360 63.020 227.545 ;
        RECT 30.800 227.130 63.020 227.360 ;
        RECT 30.800 226.945 31.420 227.130 ;
        RECT 62.400 226.945 63.020 227.130 ;
        RECT 63.250 227.360 63.870 227.545 ;
        RECT 94.850 227.360 95.470 227.545 ;
        RECT 63.250 227.130 95.470 227.360 ;
        RECT 63.250 226.945 63.870 227.130 ;
        RECT 94.850 226.945 95.470 227.130 ;
        RECT 31.650 226.495 62.170 226.875 ;
        RECT 64.100 226.495 94.620 226.875 ;
        RECT 31.650 225.785 62.170 226.155 ;
        RECT 64.100 225.785 94.620 226.155 ;
        RECT 60.320 225.775 61.940 225.785 ;
        RECT 92.770 225.775 94.390 225.785 ;
        RECT 30.800 225.520 31.420 225.705 ;
        RECT 62.400 225.520 63.020 225.705 ;
        RECT 30.800 225.290 63.020 225.520 ;
        RECT 30.800 225.105 31.420 225.290 ;
        RECT 62.400 225.105 63.020 225.290 ;
        RECT 63.250 225.520 63.870 225.705 ;
        RECT 94.850 225.520 95.470 225.705 ;
        RECT 63.250 225.290 95.470 225.520 ;
        RECT 96.400 225.355 96.770 243.285 ;
        RECT 97.420 241.990 97.790 247.610 ;
        RECT 98.440 245.115 98.810 263.625 ;
        RECT 99.460 259.990 99.830 263.625 ;
        RECT 99.455 259.610 99.835 259.990 ;
        RECT 99.460 256.990 99.830 259.610 ;
        RECT 99.455 256.610 99.835 256.990 ;
        RECT 99.460 253.990 99.830 256.610 ;
        RECT 99.455 253.610 99.835 253.990 ;
        RECT 99.460 250.990 99.830 253.610 ;
        RECT 99.455 250.610 99.835 250.990 ;
        RECT 99.460 247.990 99.830 250.610 ;
        RECT 99.455 247.610 99.835 247.990 ;
        RECT 98.440 244.735 98.820 245.115 ;
        RECT 98.440 243.665 98.810 244.735 ;
        RECT 98.440 243.285 98.820 243.665 ;
        RECT 97.415 241.610 97.795 241.990 ;
        RECT 97.420 238.990 97.790 241.610 ;
        RECT 97.415 238.610 97.795 238.990 ;
        RECT 97.420 235.990 97.790 238.610 ;
        RECT 97.415 235.610 97.795 235.990 ;
        RECT 97.420 232.990 97.790 235.610 ;
        RECT 97.415 232.610 97.795 232.990 ;
        RECT 97.420 229.990 97.790 232.610 ;
        RECT 97.415 229.610 97.795 229.990 ;
        RECT 97.420 226.990 97.790 229.610 ;
        RECT 97.415 226.610 97.795 226.990 ;
        RECT 97.420 225.355 97.790 226.610 ;
        RECT 98.440 225.355 98.810 243.285 ;
        RECT 99.460 241.990 99.830 247.610 ;
        RECT 99.455 241.610 99.835 241.990 ;
        RECT 99.460 238.990 99.830 241.610 ;
        RECT 99.455 238.610 99.835 238.990 ;
        RECT 99.460 235.990 99.830 238.610 ;
        RECT 99.455 235.610 99.835 235.990 ;
        RECT 99.460 232.990 99.830 235.610 ;
        RECT 99.455 232.610 99.835 232.990 ;
        RECT 99.460 229.990 99.830 232.610 ;
        RECT 99.455 229.610 99.835 229.990 ;
        RECT 99.460 226.990 99.830 229.610 ;
        RECT 99.455 226.610 99.835 226.990 ;
        RECT 99.460 225.355 99.830 226.610 ;
        RECT 100.480 225.355 100.860 263.625 ;
        RECT 101.210 225.365 101.650 263.615 ;
        RECT 63.250 225.105 63.870 225.290 ;
        RECT 94.850 225.105 95.470 225.290 ;
        RECT 31.650 224.655 62.170 225.035 ;
        RECT 64.100 224.655 94.620 225.035 ;
        RECT 31.650 223.935 62.170 224.315 ;
        RECT 64.100 223.935 94.620 224.315 ;
        RECT 30.800 223.680 31.420 223.865 ;
        RECT 62.400 223.680 63.020 223.865 ;
        RECT 30.800 223.450 63.020 223.680 ;
        RECT 30.800 223.265 31.420 223.450 ;
        RECT 62.400 223.265 63.020 223.450 ;
        RECT 63.250 223.680 63.870 223.865 ;
        RECT 94.850 223.680 95.470 223.865 ;
        RECT 63.250 223.450 95.470 223.680 ;
        RECT 63.250 223.265 63.870 223.450 ;
        RECT 94.850 223.265 95.470 223.450 ;
        RECT 58.400 223.185 60.020 223.195 ;
        RECT 90.850 223.185 92.470 223.195 ;
        RECT 31.650 222.815 62.170 223.185 ;
        RECT 64.100 222.815 94.620 223.185 ;
        RECT 31.650 222.095 62.170 222.475 ;
        RECT 64.100 222.095 94.620 222.475 ;
        RECT 30.800 221.840 31.420 222.025 ;
        RECT 62.400 221.840 63.020 222.025 ;
        RECT 30.800 221.610 63.020 221.840 ;
        RECT 30.800 221.425 31.420 221.610 ;
        RECT 62.400 221.425 63.020 221.610 ;
        RECT 63.250 221.840 63.870 222.025 ;
        RECT 94.850 221.840 95.470 222.025 ;
        RECT 63.250 221.610 95.470 221.840 ;
        RECT 63.250 221.425 63.870 221.610 ;
        RECT 94.850 221.425 95.470 221.610 ;
        RECT 54.560 221.345 56.180 221.355 ;
        RECT 87.010 221.345 88.630 221.355 ;
        RECT 31.650 220.975 62.170 221.345 ;
        RECT 64.100 220.975 94.620 221.345 ;
        RECT 31.660 220.180 62.160 220.620 ;
        RECT 64.110 220.180 94.610 220.620 ;
        RECT 31.650 219.450 62.170 219.830 ;
        RECT 64.100 219.450 94.620 219.830 ;
        RECT 30.800 219.195 31.420 219.380 ;
        RECT 62.400 219.195 63.020 219.380 ;
        RECT 30.800 218.965 63.020 219.195 ;
        RECT 30.800 218.780 31.420 218.965 ;
        RECT 62.400 218.780 63.020 218.965 ;
        RECT 63.250 219.195 63.870 219.380 ;
        RECT 94.850 219.195 95.470 219.380 ;
        RECT 63.250 218.965 95.470 219.195 ;
        RECT 63.250 218.780 63.870 218.965 ;
        RECT 94.850 218.780 95.470 218.965 ;
        RECT 50.720 218.700 52.340 218.710 ;
        RECT 83.170 218.700 84.790 218.710 ;
        RECT 31.650 218.330 62.170 218.700 ;
        RECT 64.100 218.330 94.620 218.700 ;
        RECT 31.650 217.610 62.170 217.990 ;
        RECT 64.100 217.610 94.620 217.990 ;
        RECT 30.800 217.355 31.420 217.540 ;
        RECT 62.400 217.355 63.020 217.540 ;
        RECT 30.800 217.125 63.020 217.355 ;
        RECT 30.800 216.940 31.420 217.125 ;
        RECT 62.400 216.940 63.020 217.125 ;
        RECT 63.250 217.355 63.870 217.540 ;
        RECT 94.850 217.355 95.470 217.540 ;
        RECT 63.250 217.125 95.470 217.355 ;
        RECT 63.250 216.940 63.870 217.125 ;
        RECT 94.850 216.940 95.470 217.125 ;
        RECT 46.880 216.860 48.500 216.870 ;
        RECT 79.330 216.860 80.950 216.870 ;
        RECT 31.650 216.490 62.170 216.860 ;
        RECT 64.100 216.490 94.620 216.860 ;
        RECT 31.650 215.770 62.170 216.150 ;
        RECT 64.100 215.770 94.620 216.150 ;
        RECT 30.800 215.515 31.420 215.700 ;
        RECT 62.400 215.515 63.020 215.700 ;
        RECT 30.800 215.285 63.020 215.515 ;
        RECT 30.800 215.100 31.420 215.285 ;
        RECT 62.400 215.100 63.020 215.285 ;
        RECT 63.250 215.515 63.870 215.700 ;
        RECT 94.850 215.515 95.470 215.700 ;
        RECT 63.250 215.285 95.470 215.515 ;
        RECT 63.250 215.100 63.870 215.285 ;
        RECT 94.850 215.100 95.470 215.285 ;
        RECT 43.040 215.020 44.660 215.030 ;
        RECT 75.490 215.020 77.110 215.030 ;
        RECT 31.650 214.650 62.170 215.020 ;
        RECT 64.100 214.650 94.620 215.020 ;
        RECT 31.660 213.855 62.160 214.295 ;
        RECT 64.110 213.855 94.610 214.295 ;
        RECT 31.650 213.125 62.170 213.505 ;
        RECT 64.100 213.125 94.620 213.505 ;
        RECT 30.800 212.870 31.420 213.055 ;
        RECT 62.400 212.870 63.020 213.055 ;
        RECT 30.800 212.640 63.020 212.870 ;
        RECT 30.800 212.455 31.420 212.640 ;
        RECT 62.400 212.455 63.020 212.640 ;
        RECT 63.250 212.870 63.870 213.055 ;
        RECT 94.850 212.870 95.470 213.055 ;
        RECT 63.250 212.640 95.470 212.870 ;
        RECT 63.250 212.455 63.870 212.640 ;
        RECT 94.850 212.455 95.470 212.640 ;
        RECT 39.200 212.375 40.820 212.385 ;
        RECT 71.650 212.375 73.270 212.385 ;
        RECT 31.650 212.005 62.170 212.375 ;
        RECT 64.100 212.005 94.620 212.375 ;
        RECT 31.650 211.285 62.170 211.665 ;
        RECT 64.100 211.285 94.620 211.665 ;
        RECT 30.800 211.030 31.420 211.215 ;
        RECT 62.400 211.030 63.020 211.215 ;
        RECT 30.800 210.800 63.020 211.030 ;
        RECT 30.800 210.615 31.420 210.800 ;
        RECT 62.400 210.615 63.020 210.800 ;
        RECT 63.250 211.030 63.870 211.215 ;
        RECT 94.850 211.030 95.470 211.215 ;
        RECT 63.250 210.800 95.470 211.030 ;
        RECT 63.250 210.615 63.870 210.800 ;
        RECT 94.850 210.615 95.470 210.800 ;
        RECT 35.360 210.535 36.980 210.545 ;
        RECT 67.810 210.535 69.430 210.545 ;
        RECT 31.650 210.165 62.170 210.535 ;
        RECT 64.100 210.165 94.620 210.535 ;
        RECT 31.650 209.445 62.170 209.825 ;
        RECT 64.100 209.445 94.620 209.825 ;
        RECT 30.800 209.190 31.420 209.375 ;
        RECT 62.400 209.190 63.020 209.375 ;
        RECT 30.800 208.960 63.020 209.190 ;
        RECT 30.800 208.775 31.420 208.960 ;
        RECT 62.400 208.775 63.020 208.960 ;
        RECT 63.250 209.190 63.870 209.375 ;
        RECT 94.850 209.190 95.470 209.375 ;
        RECT 63.250 208.960 95.470 209.190 ;
        RECT 63.250 208.775 63.870 208.960 ;
        RECT 94.850 208.775 95.470 208.960 ;
        RECT 31.650 208.325 62.170 208.695 ;
        RECT 64.100 208.325 94.620 208.695 ;
        RECT 25.090 205.975 27.380 206.315 ;
        RECT 28.125 205.975 29.610 206.315 ;
        RECT 25.090 205.340 25.690 205.975 ;
        RECT 25.090 205.110 26.670 205.340 ;
        RECT 25.090 203.070 25.690 205.110 ;
        RECT 27.100 204.880 27.460 204.965 ;
        RECT 25.970 204.650 27.460 204.880 ;
        RECT 25.970 204.500 26.330 204.650 ;
        RECT 25.920 203.865 26.870 204.270 ;
        RECT 25.090 202.840 26.380 203.070 ;
        RECT 25.090 201.880 25.690 202.840 ;
        RECT 26.610 202.520 26.870 203.865 ;
        RECT 27.100 203.215 27.460 204.650 ;
        RECT 27.690 203.315 28.040 204.515 ;
        RECT 28.400 203.905 28.780 205.550 ;
        RECT 27.480 202.520 27.830 202.580 ;
        RECT 28.400 202.520 28.740 203.125 ;
        RECT 26.610 202.260 28.740 202.520 ;
        RECT 27.480 202.200 27.830 202.260 ;
        RECT 29.010 201.980 29.610 205.975 ;
        RECT 31.455 205.540 33.205 208.325 ;
        RECT 33.845 205.540 34.655 206.540 ;
        RECT 35.295 205.540 37.045 207.835 ;
        RECT 37.685 205.540 38.495 206.540 ;
        RECT 39.135 205.540 40.885 207.835 ;
        RECT 41.525 205.540 42.335 206.540 ;
        RECT 42.975 205.540 44.725 207.835 ;
        RECT 45.365 205.540 46.175 206.540 ;
        RECT 46.815 205.540 48.565 207.835 ;
        RECT 49.205 205.540 50.015 206.540 ;
        RECT 50.655 205.540 52.405 207.835 ;
        RECT 53.045 205.540 53.855 206.540 ;
        RECT 54.495 205.540 56.245 207.835 ;
        RECT 56.885 205.540 57.695 206.540 ;
        RECT 58.335 205.540 60.085 207.835 ;
        RECT 60.725 205.540 61.535 206.540 ;
        RECT 63.905 205.540 65.655 208.325 ;
        RECT 66.295 205.540 67.105 206.540 ;
        RECT 67.745 205.540 69.495 207.835 ;
        RECT 70.135 205.540 70.945 206.540 ;
        RECT 71.585 205.540 73.335 207.835 ;
        RECT 73.975 205.540 74.785 206.540 ;
        RECT 75.425 205.540 77.175 207.835 ;
        RECT 77.815 205.540 78.625 206.540 ;
        RECT 79.265 205.540 81.015 207.835 ;
        RECT 81.655 205.540 82.465 206.540 ;
        RECT 83.105 205.540 84.855 207.835 ;
        RECT 85.495 205.540 86.305 206.540 ;
        RECT 86.945 205.540 88.695 207.835 ;
        RECT 89.335 205.540 90.145 206.540 ;
        RECT 90.785 205.540 92.535 207.835 ;
        RECT 93.175 205.540 93.985 206.540 ;
        RECT 96.400 205.730 96.770 224.240 ;
        RECT 97.420 220.605 97.790 224.240 ;
        RECT 97.415 220.225 97.795 220.605 ;
        RECT 97.420 217.605 97.790 220.225 ;
        RECT 97.415 217.225 97.795 217.605 ;
        RECT 97.420 214.605 97.790 217.225 ;
        RECT 97.415 214.225 97.795 214.605 ;
        RECT 97.420 211.605 97.790 214.225 ;
        RECT 97.415 211.225 97.795 211.605 ;
        RECT 97.420 208.605 97.790 211.225 ;
        RECT 97.415 208.225 97.795 208.605 ;
        RECT 96.400 205.350 96.780 205.730 ;
        RECT 96.400 204.280 96.770 205.350 ;
        RECT 31.925 203.090 32.735 204.090 ;
        RECT 25.090 201.650 26.780 201.880 ;
        RECT 28.150 201.750 29.610 201.980 ;
        RECT 25.090 199.640 25.690 201.650 ;
        RECT 27.110 201.190 28.110 201.515 ;
        RECT 25.920 200.630 28.780 200.960 ;
        RECT 25.090 199.410 26.780 199.640 ;
        RECT 25.090 197.400 25.690 199.410 ;
        RECT 27.495 199.275 27.760 200.630 ;
        RECT 29.010 199.740 29.610 201.750 ;
        RECT 33.375 201.260 35.125 204.090 ;
        RECT 35.765 203.090 36.575 204.090 ;
        RECT 37.215 201.795 38.965 204.090 ;
        RECT 39.605 203.090 40.415 204.090 ;
        RECT 41.055 201.795 42.805 204.090 ;
        RECT 43.445 203.090 44.255 204.090 ;
        RECT 44.895 201.795 46.645 204.090 ;
        RECT 47.285 203.090 48.095 204.090 ;
        RECT 48.735 201.795 50.485 204.090 ;
        RECT 51.125 203.090 51.935 204.090 ;
        RECT 52.575 201.795 54.325 204.090 ;
        RECT 54.965 203.090 55.775 204.090 ;
        RECT 56.415 201.795 58.165 204.090 ;
        RECT 58.805 203.090 59.615 204.090 ;
        RECT 60.255 201.795 62.005 204.090 ;
        RECT 64.375 203.090 65.185 204.090 ;
        RECT 65.825 201.260 67.575 204.090 ;
        RECT 68.215 203.090 69.025 204.090 ;
        RECT 69.665 201.795 71.415 204.090 ;
        RECT 72.055 203.090 72.865 204.090 ;
        RECT 73.505 201.795 75.255 204.090 ;
        RECT 75.895 203.090 76.705 204.090 ;
        RECT 77.345 201.795 79.095 204.090 ;
        RECT 79.735 203.090 80.545 204.090 ;
        RECT 81.185 201.795 82.935 204.090 ;
        RECT 83.575 203.090 84.385 204.090 ;
        RECT 85.025 201.795 86.775 204.090 ;
        RECT 87.415 203.090 88.225 204.090 ;
        RECT 88.865 201.795 90.615 204.090 ;
        RECT 91.255 203.090 92.065 204.090 ;
        RECT 92.705 201.795 94.455 204.090 ;
        RECT 96.400 203.900 96.780 204.280 ;
        RECT 31.650 200.890 62.170 201.260 ;
        RECT 64.100 200.890 94.620 201.260 ;
        RECT 30.800 200.625 31.420 200.810 ;
        RECT 62.400 200.625 63.020 200.810 ;
        RECT 30.800 200.395 63.020 200.625 ;
        RECT 30.800 200.210 31.420 200.395 ;
        RECT 62.400 200.210 63.020 200.395 ;
        RECT 63.250 200.625 63.870 200.810 ;
        RECT 94.850 200.625 95.470 200.810 ;
        RECT 63.250 200.395 95.470 200.625 ;
        RECT 63.250 200.210 63.870 200.395 ;
        RECT 94.850 200.210 95.470 200.395 ;
        RECT 31.650 199.760 62.170 200.140 ;
        RECT 64.100 199.760 94.620 200.140 ;
        RECT 28.150 199.510 29.610 199.740 ;
        RECT 27.110 198.950 28.110 199.275 ;
        RECT 25.920 198.390 28.780 198.720 ;
        RECT 29.010 197.500 29.610 199.510 ;
        RECT 31.650 199.050 62.170 199.420 ;
        RECT 64.100 199.050 94.620 199.420 ;
        RECT 37.280 199.040 38.900 199.050 ;
        RECT 69.730 199.040 71.350 199.050 ;
        RECT 30.800 198.785 31.420 198.970 ;
        RECT 62.400 198.785 63.020 198.970 ;
        RECT 30.800 198.555 63.020 198.785 ;
        RECT 30.800 198.370 31.420 198.555 ;
        RECT 62.400 198.370 63.020 198.555 ;
        RECT 63.250 198.785 63.870 198.970 ;
        RECT 94.850 198.785 95.470 198.970 ;
        RECT 63.250 198.555 95.470 198.785 ;
        RECT 63.250 198.370 63.870 198.555 ;
        RECT 94.850 198.370 95.470 198.555 ;
        RECT 31.650 197.920 62.170 198.300 ;
        RECT 64.100 197.920 94.620 198.300 ;
        RECT 25.090 197.170 26.780 197.400 ;
        RECT 28.150 197.270 29.610 197.500 ;
        RECT 25.090 195.115 25.690 197.170 ;
        RECT 27.110 196.710 28.110 197.035 ;
        RECT 29.010 195.115 29.610 197.270 ;
        RECT 31.650 197.205 62.170 197.575 ;
        RECT 64.100 197.205 94.620 197.575 ;
        RECT 41.120 197.195 42.740 197.205 ;
        RECT 73.570 197.195 75.190 197.205 ;
        RECT 30.800 196.940 31.420 197.125 ;
        RECT 62.400 196.940 63.020 197.125 ;
        RECT 30.800 196.710 63.020 196.940 ;
        RECT 30.800 196.525 31.420 196.710 ;
        RECT 62.400 196.525 63.020 196.710 ;
        RECT 63.250 196.940 63.870 197.125 ;
        RECT 94.850 196.940 95.470 197.125 ;
        RECT 63.250 196.710 95.470 196.940 ;
        RECT 63.250 196.525 63.870 196.710 ;
        RECT 94.850 196.525 95.470 196.710 ;
        RECT 31.650 196.075 62.170 196.455 ;
        RECT 64.100 196.075 94.620 196.455 ;
        RECT 31.660 195.285 62.160 195.725 ;
        RECT 64.110 195.285 94.610 195.725 ;
        RECT 25.090 194.775 27.380 195.115 ;
        RECT 28.125 194.775 29.610 195.115 ;
        RECT 25.090 166.930 25.690 194.775 ;
        RECT 29.010 166.930 29.610 194.775 ;
        RECT 31.650 194.565 62.170 194.935 ;
        RECT 64.100 194.565 94.620 194.935 ;
        RECT 44.960 194.555 46.580 194.565 ;
        RECT 77.410 194.555 79.030 194.565 ;
        RECT 30.800 194.300 31.420 194.485 ;
        RECT 62.400 194.300 63.020 194.485 ;
        RECT 30.800 194.070 63.020 194.300 ;
        RECT 30.800 193.885 31.420 194.070 ;
        RECT 62.400 193.885 63.020 194.070 ;
        RECT 63.250 194.300 63.870 194.485 ;
        RECT 94.850 194.300 95.470 194.485 ;
        RECT 63.250 194.070 95.470 194.300 ;
        RECT 63.250 193.885 63.870 194.070 ;
        RECT 94.850 193.885 95.470 194.070 ;
        RECT 31.650 193.435 62.170 193.815 ;
        RECT 64.100 193.435 94.620 193.815 ;
        RECT 31.650 192.725 62.170 193.095 ;
        RECT 64.100 192.725 94.620 193.095 ;
        RECT 48.800 192.715 50.420 192.725 ;
        RECT 81.250 192.715 82.870 192.725 ;
        RECT 30.800 192.460 31.420 192.645 ;
        RECT 62.400 192.460 63.020 192.645 ;
        RECT 30.800 192.230 63.020 192.460 ;
        RECT 30.800 192.045 31.420 192.230 ;
        RECT 62.400 192.045 63.020 192.230 ;
        RECT 63.250 192.460 63.870 192.645 ;
        RECT 94.850 192.460 95.470 192.645 ;
        RECT 63.250 192.230 95.470 192.460 ;
        RECT 63.250 192.045 63.870 192.230 ;
        RECT 94.850 192.045 95.470 192.230 ;
        RECT 31.650 191.595 62.170 191.975 ;
        RECT 64.100 191.595 94.620 191.975 ;
        RECT 31.650 190.880 62.170 191.250 ;
        RECT 64.100 190.880 94.620 191.250 ;
        RECT 52.640 190.870 54.260 190.880 ;
        RECT 85.090 190.870 86.710 190.880 ;
        RECT 30.800 190.615 31.420 190.800 ;
        RECT 62.400 190.615 63.020 190.800 ;
        RECT 30.800 190.385 63.020 190.615 ;
        RECT 30.800 190.200 31.420 190.385 ;
        RECT 62.400 190.200 63.020 190.385 ;
        RECT 63.250 190.615 63.870 190.800 ;
        RECT 94.850 190.615 95.470 190.800 ;
        RECT 63.250 190.385 95.470 190.615 ;
        RECT 63.250 190.200 63.870 190.385 ;
        RECT 94.850 190.200 95.470 190.385 ;
        RECT 31.650 189.750 62.170 190.130 ;
        RECT 64.100 189.750 94.620 190.130 ;
        RECT 31.660 188.960 62.160 189.400 ;
        RECT 64.110 188.960 94.610 189.400 ;
        RECT 31.650 188.240 62.170 188.610 ;
        RECT 64.100 188.240 94.620 188.610 ;
        RECT 56.480 188.230 58.100 188.240 ;
        RECT 88.930 188.230 90.550 188.240 ;
        RECT 30.800 187.975 31.420 188.160 ;
        RECT 62.400 187.975 63.020 188.160 ;
        RECT 30.800 187.745 63.020 187.975 ;
        RECT 30.800 187.560 31.420 187.745 ;
        RECT 62.400 187.560 63.020 187.745 ;
        RECT 63.250 187.975 63.870 188.160 ;
        RECT 94.850 187.975 95.470 188.160 ;
        RECT 63.250 187.745 95.470 187.975 ;
        RECT 63.250 187.560 63.870 187.745 ;
        RECT 94.850 187.560 95.470 187.745 ;
        RECT 31.650 187.110 62.170 187.490 ;
        RECT 64.100 187.110 94.620 187.490 ;
        RECT 31.650 186.400 62.170 186.770 ;
        RECT 64.100 186.400 94.620 186.770 ;
        RECT 60.320 186.390 61.940 186.400 ;
        RECT 92.770 186.390 94.390 186.400 ;
        RECT 30.800 186.135 31.420 186.320 ;
        RECT 62.400 186.135 63.020 186.320 ;
        RECT 30.800 185.905 63.020 186.135 ;
        RECT 30.800 185.720 31.420 185.905 ;
        RECT 62.400 185.720 63.020 185.905 ;
        RECT 63.250 186.135 63.870 186.320 ;
        RECT 94.850 186.135 95.470 186.320 ;
        RECT 63.250 185.905 95.470 186.135 ;
        RECT 96.400 185.970 96.770 203.900 ;
        RECT 97.420 202.605 97.790 208.225 ;
        RECT 98.440 205.730 98.810 224.240 ;
        RECT 99.460 220.605 99.830 224.240 ;
        RECT 99.455 220.225 99.835 220.605 ;
        RECT 99.460 217.605 99.830 220.225 ;
        RECT 99.455 217.225 99.835 217.605 ;
        RECT 99.460 214.605 99.830 217.225 ;
        RECT 99.455 214.225 99.835 214.605 ;
        RECT 99.460 211.605 99.830 214.225 ;
        RECT 99.455 211.225 99.835 211.605 ;
        RECT 99.460 208.605 99.830 211.225 ;
        RECT 99.455 208.225 99.835 208.605 ;
        RECT 98.440 205.350 98.820 205.730 ;
        RECT 98.440 204.280 98.810 205.350 ;
        RECT 98.440 203.900 98.820 204.280 ;
        RECT 97.415 202.225 97.795 202.605 ;
        RECT 97.420 199.605 97.790 202.225 ;
        RECT 97.415 199.225 97.795 199.605 ;
        RECT 97.420 196.605 97.790 199.225 ;
        RECT 97.415 196.225 97.795 196.605 ;
        RECT 97.420 193.605 97.790 196.225 ;
        RECT 97.415 193.225 97.795 193.605 ;
        RECT 97.420 190.605 97.790 193.225 ;
        RECT 97.415 190.225 97.795 190.605 ;
        RECT 97.420 187.605 97.790 190.225 ;
        RECT 97.415 187.225 97.795 187.605 ;
        RECT 97.420 185.970 97.790 187.225 ;
        RECT 98.440 185.970 98.810 203.900 ;
        RECT 99.460 202.605 99.830 208.225 ;
        RECT 99.455 202.225 99.835 202.605 ;
        RECT 99.460 199.605 99.830 202.225 ;
        RECT 99.455 199.225 99.835 199.605 ;
        RECT 99.460 196.605 99.830 199.225 ;
        RECT 99.455 196.225 99.835 196.605 ;
        RECT 99.460 193.605 99.830 196.225 ;
        RECT 99.455 193.225 99.835 193.605 ;
        RECT 99.460 190.605 99.830 193.225 ;
        RECT 99.455 190.225 99.835 190.605 ;
        RECT 99.460 187.605 99.830 190.225 ;
        RECT 99.455 187.225 99.835 187.605 ;
        RECT 99.460 185.970 99.830 187.225 ;
        RECT 100.480 185.970 100.860 224.240 ;
        RECT 101.210 185.980 101.650 224.230 ;
        RECT 63.250 185.720 63.870 185.905 ;
        RECT 94.850 185.720 95.470 185.905 ;
        RECT 31.650 185.270 62.170 185.650 ;
        RECT 64.100 185.270 94.620 185.650 ;
        RECT 31.650 184.550 62.170 184.930 ;
        RECT 64.100 184.550 94.620 184.930 ;
        RECT 30.800 184.295 31.420 184.480 ;
        RECT 62.400 184.295 63.020 184.480 ;
        RECT 30.800 184.065 63.020 184.295 ;
        RECT 30.800 183.880 31.420 184.065 ;
        RECT 62.400 183.880 63.020 184.065 ;
        RECT 63.250 184.295 63.870 184.480 ;
        RECT 94.850 184.295 95.470 184.480 ;
        RECT 63.250 184.065 95.470 184.295 ;
        RECT 63.250 183.880 63.870 184.065 ;
        RECT 94.850 183.880 95.470 184.065 ;
        RECT 58.400 183.800 60.020 183.810 ;
        RECT 90.850 183.800 92.470 183.810 ;
        RECT 31.650 183.430 62.170 183.800 ;
        RECT 64.100 183.430 94.620 183.800 ;
        RECT 31.650 182.710 62.170 183.090 ;
        RECT 64.100 182.710 94.620 183.090 ;
        RECT 30.800 182.455 31.420 182.640 ;
        RECT 62.400 182.455 63.020 182.640 ;
        RECT 30.800 182.225 63.020 182.455 ;
        RECT 30.800 182.040 31.420 182.225 ;
        RECT 62.400 182.040 63.020 182.225 ;
        RECT 63.250 182.455 63.870 182.640 ;
        RECT 94.850 182.455 95.470 182.640 ;
        RECT 63.250 182.225 95.470 182.455 ;
        RECT 63.250 182.040 63.870 182.225 ;
        RECT 94.850 182.040 95.470 182.225 ;
        RECT 54.560 181.960 56.180 181.970 ;
        RECT 87.010 181.960 88.630 181.970 ;
        RECT 31.650 181.590 62.170 181.960 ;
        RECT 64.100 181.590 94.620 181.960 ;
        RECT 31.660 180.795 62.160 181.235 ;
        RECT 64.110 180.795 94.610 181.235 ;
        RECT 31.650 180.065 62.170 180.445 ;
        RECT 64.100 180.065 94.620 180.445 ;
        RECT 30.800 179.810 31.420 179.995 ;
        RECT 62.400 179.810 63.020 179.995 ;
        RECT 30.800 179.580 63.020 179.810 ;
        RECT 30.800 179.395 31.420 179.580 ;
        RECT 62.400 179.395 63.020 179.580 ;
        RECT 63.250 179.810 63.870 179.995 ;
        RECT 94.850 179.810 95.470 179.995 ;
        RECT 63.250 179.580 95.470 179.810 ;
        RECT 63.250 179.395 63.870 179.580 ;
        RECT 94.850 179.395 95.470 179.580 ;
        RECT 50.720 179.315 52.340 179.325 ;
        RECT 83.170 179.315 84.790 179.325 ;
        RECT 31.650 178.945 62.170 179.315 ;
        RECT 64.100 178.945 94.620 179.315 ;
        RECT 31.650 178.225 62.170 178.605 ;
        RECT 64.100 178.225 94.620 178.605 ;
        RECT 30.800 177.970 31.420 178.155 ;
        RECT 62.400 177.970 63.020 178.155 ;
        RECT 30.800 177.740 63.020 177.970 ;
        RECT 30.800 177.555 31.420 177.740 ;
        RECT 62.400 177.555 63.020 177.740 ;
        RECT 63.250 177.970 63.870 178.155 ;
        RECT 94.850 177.970 95.470 178.155 ;
        RECT 63.250 177.740 95.470 177.970 ;
        RECT 63.250 177.555 63.870 177.740 ;
        RECT 94.850 177.555 95.470 177.740 ;
        RECT 46.880 177.475 48.500 177.485 ;
        RECT 79.330 177.475 80.950 177.485 ;
        RECT 31.650 177.105 62.170 177.475 ;
        RECT 64.100 177.105 94.620 177.475 ;
        RECT 31.650 176.385 62.170 176.765 ;
        RECT 64.100 176.385 94.620 176.765 ;
        RECT 30.800 176.130 31.420 176.315 ;
        RECT 62.400 176.130 63.020 176.315 ;
        RECT 30.800 175.900 63.020 176.130 ;
        RECT 30.800 175.715 31.420 175.900 ;
        RECT 62.400 175.715 63.020 175.900 ;
        RECT 63.250 176.130 63.870 176.315 ;
        RECT 94.850 176.130 95.470 176.315 ;
        RECT 63.250 175.900 95.470 176.130 ;
        RECT 63.250 175.715 63.870 175.900 ;
        RECT 94.850 175.715 95.470 175.900 ;
        RECT 43.040 175.635 44.660 175.645 ;
        RECT 75.490 175.635 77.110 175.645 ;
        RECT 31.650 175.265 62.170 175.635 ;
        RECT 64.100 175.265 94.620 175.635 ;
        RECT 31.660 174.470 62.160 174.910 ;
        RECT 64.110 174.470 94.610 174.910 ;
        RECT 31.650 173.740 62.170 174.120 ;
        RECT 64.100 173.740 94.620 174.120 ;
        RECT 30.800 173.485 31.420 173.670 ;
        RECT 62.400 173.485 63.020 173.670 ;
        RECT 30.800 173.255 63.020 173.485 ;
        RECT 30.800 173.070 31.420 173.255 ;
        RECT 62.400 173.070 63.020 173.255 ;
        RECT 63.250 173.485 63.870 173.670 ;
        RECT 94.850 173.485 95.470 173.670 ;
        RECT 63.250 173.255 95.470 173.485 ;
        RECT 63.250 173.070 63.870 173.255 ;
        RECT 94.850 173.070 95.470 173.255 ;
        RECT 39.200 172.990 40.820 173.000 ;
        RECT 71.650 172.990 73.270 173.000 ;
        RECT 31.650 172.620 62.170 172.990 ;
        RECT 64.100 172.620 94.620 172.990 ;
        RECT 31.650 171.900 62.170 172.280 ;
        RECT 64.100 171.900 94.620 172.280 ;
        RECT 30.800 171.645 31.420 171.830 ;
        RECT 62.400 171.645 63.020 171.830 ;
        RECT 30.800 171.415 63.020 171.645 ;
        RECT 30.800 171.230 31.420 171.415 ;
        RECT 62.400 171.230 63.020 171.415 ;
        RECT 63.250 171.645 63.870 171.830 ;
        RECT 94.850 171.645 95.470 171.830 ;
        RECT 63.250 171.415 95.470 171.645 ;
        RECT 63.250 171.230 63.870 171.415 ;
        RECT 94.850 171.230 95.470 171.415 ;
        RECT 35.360 171.150 36.980 171.160 ;
        RECT 67.810 171.150 69.430 171.160 ;
        RECT 31.650 170.780 62.170 171.150 ;
        RECT 64.100 170.780 94.620 171.150 ;
        RECT 31.650 170.060 62.170 170.440 ;
        RECT 64.100 170.060 94.620 170.440 ;
        RECT 30.800 169.805 31.420 169.990 ;
        RECT 62.400 169.805 63.020 169.990 ;
        RECT 30.800 169.575 63.020 169.805 ;
        RECT 30.800 169.390 31.420 169.575 ;
        RECT 62.400 169.390 63.020 169.575 ;
        RECT 63.250 169.805 63.870 169.990 ;
        RECT 94.850 169.805 95.470 169.990 ;
        RECT 63.250 169.575 95.470 169.805 ;
        RECT 63.250 169.390 63.870 169.575 ;
        RECT 94.850 169.390 95.470 169.575 ;
        RECT 31.650 168.940 62.170 169.310 ;
        RECT 64.100 168.940 94.620 169.310 ;
        RECT 25.090 166.590 27.380 166.930 ;
        RECT 28.125 166.590 29.610 166.930 ;
        RECT 25.090 165.955 25.690 166.590 ;
        RECT 25.090 165.725 26.670 165.955 ;
        RECT 25.090 163.685 25.690 165.725 ;
        RECT 27.100 165.495 27.460 165.580 ;
        RECT 25.970 165.265 27.460 165.495 ;
        RECT 25.970 165.115 26.330 165.265 ;
        RECT 25.920 164.480 26.870 164.885 ;
        RECT 25.090 163.455 26.380 163.685 ;
        RECT 25.090 162.495 25.690 163.455 ;
        RECT 26.610 163.135 26.870 164.480 ;
        RECT 27.100 163.830 27.460 165.265 ;
        RECT 27.690 163.930 28.040 165.130 ;
        RECT 28.400 164.520 28.780 166.165 ;
        RECT 27.480 163.135 27.830 163.195 ;
        RECT 28.400 163.135 28.740 163.740 ;
        RECT 26.610 162.875 28.740 163.135 ;
        RECT 27.480 162.815 27.830 162.875 ;
        RECT 29.010 162.595 29.610 166.590 ;
        RECT 31.455 166.155 33.205 168.940 ;
        RECT 33.845 166.155 34.655 167.155 ;
        RECT 35.295 166.155 37.045 168.450 ;
        RECT 37.685 166.155 38.495 167.155 ;
        RECT 39.135 166.155 40.885 168.450 ;
        RECT 41.525 166.155 42.335 167.155 ;
        RECT 42.975 166.155 44.725 168.450 ;
        RECT 45.365 166.155 46.175 167.155 ;
        RECT 46.815 166.155 48.565 168.450 ;
        RECT 49.205 166.155 50.015 167.155 ;
        RECT 50.655 166.155 52.405 168.450 ;
        RECT 53.045 166.155 53.855 167.155 ;
        RECT 54.495 166.155 56.245 168.450 ;
        RECT 56.885 166.155 57.695 167.155 ;
        RECT 58.335 166.155 60.085 168.450 ;
        RECT 60.725 166.155 61.535 167.155 ;
        RECT 63.905 166.155 65.655 168.940 ;
        RECT 66.295 166.155 67.105 167.155 ;
        RECT 67.745 166.155 69.495 168.450 ;
        RECT 70.135 166.155 70.945 167.155 ;
        RECT 71.585 166.155 73.335 168.450 ;
        RECT 73.975 166.155 74.785 167.155 ;
        RECT 75.425 166.155 77.175 168.450 ;
        RECT 77.815 166.155 78.625 167.155 ;
        RECT 79.265 166.155 81.015 168.450 ;
        RECT 81.655 166.155 82.465 167.155 ;
        RECT 83.105 166.155 84.855 168.450 ;
        RECT 85.495 166.155 86.305 167.155 ;
        RECT 86.945 166.155 88.695 168.450 ;
        RECT 89.335 166.155 90.145 167.155 ;
        RECT 90.785 166.155 92.535 168.450 ;
        RECT 93.175 166.155 93.985 167.155 ;
        RECT 96.400 166.345 96.770 184.855 ;
        RECT 97.420 181.220 97.790 184.855 ;
        RECT 97.415 180.840 97.795 181.220 ;
        RECT 97.420 178.220 97.790 180.840 ;
        RECT 97.415 177.840 97.795 178.220 ;
        RECT 97.420 175.220 97.790 177.840 ;
        RECT 97.415 174.840 97.795 175.220 ;
        RECT 97.420 172.220 97.790 174.840 ;
        RECT 97.415 171.840 97.795 172.220 ;
        RECT 97.420 169.220 97.790 171.840 ;
        RECT 97.415 168.840 97.795 169.220 ;
        RECT 96.400 165.965 96.780 166.345 ;
        RECT 96.400 164.895 96.770 165.965 ;
        RECT 31.925 163.705 32.735 164.705 ;
        RECT 25.090 162.265 26.780 162.495 ;
        RECT 28.150 162.365 29.610 162.595 ;
        RECT 25.090 160.255 25.690 162.265 ;
        RECT 27.110 161.805 28.110 162.130 ;
        RECT 25.920 161.245 28.780 161.575 ;
        RECT 25.090 160.025 26.780 160.255 ;
        RECT 25.090 158.015 25.690 160.025 ;
        RECT 27.495 159.890 27.760 161.245 ;
        RECT 29.010 160.355 29.610 162.365 ;
        RECT 33.375 161.875 35.125 164.705 ;
        RECT 35.765 163.705 36.575 164.705 ;
        RECT 37.215 162.410 38.965 164.705 ;
        RECT 39.605 163.705 40.415 164.705 ;
        RECT 41.055 162.410 42.805 164.705 ;
        RECT 43.445 163.705 44.255 164.705 ;
        RECT 44.895 162.410 46.645 164.705 ;
        RECT 47.285 163.705 48.095 164.705 ;
        RECT 48.735 162.410 50.485 164.705 ;
        RECT 51.125 163.705 51.935 164.705 ;
        RECT 52.575 162.410 54.325 164.705 ;
        RECT 54.965 163.705 55.775 164.705 ;
        RECT 56.415 162.410 58.165 164.705 ;
        RECT 58.805 163.705 59.615 164.705 ;
        RECT 60.255 162.410 62.005 164.705 ;
        RECT 64.375 163.705 65.185 164.705 ;
        RECT 65.825 161.875 67.575 164.705 ;
        RECT 68.215 163.705 69.025 164.705 ;
        RECT 69.665 162.410 71.415 164.705 ;
        RECT 72.055 163.705 72.865 164.705 ;
        RECT 73.505 162.410 75.255 164.705 ;
        RECT 75.895 163.705 76.705 164.705 ;
        RECT 77.345 162.410 79.095 164.705 ;
        RECT 79.735 163.705 80.545 164.705 ;
        RECT 81.185 162.410 82.935 164.705 ;
        RECT 83.575 163.705 84.385 164.705 ;
        RECT 85.025 162.410 86.775 164.705 ;
        RECT 87.415 163.705 88.225 164.705 ;
        RECT 88.865 162.410 90.615 164.705 ;
        RECT 91.255 163.705 92.065 164.705 ;
        RECT 92.705 162.410 94.455 164.705 ;
        RECT 96.400 164.515 96.780 164.895 ;
        RECT 31.650 161.505 62.170 161.875 ;
        RECT 64.100 161.505 94.620 161.875 ;
        RECT 30.800 161.240 31.420 161.425 ;
        RECT 62.400 161.240 63.020 161.425 ;
        RECT 30.800 161.010 63.020 161.240 ;
        RECT 30.800 160.825 31.420 161.010 ;
        RECT 62.400 160.825 63.020 161.010 ;
        RECT 63.250 161.240 63.870 161.425 ;
        RECT 94.850 161.240 95.470 161.425 ;
        RECT 63.250 161.010 95.470 161.240 ;
        RECT 63.250 160.825 63.870 161.010 ;
        RECT 94.850 160.825 95.470 161.010 ;
        RECT 31.650 160.375 62.170 160.755 ;
        RECT 64.100 160.375 94.620 160.755 ;
        RECT 28.150 160.125 29.610 160.355 ;
        RECT 27.110 159.565 28.110 159.890 ;
        RECT 25.920 159.005 28.780 159.335 ;
        RECT 29.010 158.115 29.610 160.125 ;
        RECT 31.650 159.665 62.170 160.035 ;
        RECT 64.100 159.665 94.620 160.035 ;
        RECT 37.280 159.655 38.900 159.665 ;
        RECT 69.730 159.655 71.350 159.665 ;
        RECT 30.800 159.400 31.420 159.585 ;
        RECT 62.400 159.400 63.020 159.585 ;
        RECT 30.800 159.170 63.020 159.400 ;
        RECT 30.800 158.985 31.420 159.170 ;
        RECT 62.400 158.985 63.020 159.170 ;
        RECT 63.250 159.400 63.870 159.585 ;
        RECT 94.850 159.400 95.470 159.585 ;
        RECT 63.250 159.170 95.470 159.400 ;
        RECT 63.250 158.985 63.870 159.170 ;
        RECT 94.850 158.985 95.470 159.170 ;
        RECT 31.650 158.535 62.170 158.915 ;
        RECT 64.100 158.535 94.620 158.915 ;
        RECT 25.090 157.785 26.780 158.015 ;
        RECT 28.150 157.885 29.610 158.115 ;
        RECT 25.090 155.730 25.690 157.785 ;
        RECT 27.110 157.325 28.110 157.650 ;
        RECT 29.010 155.730 29.610 157.885 ;
        RECT 31.650 157.820 62.170 158.190 ;
        RECT 64.100 157.820 94.620 158.190 ;
        RECT 41.120 157.810 42.740 157.820 ;
        RECT 73.570 157.810 75.190 157.820 ;
        RECT 30.800 157.555 31.420 157.740 ;
        RECT 62.400 157.555 63.020 157.740 ;
        RECT 30.800 157.325 63.020 157.555 ;
        RECT 30.800 157.140 31.420 157.325 ;
        RECT 62.400 157.140 63.020 157.325 ;
        RECT 63.250 157.555 63.870 157.740 ;
        RECT 94.850 157.555 95.470 157.740 ;
        RECT 63.250 157.325 95.470 157.555 ;
        RECT 63.250 157.140 63.870 157.325 ;
        RECT 94.850 157.140 95.470 157.325 ;
        RECT 31.650 156.690 62.170 157.070 ;
        RECT 64.100 156.690 94.620 157.070 ;
        RECT 31.660 155.900 62.160 156.340 ;
        RECT 64.110 155.900 94.610 156.340 ;
        RECT 25.090 155.390 27.380 155.730 ;
        RECT 28.125 155.390 29.610 155.730 ;
        RECT 25.090 127.545 25.690 155.390 ;
        RECT 29.010 127.545 29.610 155.390 ;
        RECT 31.650 155.180 62.170 155.550 ;
        RECT 64.100 155.180 94.620 155.550 ;
        RECT 44.960 155.170 46.580 155.180 ;
        RECT 77.410 155.170 79.030 155.180 ;
        RECT 30.800 154.915 31.420 155.100 ;
        RECT 62.400 154.915 63.020 155.100 ;
        RECT 30.800 154.685 63.020 154.915 ;
        RECT 30.800 154.500 31.420 154.685 ;
        RECT 62.400 154.500 63.020 154.685 ;
        RECT 63.250 154.915 63.870 155.100 ;
        RECT 94.850 154.915 95.470 155.100 ;
        RECT 63.250 154.685 95.470 154.915 ;
        RECT 63.250 154.500 63.870 154.685 ;
        RECT 94.850 154.500 95.470 154.685 ;
        RECT 31.650 154.050 62.170 154.430 ;
        RECT 64.100 154.050 94.620 154.430 ;
        RECT 31.650 153.340 62.170 153.710 ;
        RECT 64.100 153.340 94.620 153.710 ;
        RECT 48.800 153.330 50.420 153.340 ;
        RECT 81.250 153.330 82.870 153.340 ;
        RECT 30.800 153.075 31.420 153.260 ;
        RECT 62.400 153.075 63.020 153.260 ;
        RECT 30.800 152.845 63.020 153.075 ;
        RECT 30.800 152.660 31.420 152.845 ;
        RECT 62.400 152.660 63.020 152.845 ;
        RECT 63.250 153.075 63.870 153.260 ;
        RECT 94.850 153.075 95.470 153.260 ;
        RECT 63.250 152.845 95.470 153.075 ;
        RECT 63.250 152.660 63.870 152.845 ;
        RECT 94.850 152.660 95.470 152.845 ;
        RECT 31.650 152.210 62.170 152.590 ;
        RECT 64.100 152.210 94.620 152.590 ;
        RECT 31.650 151.495 62.170 151.865 ;
        RECT 64.100 151.495 94.620 151.865 ;
        RECT 52.640 151.485 54.260 151.495 ;
        RECT 85.090 151.485 86.710 151.495 ;
        RECT 30.800 151.230 31.420 151.415 ;
        RECT 62.400 151.230 63.020 151.415 ;
        RECT 30.800 151.000 63.020 151.230 ;
        RECT 30.800 150.815 31.420 151.000 ;
        RECT 62.400 150.815 63.020 151.000 ;
        RECT 63.250 151.230 63.870 151.415 ;
        RECT 94.850 151.230 95.470 151.415 ;
        RECT 63.250 151.000 95.470 151.230 ;
        RECT 63.250 150.815 63.870 151.000 ;
        RECT 94.850 150.815 95.470 151.000 ;
        RECT 31.650 150.365 62.170 150.745 ;
        RECT 64.100 150.365 94.620 150.745 ;
        RECT 31.660 149.575 62.160 150.015 ;
        RECT 64.110 149.575 94.610 150.015 ;
        RECT 31.650 148.855 62.170 149.225 ;
        RECT 64.100 148.855 94.620 149.225 ;
        RECT 56.480 148.845 58.100 148.855 ;
        RECT 88.930 148.845 90.550 148.855 ;
        RECT 30.800 148.590 31.420 148.775 ;
        RECT 62.400 148.590 63.020 148.775 ;
        RECT 30.800 148.360 63.020 148.590 ;
        RECT 30.800 148.175 31.420 148.360 ;
        RECT 62.400 148.175 63.020 148.360 ;
        RECT 63.250 148.590 63.870 148.775 ;
        RECT 94.850 148.590 95.470 148.775 ;
        RECT 63.250 148.360 95.470 148.590 ;
        RECT 63.250 148.175 63.870 148.360 ;
        RECT 94.850 148.175 95.470 148.360 ;
        RECT 31.650 147.725 62.170 148.105 ;
        RECT 64.100 147.725 94.620 148.105 ;
        RECT 31.650 147.015 62.170 147.385 ;
        RECT 64.100 147.015 94.620 147.385 ;
        RECT 60.320 147.005 61.940 147.015 ;
        RECT 92.770 147.005 94.390 147.015 ;
        RECT 30.800 146.750 31.420 146.935 ;
        RECT 62.400 146.750 63.020 146.935 ;
        RECT 30.800 146.520 63.020 146.750 ;
        RECT 30.800 146.335 31.420 146.520 ;
        RECT 62.400 146.335 63.020 146.520 ;
        RECT 63.250 146.750 63.870 146.935 ;
        RECT 94.850 146.750 95.470 146.935 ;
        RECT 63.250 146.520 95.470 146.750 ;
        RECT 96.400 146.585 96.770 164.515 ;
        RECT 97.420 163.220 97.790 168.840 ;
        RECT 98.440 166.345 98.810 184.855 ;
        RECT 99.460 181.220 99.830 184.855 ;
        RECT 99.455 180.840 99.835 181.220 ;
        RECT 99.460 178.220 99.830 180.840 ;
        RECT 99.455 177.840 99.835 178.220 ;
        RECT 99.460 175.220 99.830 177.840 ;
        RECT 99.455 174.840 99.835 175.220 ;
        RECT 99.460 172.220 99.830 174.840 ;
        RECT 99.455 171.840 99.835 172.220 ;
        RECT 99.460 169.220 99.830 171.840 ;
        RECT 99.455 168.840 99.835 169.220 ;
        RECT 98.440 165.965 98.820 166.345 ;
        RECT 98.440 164.895 98.810 165.965 ;
        RECT 98.440 164.515 98.820 164.895 ;
        RECT 97.415 162.840 97.795 163.220 ;
        RECT 97.420 160.220 97.790 162.840 ;
        RECT 97.415 159.840 97.795 160.220 ;
        RECT 97.420 157.220 97.790 159.840 ;
        RECT 97.415 156.840 97.795 157.220 ;
        RECT 97.420 154.220 97.790 156.840 ;
        RECT 97.415 153.840 97.795 154.220 ;
        RECT 97.420 151.220 97.790 153.840 ;
        RECT 97.415 150.840 97.795 151.220 ;
        RECT 97.420 148.220 97.790 150.840 ;
        RECT 97.415 147.840 97.795 148.220 ;
        RECT 97.420 146.585 97.790 147.840 ;
        RECT 98.440 146.585 98.810 164.515 ;
        RECT 99.460 163.220 99.830 168.840 ;
        RECT 99.455 162.840 99.835 163.220 ;
        RECT 99.460 160.220 99.830 162.840 ;
        RECT 99.455 159.840 99.835 160.220 ;
        RECT 99.460 157.220 99.830 159.840 ;
        RECT 99.455 156.840 99.835 157.220 ;
        RECT 99.460 154.220 99.830 156.840 ;
        RECT 99.455 153.840 99.835 154.220 ;
        RECT 99.460 151.220 99.830 153.840 ;
        RECT 99.455 150.840 99.835 151.220 ;
        RECT 99.460 148.220 99.830 150.840 ;
        RECT 99.455 147.840 99.835 148.220 ;
        RECT 99.460 146.585 99.830 147.840 ;
        RECT 100.480 146.585 100.860 184.855 ;
        RECT 101.210 146.595 101.650 184.845 ;
        RECT 63.250 146.335 63.870 146.520 ;
        RECT 94.850 146.335 95.470 146.520 ;
        RECT 31.650 145.885 62.170 146.265 ;
        RECT 64.100 145.885 94.620 146.265 ;
        RECT 31.650 145.165 62.170 145.545 ;
        RECT 64.100 145.165 94.620 145.545 ;
        RECT 30.800 144.910 31.420 145.095 ;
        RECT 62.400 144.910 63.020 145.095 ;
        RECT 30.800 144.680 63.020 144.910 ;
        RECT 30.800 144.495 31.420 144.680 ;
        RECT 62.400 144.495 63.020 144.680 ;
        RECT 63.250 144.910 63.870 145.095 ;
        RECT 94.850 144.910 95.470 145.095 ;
        RECT 63.250 144.680 95.470 144.910 ;
        RECT 63.250 144.495 63.870 144.680 ;
        RECT 94.850 144.495 95.470 144.680 ;
        RECT 58.400 144.415 60.020 144.425 ;
        RECT 90.850 144.415 92.470 144.425 ;
        RECT 31.650 144.045 62.170 144.415 ;
        RECT 64.100 144.045 94.620 144.415 ;
        RECT 31.650 143.325 62.170 143.705 ;
        RECT 64.100 143.325 94.620 143.705 ;
        RECT 30.800 143.070 31.420 143.255 ;
        RECT 62.400 143.070 63.020 143.255 ;
        RECT 30.800 142.840 63.020 143.070 ;
        RECT 30.800 142.655 31.420 142.840 ;
        RECT 62.400 142.655 63.020 142.840 ;
        RECT 63.250 143.070 63.870 143.255 ;
        RECT 94.850 143.070 95.470 143.255 ;
        RECT 63.250 142.840 95.470 143.070 ;
        RECT 63.250 142.655 63.870 142.840 ;
        RECT 94.850 142.655 95.470 142.840 ;
        RECT 54.560 142.575 56.180 142.585 ;
        RECT 87.010 142.575 88.630 142.585 ;
        RECT 31.650 142.205 62.170 142.575 ;
        RECT 64.100 142.205 94.620 142.575 ;
        RECT 31.660 141.410 62.160 141.850 ;
        RECT 64.110 141.410 94.610 141.850 ;
        RECT 31.650 140.680 62.170 141.060 ;
        RECT 64.100 140.680 94.620 141.060 ;
        RECT 30.800 140.425 31.420 140.610 ;
        RECT 62.400 140.425 63.020 140.610 ;
        RECT 30.800 140.195 63.020 140.425 ;
        RECT 30.800 140.010 31.420 140.195 ;
        RECT 62.400 140.010 63.020 140.195 ;
        RECT 63.250 140.425 63.870 140.610 ;
        RECT 94.850 140.425 95.470 140.610 ;
        RECT 63.250 140.195 95.470 140.425 ;
        RECT 63.250 140.010 63.870 140.195 ;
        RECT 94.850 140.010 95.470 140.195 ;
        RECT 50.720 139.930 52.340 139.940 ;
        RECT 83.170 139.930 84.790 139.940 ;
        RECT 31.650 139.560 62.170 139.930 ;
        RECT 64.100 139.560 94.620 139.930 ;
        RECT 31.650 138.840 62.170 139.220 ;
        RECT 64.100 138.840 94.620 139.220 ;
        RECT 30.800 138.585 31.420 138.770 ;
        RECT 62.400 138.585 63.020 138.770 ;
        RECT 30.800 138.355 63.020 138.585 ;
        RECT 30.800 138.170 31.420 138.355 ;
        RECT 62.400 138.170 63.020 138.355 ;
        RECT 63.250 138.585 63.870 138.770 ;
        RECT 94.850 138.585 95.470 138.770 ;
        RECT 63.250 138.355 95.470 138.585 ;
        RECT 63.250 138.170 63.870 138.355 ;
        RECT 94.850 138.170 95.470 138.355 ;
        RECT 46.880 138.090 48.500 138.100 ;
        RECT 79.330 138.090 80.950 138.100 ;
        RECT 31.650 137.720 62.170 138.090 ;
        RECT 64.100 137.720 94.620 138.090 ;
        RECT 31.650 137.000 62.170 137.380 ;
        RECT 64.100 137.000 94.620 137.380 ;
        RECT 30.800 136.745 31.420 136.930 ;
        RECT 62.400 136.745 63.020 136.930 ;
        RECT 30.800 136.515 63.020 136.745 ;
        RECT 30.800 136.330 31.420 136.515 ;
        RECT 62.400 136.330 63.020 136.515 ;
        RECT 63.250 136.745 63.870 136.930 ;
        RECT 94.850 136.745 95.470 136.930 ;
        RECT 63.250 136.515 95.470 136.745 ;
        RECT 63.250 136.330 63.870 136.515 ;
        RECT 94.850 136.330 95.470 136.515 ;
        RECT 43.040 136.250 44.660 136.260 ;
        RECT 75.490 136.250 77.110 136.260 ;
        RECT 31.650 135.880 62.170 136.250 ;
        RECT 64.100 135.880 94.620 136.250 ;
        RECT 31.660 135.085 62.160 135.525 ;
        RECT 64.110 135.085 94.610 135.525 ;
        RECT 31.650 134.355 62.170 134.735 ;
        RECT 64.100 134.355 94.620 134.735 ;
        RECT 30.800 134.100 31.420 134.285 ;
        RECT 62.400 134.100 63.020 134.285 ;
        RECT 30.800 133.870 63.020 134.100 ;
        RECT 30.800 133.685 31.420 133.870 ;
        RECT 62.400 133.685 63.020 133.870 ;
        RECT 63.250 134.100 63.870 134.285 ;
        RECT 94.850 134.100 95.470 134.285 ;
        RECT 63.250 133.870 95.470 134.100 ;
        RECT 63.250 133.685 63.870 133.870 ;
        RECT 94.850 133.685 95.470 133.870 ;
        RECT 39.200 133.605 40.820 133.615 ;
        RECT 71.650 133.605 73.270 133.615 ;
        RECT 31.650 133.235 62.170 133.605 ;
        RECT 64.100 133.235 94.620 133.605 ;
        RECT 31.650 132.515 62.170 132.895 ;
        RECT 64.100 132.515 94.620 132.895 ;
        RECT 30.800 132.260 31.420 132.445 ;
        RECT 62.400 132.260 63.020 132.445 ;
        RECT 30.800 132.030 63.020 132.260 ;
        RECT 30.800 131.845 31.420 132.030 ;
        RECT 62.400 131.845 63.020 132.030 ;
        RECT 63.250 132.260 63.870 132.445 ;
        RECT 94.850 132.260 95.470 132.445 ;
        RECT 63.250 132.030 95.470 132.260 ;
        RECT 63.250 131.845 63.870 132.030 ;
        RECT 94.850 131.845 95.470 132.030 ;
        RECT 35.360 131.765 36.980 131.775 ;
        RECT 67.810 131.765 69.430 131.775 ;
        RECT 31.650 131.395 62.170 131.765 ;
        RECT 64.100 131.395 94.620 131.765 ;
        RECT 31.650 130.675 62.170 131.055 ;
        RECT 64.100 130.675 94.620 131.055 ;
        RECT 30.800 130.420 31.420 130.605 ;
        RECT 62.400 130.420 63.020 130.605 ;
        RECT 30.800 130.190 63.020 130.420 ;
        RECT 30.800 130.005 31.420 130.190 ;
        RECT 62.400 130.005 63.020 130.190 ;
        RECT 63.250 130.420 63.870 130.605 ;
        RECT 94.850 130.420 95.470 130.605 ;
        RECT 63.250 130.190 95.470 130.420 ;
        RECT 63.250 130.005 63.870 130.190 ;
        RECT 94.850 130.005 95.470 130.190 ;
        RECT 31.650 129.555 62.170 129.925 ;
        RECT 64.100 129.555 94.620 129.925 ;
        RECT 25.090 127.205 27.380 127.545 ;
        RECT 28.125 127.205 29.610 127.545 ;
        RECT 25.090 126.570 25.690 127.205 ;
        RECT 25.090 126.340 26.670 126.570 ;
        RECT 25.090 124.300 25.690 126.340 ;
        RECT 27.100 126.110 27.460 126.195 ;
        RECT 25.970 125.880 27.460 126.110 ;
        RECT 25.970 125.730 26.330 125.880 ;
        RECT 25.920 125.095 26.870 125.500 ;
        RECT 25.090 124.070 26.380 124.300 ;
        RECT 25.090 123.110 25.690 124.070 ;
        RECT 26.610 123.750 26.870 125.095 ;
        RECT 27.100 124.445 27.460 125.880 ;
        RECT 27.690 124.545 28.040 125.745 ;
        RECT 28.400 125.135 28.780 126.780 ;
        RECT 27.480 123.750 27.830 123.810 ;
        RECT 28.400 123.750 28.740 124.355 ;
        RECT 26.610 123.490 28.740 123.750 ;
        RECT 27.480 123.430 27.830 123.490 ;
        RECT 29.010 123.210 29.610 127.205 ;
        RECT 31.455 126.770 33.205 129.555 ;
        RECT 33.845 126.770 34.655 127.770 ;
        RECT 35.295 126.770 37.045 129.065 ;
        RECT 37.685 126.770 38.495 127.770 ;
        RECT 39.135 126.770 40.885 129.065 ;
        RECT 41.525 126.770 42.335 127.770 ;
        RECT 42.975 126.770 44.725 129.065 ;
        RECT 45.365 126.770 46.175 127.770 ;
        RECT 46.815 126.770 48.565 129.065 ;
        RECT 49.205 126.770 50.015 127.770 ;
        RECT 50.655 126.770 52.405 129.065 ;
        RECT 53.045 126.770 53.855 127.770 ;
        RECT 54.495 126.770 56.245 129.065 ;
        RECT 56.885 126.770 57.695 127.770 ;
        RECT 58.335 126.770 60.085 129.065 ;
        RECT 60.725 126.770 61.535 127.770 ;
        RECT 63.905 126.770 65.655 129.555 ;
        RECT 66.295 126.770 67.105 127.770 ;
        RECT 67.745 126.770 69.495 129.065 ;
        RECT 70.135 126.770 70.945 127.770 ;
        RECT 71.585 126.770 73.335 129.065 ;
        RECT 73.975 126.770 74.785 127.770 ;
        RECT 75.425 126.770 77.175 129.065 ;
        RECT 77.815 126.770 78.625 127.770 ;
        RECT 79.265 126.770 81.015 129.065 ;
        RECT 81.655 126.770 82.465 127.770 ;
        RECT 83.105 126.770 84.855 129.065 ;
        RECT 85.495 126.770 86.305 127.770 ;
        RECT 86.945 126.770 88.695 129.065 ;
        RECT 89.335 126.770 90.145 127.770 ;
        RECT 90.785 126.770 92.535 129.065 ;
        RECT 93.175 126.770 93.985 127.770 ;
        RECT 96.400 126.960 96.770 145.470 ;
        RECT 97.420 141.835 97.790 145.470 ;
        RECT 97.415 141.455 97.795 141.835 ;
        RECT 97.420 138.835 97.790 141.455 ;
        RECT 97.415 138.455 97.795 138.835 ;
        RECT 97.420 135.835 97.790 138.455 ;
        RECT 97.415 135.455 97.795 135.835 ;
        RECT 97.420 132.835 97.790 135.455 ;
        RECT 97.415 132.455 97.795 132.835 ;
        RECT 97.420 129.835 97.790 132.455 ;
        RECT 97.415 129.455 97.795 129.835 ;
        RECT 96.400 126.580 96.780 126.960 ;
        RECT 96.400 125.510 96.770 126.580 ;
        RECT 31.925 124.320 32.735 125.320 ;
        RECT 25.090 122.880 26.780 123.110 ;
        RECT 28.150 122.980 29.610 123.210 ;
        RECT 25.090 120.870 25.690 122.880 ;
        RECT 27.110 122.420 28.110 122.745 ;
        RECT 25.920 121.860 28.780 122.190 ;
        RECT 25.090 120.640 26.780 120.870 ;
        RECT 25.090 118.630 25.690 120.640 ;
        RECT 27.495 120.505 27.760 121.860 ;
        RECT 29.010 120.970 29.610 122.980 ;
        RECT 33.375 122.490 35.125 125.320 ;
        RECT 35.765 124.320 36.575 125.320 ;
        RECT 37.215 123.025 38.965 125.320 ;
        RECT 39.605 124.320 40.415 125.320 ;
        RECT 41.055 123.025 42.805 125.320 ;
        RECT 43.445 124.320 44.255 125.320 ;
        RECT 44.895 123.025 46.645 125.320 ;
        RECT 47.285 124.320 48.095 125.320 ;
        RECT 48.735 123.025 50.485 125.320 ;
        RECT 51.125 124.320 51.935 125.320 ;
        RECT 52.575 123.025 54.325 125.320 ;
        RECT 54.965 124.320 55.775 125.320 ;
        RECT 56.415 123.025 58.165 125.320 ;
        RECT 58.805 124.320 59.615 125.320 ;
        RECT 60.255 123.025 62.005 125.320 ;
        RECT 64.375 124.320 65.185 125.320 ;
        RECT 65.825 122.490 67.575 125.320 ;
        RECT 68.215 124.320 69.025 125.320 ;
        RECT 69.665 123.025 71.415 125.320 ;
        RECT 72.055 124.320 72.865 125.320 ;
        RECT 73.505 123.025 75.255 125.320 ;
        RECT 75.895 124.320 76.705 125.320 ;
        RECT 77.345 123.025 79.095 125.320 ;
        RECT 79.735 124.320 80.545 125.320 ;
        RECT 81.185 123.025 82.935 125.320 ;
        RECT 83.575 124.320 84.385 125.320 ;
        RECT 85.025 123.025 86.775 125.320 ;
        RECT 87.415 124.320 88.225 125.320 ;
        RECT 88.865 123.025 90.615 125.320 ;
        RECT 91.255 124.320 92.065 125.320 ;
        RECT 92.705 123.025 94.455 125.320 ;
        RECT 96.400 125.130 96.780 125.510 ;
        RECT 31.650 122.120 62.170 122.490 ;
        RECT 64.100 122.120 94.620 122.490 ;
        RECT 30.800 121.855 31.420 122.040 ;
        RECT 62.400 121.855 63.020 122.040 ;
        RECT 30.800 121.625 63.020 121.855 ;
        RECT 30.800 121.440 31.420 121.625 ;
        RECT 62.400 121.440 63.020 121.625 ;
        RECT 63.250 121.855 63.870 122.040 ;
        RECT 94.850 121.855 95.470 122.040 ;
        RECT 63.250 121.625 95.470 121.855 ;
        RECT 63.250 121.440 63.870 121.625 ;
        RECT 94.850 121.440 95.470 121.625 ;
        RECT 31.650 120.990 62.170 121.370 ;
        RECT 64.100 120.990 94.620 121.370 ;
        RECT 28.150 120.740 29.610 120.970 ;
        RECT 27.110 120.180 28.110 120.505 ;
        RECT 25.920 119.620 28.780 119.950 ;
        RECT 29.010 118.730 29.610 120.740 ;
        RECT 31.650 120.280 62.170 120.650 ;
        RECT 64.100 120.280 94.620 120.650 ;
        RECT 37.280 120.270 38.900 120.280 ;
        RECT 69.730 120.270 71.350 120.280 ;
        RECT 30.800 120.015 31.420 120.200 ;
        RECT 62.400 120.015 63.020 120.200 ;
        RECT 30.800 119.785 63.020 120.015 ;
        RECT 30.800 119.600 31.420 119.785 ;
        RECT 62.400 119.600 63.020 119.785 ;
        RECT 63.250 120.015 63.870 120.200 ;
        RECT 94.850 120.015 95.470 120.200 ;
        RECT 63.250 119.785 95.470 120.015 ;
        RECT 63.250 119.600 63.870 119.785 ;
        RECT 94.850 119.600 95.470 119.785 ;
        RECT 31.650 119.150 62.170 119.530 ;
        RECT 64.100 119.150 94.620 119.530 ;
        RECT 25.090 118.400 26.780 118.630 ;
        RECT 28.150 118.500 29.610 118.730 ;
        RECT 25.090 116.345 25.690 118.400 ;
        RECT 27.110 117.940 28.110 118.265 ;
        RECT 29.010 116.345 29.610 118.500 ;
        RECT 31.650 118.435 62.170 118.805 ;
        RECT 64.100 118.435 94.620 118.805 ;
        RECT 41.120 118.425 42.740 118.435 ;
        RECT 73.570 118.425 75.190 118.435 ;
        RECT 30.800 118.170 31.420 118.355 ;
        RECT 62.400 118.170 63.020 118.355 ;
        RECT 30.800 117.940 63.020 118.170 ;
        RECT 30.800 117.755 31.420 117.940 ;
        RECT 62.400 117.755 63.020 117.940 ;
        RECT 63.250 118.170 63.870 118.355 ;
        RECT 94.850 118.170 95.470 118.355 ;
        RECT 63.250 117.940 95.470 118.170 ;
        RECT 63.250 117.755 63.870 117.940 ;
        RECT 94.850 117.755 95.470 117.940 ;
        RECT 31.650 117.305 62.170 117.685 ;
        RECT 64.100 117.305 94.620 117.685 ;
        RECT 31.660 116.515 62.160 116.955 ;
        RECT 64.110 116.515 94.610 116.955 ;
        RECT 25.090 116.005 27.380 116.345 ;
        RECT 28.125 116.005 29.610 116.345 ;
        RECT 25.090 88.160 25.690 116.005 ;
        RECT 29.010 88.160 29.610 116.005 ;
        RECT 31.650 115.795 62.170 116.165 ;
        RECT 64.100 115.795 94.620 116.165 ;
        RECT 44.960 115.785 46.580 115.795 ;
        RECT 77.410 115.785 79.030 115.795 ;
        RECT 30.800 115.530 31.420 115.715 ;
        RECT 62.400 115.530 63.020 115.715 ;
        RECT 30.800 115.300 63.020 115.530 ;
        RECT 30.800 115.115 31.420 115.300 ;
        RECT 62.400 115.115 63.020 115.300 ;
        RECT 63.250 115.530 63.870 115.715 ;
        RECT 94.850 115.530 95.470 115.715 ;
        RECT 63.250 115.300 95.470 115.530 ;
        RECT 63.250 115.115 63.870 115.300 ;
        RECT 94.850 115.115 95.470 115.300 ;
        RECT 31.650 114.665 62.170 115.045 ;
        RECT 64.100 114.665 94.620 115.045 ;
        RECT 31.650 113.955 62.170 114.325 ;
        RECT 64.100 113.955 94.620 114.325 ;
        RECT 48.800 113.945 50.420 113.955 ;
        RECT 81.250 113.945 82.870 113.955 ;
        RECT 30.800 113.690 31.420 113.875 ;
        RECT 62.400 113.690 63.020 113.875 ;
        RECT 30.800 113.460 63.020 113.690 ;
        RECT 30.800 113.275 31.420 113.460 ;
        RECT 62.400 113.275 63.020 113.460 ;
        RECT 63.250 113.690 63.870 113.875 ;
        RECT 94.850 113.690 95.470 113.875 ;
        RECT 63.250 113.460 95.470 113.690 ;
        RECT 63.250 113.275 63.870 113.460 ;
        RECT 94.850 113.275 95.470 113.460 ;
        RECT 31.650 112.825 62.170 113.205 ;
        RECT 64.100 112.825 94.620 113.205 ;
        RECT 31.650 112.110 62.170 112.480 ;
        RECT 64.100 112.110 94.620 112.480 ;
        RECT 52.640 112.100 54.260 112.110 ;
        RECT 85.090 112.100 86.710 112.110 ;
        RECT 30.800 111.845 31.420 112.030 ;
        RECT 62.400 111.845 63.020 112.030 ;
        RECT 30.800 111.615 63.020 111.845 ;
        RECT 30.800 111.430 31.420 111.615 ;
        RECT 62.400 111.430 63.020 111.615 ;
        RECT 63.250 111.845 63.870 112.030 ;
        RECT 94.850 111.845 95.470 112.030 ;
        RECT 63.250 111.615 95.470 111.845 ;
        RECT 63.250 111.430 63.870 111.615 ;
        RECT 94.850 111.430 95.470 111.615 ;
        RECT 31.650 110.980 62.170 111.360 ;
        RECT 64.100 110.980 94.620 111.360 ;
        RECT 31.660 110.190 62.160 110.630 ;
        RECT 64.110 110.190 94.610 110.630 ;
        RECT 31.650 109.470 62.170 109.840 ;
        RECT 64.100 109.470 94.620 109.840 ;
        RECT 56.480 109.460 58.100 109.470 ;
        RECT 88.930 109.460 90.550 109.470 ;
        RECT 30.800 109.205 31.420 109.390 ;
        RECT 62.400 109.205 63.020 109.390 ;
        RECT 30.800 108.975 63.020 109.205 ;
        RECT 30.800 108.790 31.420 108.975 ;
        RECT 62.400 108.790 63.020 108.975 ;
        RECT 63.250 109.205 63.870 109.390 ;
        RECT 94.850 109.205 95.470 109.390 ;
        RECT 63.250 108.975 95.470 109.205 ;
        RECT 63.250 108.790 63.870 108.975 ;
        RECT 94.850 108.790 95.470 108.975 ;
        RECT 31.650 108.340 62.170 108.720 ;
        RECT 64.100 108.340 94.620 108.720 ;
        RECT 31.650 107.630 62.170 108.000 ;
        RECT 64.100 107.630 94.620 108.000 ;
        RECT 60.320 107.620 61.940 107.630 ;
        RECT 92.770 107.620 94.390 107.630 ;
        RECT 30.800 107.365 31.420 107.550 ;
        RECT 62.400 107.365 63.020 107.550 ;
        RECT 30.800 107.135 63.020 107.365 ;
        RECT 30.800 106.950 31.420 107.135 ;
        RECT 62.400 106.950 63.020 107.135 ;
        RECT 63.250 107.365 63.870 107.550 ;
        RECT 94.850 107.365 95.470 107.550 ;
        RECT 63.250 107.135 95.470 107.365 ;
        RECT 96.400 107.200 96.770 125.130 ;
        RECT 97.420 123.835 97.790 129.455 ;
        RECT 98.440 126.960 98.810 145.470 ;
        RECT 99.460 141.835 99.830 145.470 ;
        RECT 99.455 141.455 99.835 141.835 ;
        RECT 99.460 138.835 99.830 141.455 ;
        RECT 99.455 138.455 99.835 138.835 ;
        RECT 99.460 135.835 99.830 138.455 ;
        RECT 99.455 135.455 99.835 135.835 ;
        RECT 99.460 132.835 99.830 135.455 ;
        RECT 99.455 132.455 99.835 132.835 ;
        RECT 99.460 129.835 99.830 132.455 ;
        RECT 99.455 129.455 99.835 129.835 ;
        RECT 98.440 126.580 98.820 126.960 ;
        RECT 98.440 125.510 98.810 126.580 ;
        RECT 98.440 125.130 98.820 125.510 ;
        RECT 97.415 123.455 97.795 123.835 ;
        RECT 97.420 120.835 97.790 123.455 ;
        RECT 97.415 120.455 97.795 120.835 ;
        RECT 97.420 117.835 97.790 120.455 ;
        RECT 97.415 117.455 97.795 117.835 ;
        RECT 97.420 114.835 97.790 117.455 ;
        RECT 97.415 114.455 97.795 114.835 ;
        RECT 97.420 111.835 97.790 114.455 ;
        RECT 97.415 111.455 97.795 111.835 ;
        RECT 97.420 108.835 97.790 111.455 ;
        RECT 97.415 108.455 97.795 108.835 ;
        RECT 97.420 107.200 97.790 108.455 ;
        RECT 98.440 107.200 98.810 125.130 ;
        RECT 99.460 123.835 99.830 129.455 ;
        RECT 99.455 123.455 99.835 123.835 ;
        RECT 99.460 120.835 99.830 123.455 ;
        RECT 99.455 120.455 99.835 120.835 ;
        RECT 99.460 117.835 99.830 120.455 ;
        RECT 99.455 117.455 99.835 117.835 ;
        RECT 99.460 114.835 99.830 117.455 ;
        RECT 99.455 114.455 99.835 114.835 ;
        RECT 99.460 111.835 99.830 114.455 ;
        RECT 99.455 111.455 99.835 111.835 ;
        RECT 99.460 108.835 99.830 111.455 ;
        RECT 99.455 108.455 99.835 108.835 ;
        RECT 99.460 107.200 99.830 108.455 ;
        RECT 100.480 107.200 100.860 145.470 ;
        RECT 101.210 107.210 101.650 145.460 ;
        RECT 63.250 106.950 63.870 107.135 ;
        RECT 94.850 106.950 95.470 107.135 ;
        RECT 31.650 106.500 62.170 106.880 ;
        RECT 64.100 106.500 94.620 106.880 ;
        RECT 31.650 105.780 62.170 106.160 ;
        RECT 64.100 105.780 94.620 106.160 ;
        RECT 30.800 105.525 31.420 105.710 ;
        RECT 62.400 105.525 63.020 105.710 ;
        RECT 30.800 105.295 63.020 105.525 ;
        RECT 30.800 105.110 31.420 105.295 ;
        RECT 62.400 105.110 63.020 105.295 ;
        RECT 63.250 105.525 63.870 105.710 ;
        RECT 94.850 105.525 95.470 105.710 ;
        RECT 63.250 105.295 95.470 105.525 ;
        RECT 63.250 105.110 63.870 105.295 ;
        RECT 94.850 105.110 95.470 105.295 ;
        RECT 58.400 105.030 60.020 105.040 ;
        RECT 90.850 105.030 92.470 105.040 ;
        RECT 31.650 104.660 62.170 105.030 ;
        RECT 64.100 104.660 94.620 105.030 ;
        RECT 31.650 103.940 62.170 104.320 ;
        RECT 64.100 103.940 94.620 104.320 ;
        RECT 30.800 103.685 31.420 103.870 ;
        RECT 62.400 103.685 63.020 103.870 ;
        RECT 30.800 103.455 63.020 103.685 ;
        RECT 30.800 103.270 31.420 103.455 ;
        RECT 62.400 103.270 63.020 103.455 ;
        RECT 63.250 103.685 63.870 103.870 ;
        RECT 94.850 103.685 95.470 103.870 ;
        RECT 63.250 103.455 95.470 103.685 ;
        RECT 63.250 103.270 63.870 103.455 ;
        RECT 94.850 103.270 95.470 103.455 ;
        RECT 54.560 103.190 56.180 103.200 ;
        RECT 87.010 103.190 88.630 103.200 ;
        RECT 31.650 102.820 62.170 103.190 ;
        RECT 64.100 102.820 94.620 103.190 ;
        RECT 31.660 102.025 62.160 102.465 ;
        RECT 64.110 102.025 94.610 102.465 ;
        RECT 31.650 101.295 62.170 101.675 ;
        RECT 64.100 101.295 94.620 101.675 ;
        RECT 30.800 101.040 31.420 101.225 ;
        RECT 62.400 101.040 63.020 101.225 ;
        RECT 30.800 100.810 63.020 101.040 ;
        RECT 30.800 100.625 31.420 100.810 ;
        RECT 62.400 100.625 63.020 100.810 ;
        RECT 63.250 101.040 63.870 101.225 ;
        RECT 94.850 101.040 95.470 101.225 ;
        RECT 63.250 100.810 95.470 101.040 ;
        RECT 63.250 100.625 63.870 100.810 ;
        RECT 94.850 100.625 95.470 100.810 ;
        RECT 50.720 100.545 52.340 100.555 ;
        RECT 83.170 100.545 84.790 100.555 ;
        RECT 31.650 100.175 62.170 100.545 ;
        RECT 64.100 100.175 94.620 100.545 ;
        RECT 31.650 99.455 62.170 99.835 ;
        RECT 64.100 99.455 94.620 99.835 ;
        RECT 30.800 99.200 31.420 99.385 ;
        RECT 62.400 99.200 63.020 99.385 ;
        RECT 30.800 98.970 63.020 99.200 ;
        RECT 30.800 98.785 31.420 98.970 ;
        RECT 62.400 98.785 63.020 98.970 ;
        RECT 63.250 99.200 63.870 99.385 ;
        RECT 94.850 99.200 95.470 99.385 ;
        RECT 63.250 98.970 95.470 99.200 ;
        RECT 63.250 98.785 63.870 98.970 ;
        RECT 94.850 98.785 95.470 98.970 ;
        RECT 46.880 98.705 48.500 98.715 ;
        RECT 79.330 98.705 80.950 98.715 ;
        RECT 31.650 98.335 62.170 98.705 ;
        RECT 64.100 98.335 94.620 98.705 ;
        RECT 31.650 97.615 62.170 97.995 ;
        RECT 64.100 97.615 94.620 97.995 ;
        RECT 30.800 97.360 31.420 97.545 ;
        RECT 62.400 97.360 63.020 97.545 ;
        RECT 30.800 97.130 63.020 97.360 ;
        RECT 30.800 96.945 31.420 97.130 ;
        RECT 62.400 96.945 63.020 97.130 ;
        RECT 63.250 97.360 63.870 97.545 ;
        RECT 94.850 97.360 95.470 97.545 ;
        RECT 63.250 97.130 95.470 97.360 ;
        RECT 63.250 96.945 63.870 97.130 ;
        RECT 94.850 96.945 95.470 97.130 ;
        RECT 43.040 96.865 44.660 96.875 ;
        RECT 75.490 96.865 77.110 96.875 ;
        RECT 31.650 96.495 62.170 96.865 ;
        RECT 64.100 96.495 94.620 96.865 ;
        RECT 31.660 95.700 62.160 96.140 ;
        RECT 64.110 95.700 94.610 96.140 ;
        RECT 31.650 94.970 62.170 95.350 ;
        RECT 64.100 94.970 94.620 95.350 ;
        RECT 30.800 94.715 31.420 94.900 ;
        RECT 62.400 94.715 63.020 94.900 ;
        RECT 30.800 94.485 63.020 94.715 ;
        RECT 30.800 94.300 31.420 94.485 ;
        RECT 62.400 94.300 63.020 94.485 ;
        RECT 63.250 94.715 63.870 94.900 ;
        RECT 94.850 94.715 95.470 94.900 ;
        RECT 63.250 94.485 95.470 94.715 ;
        RECT 63.250 94.300 63.870 94.485 ;
        RECT 94.850 94.300 95.470 94.485 ;
        RECT 39.200 94.220 40.820 94.230 ;
        RECT 71.650 94.220 73.270 94.230 ;
        RECT 31.650 93.850 62.170 94.220 ;
        RECT 64.100 93.850 94.620 94.220 ;
        RECT 31.650 93.130 62.170 93.510 ;
        RECT 64.100 93.130 94.620 93.510 ;
        RECT 30.800 92.875 31.420 93.060 ;
        RECT 62.400 92.875 63.020 93.060 ;
        RECT 30.800 92.645 63.020 92.875 ;
        RECT 30.800 92.460 31.420 92.645 ;
        RECT 62.400 92.460 63.020 92.645 ;
        RECT 63.250 92.875 63.870 93.060 ;
        RECT 94.850 92.875 95.470 93.060 ;
        RECT 63.250 92.645 95.470 92.875 ;
        RECT 63.250 92.460 63.870 92.645 ;
        RECT 94.850 92.460 95.470 92.645 ;
        RECT 35.360 92.380 36.980 92.390 ;
        RECT 67.810 92.380 69.430 92.390 ;
        RECT 31.650 92.010 62.170 92.380 ;
        RECT 64.100 92.010 94.620 92.380 ;
        RECT 31.650 91.290 62.170 91.670 ;
        RECT 64.100 91.290 94.620 91.670 ;
        RECT 30.800 91.035 31.420 91.220 ;
        RECT 62.400 91.035 63.020 91.220 ;
        RECT 30.800 90.805 63.020 91.035 ;
        RECT 30.800 90.620 31.420 90.805 ;
        RECT 62.400 90.620 63.020 90.805 ;
        RECT 63.250 91.035 63.870 91.220 ;
        RECT 94.850 91.035 95.470 91.220 ;
        RECT 63.250 90.805 95.470 91.035 ;
        RECT 63.250 90.620 63.870 90.805 ;
        RECT 94.850 90.620 95.470 90.805 ;
        RECT 31.650 90.170 62.170 90.540 ;
        RECT 64.100 90.170 94.620 90.540 ;
        RECT 25.090 87.820 27.380 88.160 ;
        RECT 28.125 87.820 29.610 88.160 ;
        RECT 25.090 87.185 25.690 87.820 ;
        RECT 25.090 86.955 26.670 87.185 ;
        RECT 25.090 84.915 25.690 86.955 ;
        RECT 27.100 86.725 27.460 86.810 ;
        RECT 25.970 86.495 27.460 86.725 ;
        RECT 25.970 86.345 26.330 86.495 ;
        RECT 25.920 85.710 26.870 86.115 ;
        RECT 25.090 84.685 26.380 84.915 ;
        RECT 25.090 83.725 25.690 84.685 ;
        RECT 26.610 84.365 26.870 85.710 ;
        RECT 27.100 85.060 27.460 86.495 ;
        RECT 27.690 85.160 28.040 86.360 ;
        RECT 28.400 85.750 28.780 87.395 ;
        RECT 27.480 84.365 27.830 84.425 ;
        RECT 28.400 84.365 28.740 84.970 ;
        RECT 26.610 84.105 28.740 84.365 ;
        RECT 27.480 84.045 27.830 84.105 ;
        RECT 29.010 83.825 29.610 87.820 ;
        RECT 31.455 87.385 33.205 90.170 ;
        RECT 33.845 87.385 34.655 88.385 ;
        RECT 35.295 87.385 37.045 89.680 ;
        RECT 37.685 87.385 38.495 88.385 ;
        RECT 39.135 87.385 40.885 89.680 ;
        RECT 41.525 87.385 42.335 88.385 ;
        RECT 42.975 87.385 44.725 89.680 ;
        RECT 45.365 87.385 46.175 88.385 ;
        RECT 46.815 87.385 48.565 89.680 ;
        RECT 49.205 87.385 50.015 88.385 ;
        RECT 50.655 87.385 52.405 89.680 ;
        RECT 53.045 87.385 53.855 88.385 ;
        RECT 54.495 87.385 56.245 89.680 ;
        RECT 56.885 87.385 57.695 88.385 ;
        RECT 58.335 87.385 60.085 89.680 ;
        RECT 60.725 87.385 61.535 88.385 ;
        RECT 63.905 87.385 65.655 90.170 ;
        RECT 66.295 87.385 67.105 88.385 ;
        RECT 67.745 87.385 69.495 89.680 ;
        RECT 70.135 87.385 70.945 88.385 ;
        RECT 71.585 87.385 73.335 89.680 ;
        RECT 73.975 87.385 74.785 88.385 ;
        RECT 75.425 87.385 77.175 89.680 ;
        RECT 77.815 87.385 78.625 88.385 ;
        RECT 79.265 87.385 81.015 89.680 ;
        RECT 81.655 87.385 82.465 88.385 ;
        RECT 83.105 87.385 84.855 89.680 ;
        RECT 85.495 87.385 86.305 88.385 ;
        RECT 86.945 87.385 88.695 89.680 ;
        RECT 89.335 87.385 90.145 88.385 ;
        RECT 90.785 87.385 92.535 89.680 ;
        RECT 93.175 87.385 93.985 88.385 ;
        RECT 96.400 87.575 96.770 106.085 ;
        RECT 97.420 102.450 97.790 106.085 ;
        RECT 97.415 102.070 97.795 102.450 ;
        RECT 97.420 99.450 97.790 102.070 ;
        RECT 97.415 99.070 97.795 99.450 ;
        RECT 97.420 96.450 97.790 99.070 ;
        RECT 97.415 96.070 97.795 96.450 ;
        RECT 97.420 93.450 97.790 96.070 ;
        RECT 97.415 93.070 97.795 93.450 ;
        RECT 97.420 90.450 97.790 93.070 ;
        RECT 97.415 90.070 97.795 90.450 ;
        RECT 96.400 87.195 96.780 87.575 ;
        RECT 96.400 86.125 96.770 87.195 ;
        RECT 31.925 84.935 32.735 85.935 ;
        RECT 25.090 83.495 26.780 83.725 ;
        RECT 28.150 83.595 29.610 83.825 ;
        RECT 25.090 81.485 25.690 83.495 ;
        RECT 27.110 83.035 28.110 83.360 ;
        RECT 25.920 82.475 28.780 82.805 ;
        RECT 25.090 81.255 26.780 81.485 ;
        RECT 25.090 79.245 25.690 81.255 ;
        RECT 27.495 81.120 27.760 82.475 ;
        RECT 29.010 81.585 29.610 83.595 ;
        RECT 33.375 83.105 35.125 85.935 ;
        RECT 35.765 84.935 36.575 85.935 ;
        RECT 37.215 83.640 38.965 85.935 ;
        RECT 39.605 84.935 40.415 85.935 ;
        RECT 41.055 83.640 42.805 85.935 ;
        RECT 43.445 84.935 44.255 85.935 ;
        RECT 44.895 83.640 46.645 85.935 ;
        RECT 47.285 84.935 48.095 85.935 ;
        RECT 48.735 83.640 50.485 85.935 ;
        RECT 51.125 84.935 51.935 85.935 ;
        RECT 52.575 83.640 54.325 85.935 ;
        RECT 54.965 84.935 55.775 85.935 ;
        RECT 56.415 83.640 58.165 85.935 ;
        RECT 58.805 84.935 59.615 85.935 ;
        RECT 60.255 83.640 62.005 85.935 ;
        RECT 64.375 84.935 65.185 85.935 ;
        RECT 65.825 83.105 67.575 85.935 ;
        RECT 68.215 84.935 69.025 85.935 ;
        RECT 69.665 83.640 71.415 85.935 ;
        RECT 72.055 84.935 72.865 85.935 ;
        RECT 73.505 83.640 75.255 85.935 ;
        RECT 75.895 84.935 76.705 85.935 ;
        RECT 77.345 83.640 79.095 85.935 ;
        RECT 79.735 84.935 80.545 85.935 ;
        RECT 81.185 83.640 82.935 85.935 ;
        RECT 83.575 84.935 84.385 85.935 ;
        RECT 85.025 83.640 86.775 85.935 ;
        RECT 87.415 84.935 88.225 85.935 ;
        RECT 88.865 83.640 90.615 85.935 ;
        RECT 91.255 84.935 92.065 85.935 ;
        RECT 92.705 83.640 94.455 85.935 ;
        RECT 96.400 85.745 96.780 86.125 ;
        RECT 31.650 82.735 62.170 83.105 ;
        RECT 64.100 82.735 94.620 83.105 ;
        RECT 30.800 82.470 31.420 82.655 ;
        RECT 62.400 82.470 63.020 82.655 ;
        RECT 30.800 82.240 63.020 82.470 ;
        RECT 30.800 82.055 31.420 82.240 ;
        RECT 62.400 82.055 63.020 82.240 ;
        RECT 63.250 82.470 63.870 82.655 ;
        RECT 94.850 82.470 95.470 82.655 ;
        RECT 63.250 82.240 95.470 82.470 ;
        RECT 63.250 82.055 63.870 82.240 ;
        RECT 94.850 82.055 95.470 82.240 ;
        RECT 31.650 81.605 62.170 81.985 ;
        RECT 64.100 81.605 94.620 81.985 ;
        RECT 28.150 81.355 29.610 81.585 ;
        RECT 27.110 80.795 28.110 81.120 ;
        RECT 25.920 80.235 28.780 80.565 ;
        RECT 29.010 79.345 29.610 81.355 ;
        RECT 31.650 80.895 62.170 81.265 ;
        RECT 64.100 80.895 94.620 81.265 ;
        RECT 37.280 80.885 38.900 80.895 ;
        RECT 69.730 80.885 71.350 80.895 ;
        RECT 30.800 80.630 31.420 80.815 ;
        RECT 62.400 80.630 63.020 80.815 ;
        RECT 30.800 80.400 63.020 80.630 ;
        RECT 30.800 80.215 31.420 80.400 ;
        RECT 62.400 80.215 63.020 80.400 ;
        RECT 63.250 80.630 63.870 80.815 ;
        RECT 94.850 80.630 95.470 80.815 ;
        RECT 63.250 80.400 95.470 80.630 ;
        RECT 63.250 80.215 63.870 80.400 ;
        RECT 94.850 80.215 95.470 80.400 ;
        RECT 31.650 79.765 62.170 80.145 ;
        RECT 64.100 79.765 94.620 80.145 ;
        RECT 25.090 79.015 26.780 79.245 ;
        RECT 28.150 79.115 29.610 79.345 ;
        RECT 25.090 76.960 25.690 79.015 ;
        RECT 27.110 78.555 28.110 78.880 ;
        RECT 29.010 76.960 29.610 79.115 ;
        RECT 31.650 79.050 62.170 79.420 ;
        RECT 64.100 79.050 94.620 79.420 ;
        RECT 41.120 79.040 42.740 79.050 ;
        RECT 73.570 79.040 75.190 79.050 ;
        RECT 30.800 78.785 31.420 78.970 ;
        RECT 62.400 78.785 63.020 78.970 ;
        RECT 30.800 78.555 63.020 78.785 ;
        RECT 30.800 78.370 31.420 78.555 ;
        RECT 62.400 78.370 63.020 78.555 ;
        RECT 63.250 78.785 63.870 78.970 ;
        RECT 94.850 78.785 95.470 78.970 ;
        RECT 63.250 78.555 95.470 78.785 ;
        RECT 63.250 78.370 63.870 78.555 ;
        RECT 94.850 78.370 95.470 78.555 ;
        RECT 31.650 77.920 62.170 78.300 ;
        RECT 64.100 77.920 94.620 78.300 ;
        RECT 31.660 77.130 62.160 77.570 ;
        RECT 64.110 77.130 94.610 77.570 ;
        RECT 25.090 76.620 27.380 76.960 ;
        RECT 28.125 76.620 29.610 76.960 ;
        RECT 25.090 66.885 25.690 76.620 ;
        RECT 29.010 66.885 29.610 76.620 ;
        RECT 31.650 76.410 62.170 76.780 ;
        RECT 64.100 76.410 94.620 76.780 ;
        RECT 44.960 76.400 46.580 76.410 ;
        RECT 77.410 76.400 79.030 76.410 ;
        RECT 30.800 76.145 31.420 76.330 ;
        RECT 62.400 76.145 63.020 76.330 ;
        RECT 30.800 75.915 63.020 76.145 ;
        RECT 30.800 75.730 31.420 75.915 ;
        RECT 62.400 75.730 63.020 75.915 ;
        RECT 63.250 76.145 63.870 76.330 ;
        RECT 94.850 76.145 95.470 76.330 ;
        RECT 63.250 75.915 95.470 76.145 ;
        RECT 63.250 75.730 63.870 75.915 ;
        RECT 94.850 75.730 95.470 75.915 ;
        RECT 31.650 75.280 62.170 75.660 ;
        RECT 64.100 75.280 94.620 75.660 ;
        RECT 31.650 74.570 62.170 74.940 ;
        RECT 64.100 74.570 94.620 74.940 ;
        RECT 48.800 74.560 50.420 74.570 ;
        RECT 81.250 74.560 82.870 74.570 ;
        RECT 30.800 74.305 31.420 74.490 ;
        RECT 62.400 74.305 63.020 74.490 ;
        RECT 30.800 74.075 63.020 74.305 ;
        RECT 30.800 73.890 31.420 74.075 ;
        RECT 62.400 73.890 63.020 74.075 ;
        RECT 63.250 74.305 63.870 74.490 ;
        RECT 94.850 74.305 95.470 74.490 ;
        RECT 63.250 74.075 95.470 74.305 ;
        RECT 63.250 73.890 63.870 74.075 ;
        RECT 94.850 73.890 95.470 74.075 ;
        RECT 31.650 73.440 62.170 73.820 ;
        RECT 64.100 73.440 94.620 73.820 ;
        RECT 31.650 72.725 62.170 73.095 ;
        RECT 64.100 72.725 94.620 73.095 ;
        RECT 52.640 72.715 54.260 72.725 ;
        RECT 85.090 72.715 86.710 72.725 ;
        RECT 30.800 72.460 31.420 72.645 ;
        RECT 62.400 72.460 63.020 72.645 ;
        RECT 30.800 72.230 63.020 72.460 ;
        RECT 30.800 72.045 31.420 72.230 ;
        RECT 62.400 72.045 63.020 72.230 ;
        RECT 63.250 72.460 63.870 72.645 ;
        RECT 94.850 72.460 95.470 72.645 ;
        RECT 63.250 72.230 95.470 72.460 ;
        RECT 63.250 72.045 63.870 72.230 ;
        RECT 94.850 72.045 95.470 72.230 ;
        RECT 31.650 71.595 62.170 71.975 ;
        RECT 64.100 71.595 94.620 71.975 ;
        RECT 31.660 70.805 62.160 71.245 ;
        RECT 64.110 70.805 94.610 71.245 ;
        RECT 31.650 70.085 62.170 70.455 ;
        RECT 64.100 70.085 94.620 70.455 ;
        RECT 56.480 70.075 58.100 70.085 ;
        RECT 88.930 70.075 90.550 70.085 ;
        RECT 30.800 69.820 31.420 70.005 ;
        RECT 62.400 69.820 63.020 70.005 ;
        RECT 30.800 69.590 63.020 69.820 ;
        RECT 30.800 69.405 31.420 69.590 ;
        RECT 62.400 69.405 63.020 69.590 ;
        RECT 63.250 69.820 63.870 70.005 ;
        RECT 94.850 69.820 95.470 70.005 ;
        RECT 63.250 69.590 95.470 69.820 ;
        RECT 63.250 69.405 63.870 69.590 ;
        RECT 94.850 69.405 95.470 69.590 ;
        RECT 31.650 68.955 62.170 69.335 ;
        RECT 64.100 68.955 94.620 69.335 ;
        RECT 31.650 68.245 62.170 68.615 ;
        RECT 64.100 68.245 94.620 68.615 ;
        RECT 60.320 68.235 61.940 68.245 ;
        RECT 92.770 68.235 94.390 68.245 ;
        RECT 30.800 67.980 31.420 68.165 ;
        RECT 62.400 67.980 63.020 68.165 ;
        RECT 30.800 67.750 63.020 67.980 ;
        RECT 30.800 67.565 31.420 67.750 ;
        RECT 62.400 67.565 63.020 67.750 ;
        RECT 63.250 67.980 63.870 68.165 ;
        RECT 94.850 67.980 95.470 68.165 ;
        RECT 63.250 67.750 95.470 67.980 ;
        RECT 96.400 67.815 96.770 85.745 ;
        RECT 97.420 84.450 97.790 90.070 ;
        RECT 98.440 87.575 98.810 106.085 ;
        RECT 99.460 102.450 99.830 106.085 ;
        RECT 99.455 102.070 99.835 102.450 ;
        RECT 99.460 99.450 99.830 102.070 ;
        RECT 99.455 99.070 99.835 99.450 ;
        RECT 99.460 96.450 99.830 99.070 ;
        RECT 99.455 96.070 99.835 96.450 ;
        RECT 99.460 93.450 99.830 96.070 ;
        RECT 99.455 93.070 99.835 93.450 ;
        RECT 99.460 90.450 99.830 93.070 ;
        RECT 99.455 90.070 99.835 90.450 ;
        RECT 98.440 87.195 98.820 87.575 ;
        RECT 98.440 86.125 98.810 87.195 ;
        RECT 98.440 85.745 98.820 86.125 ;
        RECT 97.415 84.070 97.795 84.450 ;
        RECT 97.420 81.450 97.790 84.070 ;
        RECT 97.415 81.070 97.795 81.450 ;
        RECT 97.420 78.450 97.790 81.070 ;
        RECT 97.415 78.070 97.795 78.450 ;
        RECT 97.420 75.450 97.790 78.070 ;
        RECT 97.415 75.070 97.795 75.450 ;
        RECT 97.420 72.450 97.790 75.070 ;
        RECT 97.415 72.070 97.795 72.450 ;
        RECT 97.420 69.450 97.790 72.070 ;
        RECT 97.415 69.070 97.795 69.450 ;
        RECT 97.420 67.815 97.790 69.070 ;
        RECT 98.440 67.815 98.810 85.745 ;
        RECT 99.460 84.450 99.830 90.070 ;
        RECT 99.455 84.070 99.835 84.450 ;
        RECT 99.460 81.450 99.830 84.070 ;
        RECT 99.455 81.070 99.835 81.450 ;
        RECT 99.460 78.450 99.830 81.070 ;
        RECT 99.455 78.070 99.835 78.450 ;
        RECT 99.460 75.450 99.830 78.070 ;
        RECT 99.455 75.070 99.835 75.450 ;
        RECT 99.460 72.450 99.830 75.070 ;
        RECT 99.455 72.070 99.835 72.450 ;
        RECT 99.460 69.450 99.830 72.070 ;
        RECT 99.455 69.070 99.835 69.450 ;
        RECT 99.460 67.815 99.830 69.070 ;
        RECT 100.480 67.815 100.860 106.085 ;
        RECT 101.210 67.825 101.650 106.075 ;
        RECT 63.250 67.565 63.870 67.750 ;
        RECT 94.850 67.565 95.470 67.750 ;
        RECT 31.650 67.115 62.170 67.495 ;
        RECT 64.100 67.115 94.620 67.495 ;
      LAYER Metal2 ;
        RECT 31.920 381.475 34.160 381.855 ;
        RECT 64.370 381.475 66.610 381.855 ;
        RECT 62.520 380.915 62.900 381.295 ;
        RECT 94.970 380.915 95.350 381.295 ;
        RECT 25.200 379.265 25.580 379.645 ;
        RECT 29.120 379.265 29.500 379.645 ;
        RECT 31.920 379.635 34.160 380.015 ;
        RECT 31.925 377.750 34.165 378.130 ;
        RECT 31.920 376.990 34.160 377.370 ;
        RECT 25.200 376.265 25.580 376.645 ;
        RECT 29.120 376.265 29.500 376.645 ;
        RECT 31.920 375.150 34.160 375.530 ;
        RECT 25.200 373.265 25.580 373.645 ;
        RECT 29.120 373.265 29.500 373.645 ;
        RECT 31.920 373.310 34.160 373.690 ;
        RECT 31.925 371.425 34.165 371.805 ;
        RECT 31.920 370.665 34.160 371.045 ;
        RECT 25.200 370.265 25.580 370.645 ;
        RECT 29.120 370.265 29.500 370.645 ;
        RECT 31.920 368.825 34.160 369.205 ;
        RECT 25.200 367.265 25.580 367.645 ;
        RECT 29.120 367.265 29.500 367.645 ;
        RECT 31.920 366.985 34.160 367.365 ;
        RECT 25.200 364.265 25.580 364.645 ;
        RECT 29.120 364.265 29.500 364.645 ;
        RECT 35.295 364.275 37.045 368.085 ;
        RECT 39.135 364.275 40.885 369.925 ;
        RECT 42.975 364.275 44.725 372.570 ;
        RECT 46.815 364.275 48.565 374.410 ;
        RECT 50.655 364.275 52.405 376.250 ;
        RECT 54.495 364.275 56.245 378.895 ;
        RECT 58.335 364.275 60.085 380.735 ;
        RECT 64.370 379.635 66.610 380.015 ;
        RECT 62.520 379.075 62.900 379.455 ;
        RECT 64.375 377.750 66.615 378.130 ;
        RECT 64.370 376.990 66.610 377.370 ;
        RECT 62.520 376.430 62.900 376.810 ;
        RECT 64.370 375.150 66.610 375.530 ;
        RECT 62.520 374.590 62.900 374.970 ;
        RECT 64.370 373.310 66.610 373.690 ;
        RECT 62.520 372.750 62.900 373.130 ;
        RECT 64.375 371.425 66.615 371.805 ;
        RECT 64.370 370.665 66.610 371.045 ;
        RECT 62.520 370.105 62.900 370.485 ;
        RECT 64.370 368.825 66.610 369.205 ;
        RECT 62.520 368.265 62.900 368.645 ;
        RECT 64.370 366.985 66.610 367.365 ;
        RECT 62.520 366.425 62.900 366.805 ;
        RECT 67.745 364.275 69.495 368.085 ;
        RECT 71.585 364.275 73.335 369.925 ;
        RECT 75.425 364.275 77.175 372.570 ;
        RECT 79.265 364.275 81.015 374.410 ;
        RECT 83.105 364.275 84.855 376.250 ;
        RECT 86.945 364.275 88.695 378.895 ;
        RECT 90.785 364.275 92.535 380.735 ;
        RECT 94.970 379.075 95.350 379.455 ;
        RECT 97.415 377.765 97.795 378.145 ;
        RECT 99.455 377.765 99.835 378.145 ;
        RECT 101.240 377.765 101.620 378.145 ;
        RECT 94.970 376.430 95.350 376.810 ;
        RECT 94.970 374.590 95.350 374.970 ;
        RECT 97.415 374.765 97.795 375.145 ;
        RECT 99.455 374.765 99.835 375.145 ;
        RECT 101.240 374.765 101.620 375.145 ;
        RECT 94.970 372.750 95.350 373.130 ;
        RECT 97.415 371.765 97.795 372.145 ;
        RECT 99.455 371.765 99.835 372.145 ;
        RECT 101.240 371.765 101.620 372.145 ;
        RECT 94.970 370.105 95.350 370.485 ;
        RECT 97.415 368.765 97.795 369.145 ;
        RECT 99.455 368.765 99.835 369.145 ;
        RECT 101.240 368.765 101.620 369.145 ;
        RECT 94.970 368.265 95.350 368.645 ;
        RECT 94.970 366.425 95.350 366.805 ;
        RECT 97.415 365.765 97.795 366.145 ;
        RECT 99.455 365.765 99.835 366.145 ;
        RECT 101.240 365.765 101.620 366.145 ;
        RECT 34.060 363.890 34.440 364.080 ;
        RECT 37.900 363.890 38.280 364.080 ;
        RECT 41.740 363.890 42.120 364.080 ;
        RECT 45.580 363.890 45.960 364.080 ;
        RECT 49.420 363.890 49.800 364.080 ;
        RECT 53.260 363.890 53.640 364.080 ;
        RECT 57.100 363.890 57.480 364.080 ;
        RECT 60.940 363.890 61.320 364.080 ;
        RECT 66.510 363.890 66.890 364.080 ;
        RECT 70.350 363.890 70.730 364.080 ;
        RECT 74.190 363.890 74.570 364.080 ;
        RECT 78.030 363.890 78.410 364.080 ;
        RECT 81.870 363.890 82.250 364.080 ;
        RECT 85.710 363.890 86.090 364.080 ;
        RECT 89.550 363.890 89.930 364.080 ;
        RECT 93.390 363.890 93.770 364.080 ;
        RECT 28.390 363.080 101.890 363.890 ;
        RECT 25.200 361.265 25.580 361.645 ;
        RECT 28.390 361.630 29.200 363.080 ;
        RECT 96.400 362.890 96.780 363.080 ;
        RECT 98.440 362.890 98.820 363.080 ;
        RECT 100.480 362.890 100.860 363.080 ;
        RECT 96.400 361.630 96.780 361.820 ;
        RECT 98.440 361.630 98.820 361.820 ;
        RECT 100.480 361.630 100.860 361.820 ;
        RECT 28.390 360.820 101.890 361.630 ;
        RECT 32.140 360.630 32.520 360.820 ;
        RECT 35.980 360.630 36.360 360.820 ;
        RECT 39.820 360.630 40.200 360.820 ;
        RECT 43.660 360.630 44.040 360.820 ;
        RECT 47.500 360.630 47.880 360.820 ;
        RECT 51.340 360.630 51.720 360.820 ;
        RECT 55.180 360.630 55.560 360.820 ;
        RECT 59.020 360.630 59.400 360.820 ;
        RECT 64.590 360.630 64.970 360.820 ;
        RECT 68.430 360.630 68.810 360.820 ;
        RECT 72.270 360.630 72.650 360.820 ;
        RECT 76.110 360.630 76.490 360.820 ;
        RECT 79.950 360.630 80.330 360.820 ;
        RECT 83.790 360.630 84.170 360.820 ;
        RECT 87.630 360.630 88.010 360.820 ;
        RECT 91.470 360.630 91.850 360.820 ;
        RECT 25.200 358.265 25.580 358.645 ;
        RECT 27.480 355.930 27.830 360.120 ;
        RECT 25.200 355.265 25.580 355.645 ;
        RECT 28.110 354.575 28.460 358.490 ;
        RECT 29.120 358.265 29.500 358.645 ;
        RECT 31.920 357.300 34.160 357.680 ;
        RECT 37.215 356.580 38.965 360.435 ;
        RECT 29.120 355.265 29.500 355.645 ;
        RECT 31.920 355.460 34.160 355.840 ;
        RECT 41.055 354.735 42.805 360.435 ;
        RECT 27.705 354.250 28.460 354.575 ;
        RECT 28.110 354.245 28.460 354.250 ;
        RECT 31.920 353.615 34.160 353.995 ;
        RECT 31.925 352.855 34.165 353.235 ;
        RECT 25.200 352.265 25.580 352.645 ;
        RECT 29.120 352.265 29.500 352.645 ;
        RECT 44.895 352.095 46.645 360.435 ;
        RECT 31.920 350.975 34.160 351.355 ;
        RECT 48.735 350.255 50.485 360.435 ;
        RECT 25.200 349.265 25.580 349.645 ;
        RECT 29.120 349.265 29.500 349.645 ;
        RECT 31.920 349.135 34.160 349.515 ;
        RECT 52.575 348.410 54.325 360.435 ;
        RECT 31.920 347.290 34.160 347.670 ;
        RECT 25.200 346.265 25.580 346.645 ;
        RECT 29.120 346.265 29.500 346.645 ;
        RECT 31.925 346.530 34.165 346.910 ;
        RECT 56.415 345.770 58.165 360.435 ;
        RECT 31.920 344.650 34.160 345.030 ;
        RECT 60.255 343.930 62.005 360.435 ;
        RECT 62.520 357.860 62.900 358.240 ;
        RECT 64.370 357.300 66.610 357.680 ;
        RECT 69.665 356.580 71.415 360.435 ;
        RECT 62.520 356.020 62.900 356.400 ;
        RECT 64.370 355.460 66.610 355.840 ;
        RECT 73.505 354.735 75.255 360.435 ;
        RECT 62.520 354.175 62.900 354.555 ;
        RECT 64.370 353.615 66.610 353.995 ;
        RECT 64.375 352.855 66.615 353.235 ;
        RECT 77.345 352.095 79.095 360.435 ;
        RECT 62.520 351.535 62.900 351.915 ;
        RECT 64.370 350.975 66.610 351.355 ;
        RECT 81.185 350.255 82.935 360.435 ;
        RECT 62.520 349.695 62.900 350.075 ;
        RECT 64.370 349.135 66.610 349.515 ;
        RECT 85.025 348.410 86.775 360.435 ;
        RECT 62.520 347.850 62.900 348.230 ;
        RECT 64.370 347.290 66.610 347.670 ;
        RECT 64.375 346.530 66.615 346.910 ;
        RECT 88.865 345.770 90.615 360.435 ;
        RECT 62.520 345.210 62.900 345.590 ;
        RECT 64.370 344.650 66.610 345.030 ;
        RECT 92.705 343.930 94.455 360.435 ;
        RECT 97.415 359.765 97.795 360.145 ;
        RECT 99.455 359.765 99.835 360.145 ;
        RECT 101.240 359.765 101.620 360.145 ;
        RECT 94.970 357.860 95.350 358.240 ;
        RECT 97.415 356.765 97.795 357.145 ;
        RECT 99.455 356.765 99.835 357.145 ;
        RECT 101.240 356.765 101.620 357.145 ;
        RECT 94.970 356.020 95.350 356.400 ;
        RECT 94.970 354.175 95.350 354.555 ;
        RECT 97.415 353.765 97.795 354.145 ;
        RECT 99.455 353.765 99.835 354.145 ;
        RECT 101.240 353.765 101.620 354.145 ;
        RECT 94.970 351.535 95.350 351.915 ;
        RECT 97.415 350.765 97.795 351.145 ;
        RECT 99.455 350.765 99.835 351.145 ;
        RECT 101.240 350.765 101.620 351.145 ;
        RECT 94.970 349.695 95.350 350.075 ;
        RECT 94.970 347.850 95.350 348.230 ;
        RECT 97.415 347.765 97.795 348.145 ;
        RECT 99.455 347.765 99.835 348.145 ;
        RECT 101.240 347.765 101.620 348.145 ;
        RECT 94.970 345.210 95.350 345.590 ;
        RECT 97.415 344.765 97.795 345.145 ;
        RECT 99.455 344.765 99.835 345.145 ;
        RECT 101.240 344.765 101.620 345.145 ;
        RECT 25.200 343.265 25.580 343.645 ;
        RECT 29.120 343.265 29.500 343.645 ;
        RECT 62.520 343.370 62.900 343.750 ;
        RECT 94.970 343.370 95.350 343.750 ;
        RECT 31.920 342.810 34.160 343.190 ;
        RECT 64.370 342.810 66.610 343.190 ;
        RECT 31.920 342.090 34.160 342.470 ;
        RECT 64.370 342.090 66.610 342.470 ;
        RECT 62.520 341.530 62.900 341.910 ;
        RECT 94.970 341.530 95.350 341.910 ;
        RECT 25.200 339.880 25.580 340.260 ;
        RECT 29.120 339.880 29.500 340.260 ;
        RECT 31.920 340.250 34.160 340.630 ;
        RECT 31.925 338.365 34.165 338.745 ;
        RECT 31.920 337.605 34.160 337.985 ;
        RECT 25.200 336.880 25.580 337.260 ;
        RECT 29.120 336.880 29.500 337.260 ;
        RECT 31.920 335.765 34.160 336.145 ;
        RECT 25.200 333.880 25.580 334.260 ;
        RECT 29.120 333.880 29.500 334.260 ;
        RECT 31.920 333.925 34.160 334.305 ;
        RECT 31.925 332.040 34.165 332.420 ;
        RECT 31.920 331.280 34.160 331.660 ;
        RECT 25.200 330.880 25.580 331.260 ;
        RECT 29.120 330.880 29.500 331.260 ;
        RECT 31.920 329.440 34.160 329.820 ;
        RECT 25.200 327.880 25.580 328.260 ;
        RECT 29.120 327.880 29.500 328.260 ;
        RECT 31.920 327.600 34.160 327.980 ;
        RECT 25.200 324.880 25.580 325.260 ;
        RECT 29.120 324.880 29.500 325.260 ;
        RECT 35.295 324.890 37.045 328.700 ;
        RECT 39.135 324.890 40.885 330.540 ;
        RECT 42.975 324.890 44.725 333.185 ;
        RECT 46.815 324.890 48.565 335.025 ;
        RECT 50.655 324.890 52.405 336.865 ;
        RECT 54.495 324.890 56.245 339.510 ;
        RECT 58.335 324.890 60.085 341.350 ;
        RECT 64.370 340.250 66.610 340.630 ;
        RECT 62.520 339.690 62.900 340.070 ;
        RECT 64.375 338.365 66.615 338.745 ;
        RECT 64.370 337.605 66.610 337.985 ;
        RECT 62.520 337.045 62.900 337.425 ;
        RECT 64.370 335.765 66.610 336.145 ;
        RECT 62.520 335.205 62.900 335.585 ;
        RECT 64.370 333.925 66.610 334.305 ;
        RECT 62.520 333.365 62.900 333.745 ;
        RECT 64.375 332.040 66.615 332.420 ;
        RECT 64.370 331.280 66.610 331.660 ;
        RECT 62.520 330.720 62.900 331.100 ;
        RECT 64.370 329.440 66.610 329.820 ;
        RECT 62.520 328.880 62.900 329.260 ;
        RECT 64.370 327.600 66.610 327.980 ;
        RECT 62.520 327.040 62.900 327.420 ;
        RECT 67.745 324.890 69.495 328.700 ;
        RECT 71.585 324.890 73.335 330.540 ;
        RECT 75.425 324.890 77.175 333.185 ;
        RECT 79.265 324.890 81.015 335.025 ;
        RECT 83.105 324.890 84.855 336.865 ;
        RECT 86.945 324.890 88.695 339.510 ;
        RECT 90.785 324.890 92.535 341.350 ;
        RECT 94.970 339.690 95.350 340.070 ;
        RECT 97.415 338.380 97.795 338.760 ;
        RECT 99.455 338.380 99.835 338.760 ;
        RECT 101.240 338.380 101.620 338.760 ;
        RECT 94.970 337.045 95.350 337.425 ;
        RECT 94.970 335.205 95.350 335.585 ;
        RECT 97.415 335.380 97.795 335.760 ;
        RECT 99.455 335.380 99.835 335.760 ;
        RECT 101.240 335.380 101.620 335.760 ;
        RECT 94.970 333.365 95.350 333.745 ;
        RECT 97.415 332.380 97.795 332.760 ;
        RECT 99.455 332.380 99.835 332.760 ;
        RECT 101.240 332.380 101.620 332.760 ;
        RECT 94.970 330.720 95.350 331.100 ;
        RECT 97.415 329.380 97.795 329.760 ;
        RECT 99.455 329.380 99.835 329.760 ;
        RECT 101.240 329.380 101.620 329.760 ;
        RECT 94.970 328.880 95.350 329.260 ;
        RECT 94.970 327.040 95.350 327.420 ;
        RECT 97.415 326.380 97.795 326.760 ;
        RECT 99.455 326.380 99.835 326.760 ;
        RECT 101.240 326.380 101.620 326.760 ;
        RECT 34.060 324.505 34.440 324.695 ;
        RECT 37.900 324.505 38.280 324.695 ;
        RECT 41.740 324.505 42.120 324.695 ;
        RECT 45.580 324.505 45.960 324.695 ;
        RECT 49.420 324.505 49.800 324.695 ;
        RECT 53.260 324.505 53.640 324.695 ;
        RECT 57.100 324.505 57.480 324.695 ;
        RECT 60.940 324.505 61.320 324.695 ;
        RECT 66.510 324.505 66.890 324.695 ;
        RECT 70.350 324.505 70.730 324.695 ;
        RECT 74.190 324.505 74.570 324.695 ;
        RECT 78.030 324.505 78.410 324.695 ;
        RECT 81.870 324.505 82.250 324.695 ;
        RECT 85.710 324.505 86.090 324.695 ;
        RECT 89.550 324.505 89.930 324.695 ;
        RECT 93.390 324.505 93.770 324.695 ;
        RECT 28.390 323.695 101.890 324.505 ;
        RECT 25.200 321.880 25.580 322.260 ;
        RECT 28.390 322.245 29.200 323.695 ;
        RECT 96.400 323.505 96.780 323.695 ;
        RECT 98.440 323.505 98.820 323.695 ;
        RECT 100.480 323.505 100.860 323.695 ;
        RECT 96.400 322.245 96.780 322.435 ;
        RECT 98.440 322.245 98.820 322.435 ;
        RECT 100.480 322.245 100.860 322.435 ;
        RECT 28.390 321.435 101.890 322.245 ;
        RECT 32.140 321.245 32.520 321.435 ;
        RECT 35.980 321.245 36.360 321.435 ;
        RECT 39.820 321.245 40.200 321.435 ;
        RECT 43.660 321.245 44.040 321.435 ;
        RECT 47.500 321.245 47.880 321.435 ;
        RECT 51.340 321.245 51.720 321.435 ;
        RECT 55.180 321.245 55.560 321.435 ;
        RECT 59.020 321.245 59.400 321.435 ;
        RECT 64.590 321.245 64.970 321.435 ;
        RECT 68.430 321.245 68.810 321.435 ;
        RECT 72.270 321.245 72.650 321.435 ;
        RECT 76.110 321.245 76.490 321.435 ;
        RECT 79.950 321.245 80.330 321.435 ;
        RECT 83.790 321.245 84.170 321.435 ;
        RECT 87.630 321.245 88.010 321.435 ;
        RECT 91.470 321.245 91.850 321.435 ;
        RECT 25.200 318.880 25.580 319.260 ;
        RECT 27.480 316.545 27.830 320.735 ;
        RECT 25.200 315.880 25.580 316.260 ;
        RECT 28.110 315.190 28.460 319.105 ;
        RECT 29.120 318.880 29.500 319.260 ;
        RECT 31.920 317.915 34.160 318.295 ;
        RECT 37.215 317.195 38.965 321.050 ;
        RECT 29.120 315.880 29.500 316.260 ;
        RECT 31.920 316.075 34.160 316.455 ;
        RECT 41.055 315.350 42.805 321.050 ;
        RECT 27.705 314.865 28.460 315.190 ;
        RECT 28.110 314.860 28.460 314.865 ;
        RECT 31.920 314.230 34.160 314.610 ;
        RECT 31.925 313.470 34.165 313.850 ;
        RECT 25.200 312.880 25.580 313.260 ;
        RECT 29.120 312.880 29.500 313.260 ;
        RECT 44.895 312.710 46.645 321.050 ;
        RECT 31.920 311.590 34.160 311.970 ;
        RECT 48.735 310.870 50.485 321.050 ;
        RECT 25.200 309.880 25.580 310.260 ;
        RECT 29.120 309.880 29.500 310.260 ;
        RECT 31.920 309.750 34.160 310.130 ;
        RECT 52.575 309.025 54.325 321.050 ;
        RECT 31.920 307.905 34.160 308.285 ;
        RECT 25.200 306.880 25.580 307.260 ;
        RECT 29.120 306.880 29.500 307.260 ;
        RECT 31.925 307.145 34.165 307.525 ;
        RECT 56.415 306.385 58.165 321.050 ;
        RECT 31.920 305.265 34.160 305.645 ;
        RECT 60.255 304.545 62.005 321.050 ;
        RECT 62.520 318.475 62.900 318.855 ;
        RECT 64.370 317.915 66.610 318.295 ;
        RECT 69.665 317.195 71.415 321.050 ;
        RECT 62.520 316.635 62.900 317.015 ;
        RECT 64.370 316.075 66.610 316.455 ;
        RECT 73.505 315.350 75.255 321.050 ;
        RECT 62.520 314.790 62.900 315.170 ;
        RECT 64.370 314.230 66.610 314.610 ;
        RECT 64.375 313.470 66.615 313.850 ;
        RECT 77.345 312.710 79.095 321.050 ;
        RECT 62.520 312.150 62.900 312.530 ;
        RECT 64.370 311.590 66.610 311.970 ;
        RECT 81.185 310.870 82.935 321.050 ;
        RECT 62.520 310.310 62.900 310.690 ;
        RECT 64.370 309.750 66.610 310.130 ;
        RECT 85.025 309.025 86.775 321.050 ;
        RECT 62.520 308.465 62.900 308.845 ;
        RECT 64.370 307.905 66.610 308.285 ;
        RECT 64.375 307.145 66.615 307.525 ;
        RECT 88.865 306.385 90.615 321.050 ;
        RECT 62.520 305.825 62.900 306.205 ;
        RECT 64.370 305.265 66.610 305.645 ;
        RECT 92.705 304.545 94.455 321.050 ;
        RECT 97.415 320.380 97.795 320.760 ;
        RECT 99.455 320.380 99.835 320.760 ;
        RECT 101.240 320.380 101.620 320.760 ;
        RECT 94.970 318.475 95.350 318.855 ;
        RECT 97.415 317.380 97.795 317.760 ;
        RECT 99.455 317.380 99.835 317.760 ;
        RECT 101.240 317.380 101.620 317.760 ;
        RECT 94.970 316.635 95.350 317.015 ;
        RECT 94.970 314.790 95.350 315.170 ;
        RECT 97.415 314.380 97.795 314.760 ;
        RECT 99.455 314.380 99.835 314.760 ;
        RECT 101.240 314.380 101.620 314.760 ;
        RECT 94.970 312.150 95.350 312.530 ;
        RECT 97.415 311.380 97.795 311.760 ;
        RECT 99.455 311.380 99.835 311.760 ;
        RECT 101.240 311.380 101.620 311.760 ;
        RECT 94.970 310.310 95.350 310.690 ;
        RECT 94.970 308.465 95.350 308.845 ;
        RECT 97.415 308.380 97.795 308.760 ;
        RECT 99.455 308.380 99.835 308.760 ;
        RECT 101.240 308.380 101.620 308.760 ;
        RECT 94.970 305.825 95.350 306.205 ;
        RECT 97.415 305.380 97.795 305.760 ;
        RECT 99.455 305.380 99.835 305.760 ;
        RECT 101.240 305.380 101.620 305.760 ;
        RECT 25.200 303.880 25.580 304.260 ;
        RECT 29.120 303.880 29.500 304.260 ;
        RECT 62.520 303.985 62.900 304.365 ;
        RECT 94.970 303.985 95.350 304.365 ;
        RECT 31.920 303.425 34.160 303.805 ;
        RECT 64.370 303.425 66.610 303.805 ;
        RECT 31.920 302.705 34.160 303.085 ;
        RECT 64.370 302.705 66.610 303.085 ;
        RECT 62.520 302.145 62.900 302.525 ;
        RECT 94.970 302.145 95.350 302.525 ;
        RECT 25.200 300.495 25.580 300.875 ;
        RECT 29.120 300.495 29.500 300.875 ;
        RECT 31.920 300.865 34.160 301.245 ;
        RECT 31.925 298.980 34.165 299.360 ;
        RECT 31.920 298.220 34.160 298.600 ;
        RECT 25.200 297.495 25.580 297.875 ;
        RECT 29.120 297.495 29.500 297.875 ;
        RECT 31.920 296.380 34.160 296.760 ;
        RECT 25.200 294.495 25.580 294.875 ;
        RECT 29.120 294.495 29.500 294.875 ;
        RECT 31.920 294.540 34.160 294.920 ;
        RECT 31.925 292.655 34.165 293.035 ;
        RECT 31.920 291.895 34.160 292.275 ;
        RECT 25.200 291.495 25.580 291.875 ;
        RECT 29.120 291.495 29.500 291.875 ;
        RECT 31.920 290.055 34.160 290.435 ;
        RECT 25.200 288.495 25.580 288.875 ;
        RECT 29.120 288.495 29.500 288.875 ;
        RECT 31.920 288.215 34.160 288.595 ;
        RECT 25.200 285.495 25.580 285.875 ;
        RECT 29.120 285.495 29.500 285.875 ;
        RECT 35.295 285.505 37.045 289.315 ;
        RECT 39.135 285.505 40.885 291.155 ;
        RECT 42.975 285.505 44.725 293.800 ;
        RECT 46.815 285.505 48.565 295.640 ;
        RECT 50.655 285.505 52.405 297.480 ;
        RECT 54.495 285.505 56.245 300.125 ;
        RECT 58.335 285.505 60.085 301.965 ;
        RECT 64.370 300.865 66.610 301.245 ;
        RECT 62.520 300.305 62.900 300.685 ;
        RECT 64.375 298.980 66.615 299.360 ;
        RECT 64.370 298.220 66.610 298.600 ;
        RECT 62.520 297.660 62.900 298.040 ;
        RECT 64.370 296.380 66.610 296.760 ;
        RECT 62.520 295.820 62.900 296.200 ;
        RECT 64.370 294.540 66.610 294.920 ;
        RECT 62.520 293.980 62.900 294.360 ;
        RECT 64.375 292.655 66.615 293.035 ;
        RECT 64.370 291.895 66.610 292.275 ;
        RECT 62.520 291.335 62.900 291.715 ;
        RECT 64.370 290.055 66.610 290.435 ;
        RECT 62.520 289.495 62.900 289.875 ;
        RECT 64.370 288.215 66.610 288.595 ;
        RECT 62.520 287.655 62.900 288.035 ;
        RECT 67.745 285.505 69.495 289.315 ;
        RECT 71.585 285.505 73.335 291.155 ;
        RECT 75.425 285.505 77.175 293.800 ;
        RECT 79.265 285.505 81.015 295.640 ;
        RECT 83.105 285.505 84.855 297.480 ;
        RECT 86.945 285.505 88.695 300.125 ;
        RECT 90.785 285.505 92.535 301.965 ;
        RECT 94.970 300.305 95.350 300.685 ;
        RECT 97.415 298.995 97.795 299.375 ;
        RECT 99.455 298.995 99.835 299.375 ;
        RECT 101.240 298.995 101.620 299.375 ;
        RECT 94.970 297.660 95.350 298.040 ;
        RECT 94.970 295.820 95.350 296.200 ;
        RECT 97.415 295.995 97.795 296.375 ;
        RECT 99.455 295.995 99.835 296.375 ;
        RECT 101.240 295.995 101.620 296.375 ;
        RECT 94.970 293.980 95.350 294.360 ;
        RECT 97.415 292.995 97.795 293.375 ;
        RECT 99.455 292.995 99.835 293.375 ;
        RECT 101.240 292.995 101.620 293.375 ;
        RECT 94.970 291.335 95.350 291.715 ;
        RECT 97.415 289.995 97.795 290.375 ;
        RECT 99.455 289.995 99.835 290.375 ;
        RECT 101.240 289.995 101.620 290.375 ;
        RECT 94.970 289.495 95.350 289.875 ;
        RECT 94.970 287.655 95.350 288.035 ;
        RECT 97.415 286.995 97.795 287.375 ;
        RECT 99.455 286.995 99.835 287.375 ;
        RECT 101.240 286.995 101.620 287.375 ;
        RECT 34.060 285.120 34.440 285.310 ;
        RECT 37.900 285.120 38.280 285.310 ;
        RECT 41.740 285.120 42.120 285.310 ;
        RECT 45.580 285.120 45.960 285.310 ;
        RECT 49.420 285.120 49.800 285.310 ;
        RECT 53.260 285.120 53.640 285.310 ;
        RECT 57.100 285.120 57.480 285.310 ;
        RECT 60.940 285.120 61.320 285.310 ;
        RECT 66.510 285.120 66.890 285.310 ;
        RECT 70.350 285.120 70.730 285.310 ;
        RECT 74.190 285.120 74.570 285.310 ;
        RECT 78.030 285.120 78.410 285.310 ;
        RECT 81.870 285.120 82.250 285.310 ;
        RECT 85.710 285.120 86.090 285.310 ;
        RECT 89.550 285.120 89.930 285.310 ;
        RECT 93.390 285.120 93.770 285.310 ;
        RECT 28.390 284.310 101.890 285.120 ;
        RECT 25.200 282.495 25.580 282.875 ;
        RECT 28.390 282.860 29.200 284.310 ;
        RECT 96.400 284.120 96.780 284.310 ;
        RECT 98.440 284.120 98.820 284.310 ;
        RECT 100.480 284.120 100.860 284.310 ;
        RECT 96.400 282.860 96.780 283.050 ;
        RECT 98.440 282.860 98.820 283.050 ;
        RECT 100.480 282.860 100.860 283.050 ;
        RECT 28.390 282.050 101.890 282.860 ;
        RECT 32.140 281.860 32.520 282.050 ;
        RECT 35.980 281.860 36.360 282.050 ;
        RECT 39.820 281.860 40.200 282.050 ;
        RECT 43.660 281.860 44.040 282.050 ;
        RECT 47.500 281.860 47.880 282.050 ;
        RECT 51.340 281.860 51.720 282.050 ;
        RECT 55.180 281.860 55.560 282.050 ;
        RECT 59.020 281.860 59.400 282.050 ;
        RECT 64.590 281.860 64.970 282.050 ;
        RECT 68.430 281.860 68.810 282.050 ;
        RECT 72.270 281.860 72.650 282.050 ;
        RECT 76.110 281.860 76.490 282.050 ;
        RECT 79.950 281.860 80.330 282.050 ;
        RECT 83.790 281.860 84.170 282.050 ;
        RECT 87.630 281.860 88.010 282.050 ;
        RECT 91.470 281.860 91.850 282.050 ;
        RECT 25.200 279.495 25.580 279.875 ;
        RECT 27.480 277.160 27.830 281.350 ;
        RECT 25.200 276.495 25.580 276.875 ;
        RECT 28.110 275.805 28.460 279.720 ;
        RECT 29.120 279.495 29.500 279.875 ;
        RECT 31.920 278.530 34.160 278.910 ;
        RECT 37.215 277.810 38.965 281.665 ;
        RECT 29.120 276.495 29.500 276.875 ;
        RECT 31.920 276.690 34.160 277.070 ;
        RECT 41.055 275.965 42.805 281.665 ;
        RECT 27.705 275.480 28.460 275.805 ;
        RECT 28.110 275.475 28.460 275.480 ;
        RECT 31.920 274.845 34.160 275.225 ;
        RECT 31.925 274.085 34.165 274.465 ;
        RECT 25.200 273.495 25.580 273.875 ;
        RECT 29.120 273.495 29.500 273.875 ;
        RECT 44.895 273.325 46.645 281.665 ;
        RECT 31.920 272.205 34.160 272.585 ;
        RECT 48.735 271.485 50.485 281.665 ;
        RECT 25.200 270.495 25.580 270.875 ;
        RECT 29.120 270.495 29.500 270.875 ;
        RECT 31.920 270.365 34.160 270.745 ;
        RECT 52.575 269.640 54.325 281.665 ;
        RECT 31.920 268.520 34.160 268.900 ;
        RECT 25.200 267.495 25.580 267.875 ;
        RECT 29.120 267.495 29.500 267.875 ;
        RECT 31.925 267.760 34.165 268.140 ;
        RECT 56.415 267.000 58.165 281.665 ;
        RECT 31.920 265.880 34.160 266.260 ;
        RECT 60.255 265.160 62.005 281.665 ;
        RECT 62.520 279.090 62.900 279.470 ;
        RECT 64.370 278.530 66.610 278.910 ;
        RECT 69.665 277.810 71.415 281.665 ;
        RECT 62.520 277.250 62.900 277.630 ;
        RECT 64.370 276.690 66.610 277.070 ;
        RECT 73.505 275.965 75.255 281.665 ;
        RECT 62.520 275.405 62.900 275.785 ;
        RECT 64.370 274.845 66.610 275.225 ;
        RECT 64.375 274.085 66.615 274.465 ;
        RECT 77.345 273.325 79.095 281.665 ;
        RECT 62.520 272.765 62.900 273.145 ;
        RECT 64.370 272.205 66.610 272.585 ;
        RECT 81.185 271.485 82.935 281.665 ;
        RECT 62.520 270.925 62.900 271.305 ;
        RECT 64.370 270.365 66.610 270.745 ;
        RECT 85.025 269.640 86.775 281.665 ;
        RECT 62.520 269.080 62.900 269.460 ;
        RECT 64.370 268.520 66.610 268.900 ;
        RECT 64.375 267.760 66.615 268.140 ;
        RECT 88.865 267.000 90.615 281.665 ;
        RECT 62.520 266.440 62.900 266.820 ;
        RECT 64.370 265.880 66.610 266.260 ;
        RECT 92.705 265.160 94.455 281.665 ;
        RECT 97.415 280.995 97.795 281.375 ;
        RECT 99.455 280.995 99.835 281.375 ;
        RECT 101.240 280.995 101.620 281.375 ;
        RECT 94.970 279.090 95.350 279.470 ;
        RECT 97.415 277.995 97.795 278.375 ;
        RECT 99.455 277.995 99.835 278.375 ;
        RECT 101.240 277.995 101.620 278.375 ;
        RECT 94.970 277.250 95.350 277.630 ;
        RECT 94.970 275.405 95.350 275.785 ;
        RECT 97.415 274.995 97.795 275.375 ;
        RECT 99.455 274.995 99.835 275.375 ;
        RECT 101.240 274.995 101.620 275.375 ;
        RECT 94.970 272.765 95.350 273.145 ;
        RECT 97.415 271.995 97.795 272.375 ;
        RECT 99.455 271.995 99.835 272.375 ;
        RECT 101.240 271.995 101.620 272.375 ;
        RECT 94.970 270.925 95.350 271.305 ;
        RECT 94.970 269.080 95.350 269.460 ;
        RECT 97.415 268.995 97.795 269.375 ;
        RECT 99.455 268.995 99.835 269.375 ;
        RECT 101.240 268.995 101.620 269.375 ;
        RECT 94.970 266.440 95.350 266.820 ;
        RECT 97.415 265.995 97.795 266.375 ;
        RECT 99.455 265.995 99.835 266.375 ;
        RECT 101.240 265.995 101.620 266.375 ;
        RECT 25.200 264.495 25.580 264.875 ;
        RECT 29.120 264.495 29.500 264.875 ;
        RECT 62.520 264.600 62.900 264.980 ;
        RECT 94.970 264.600 95.350 264.980 ;
        RECT 31.920 264.040 34.160 264.420 ;
        RECT 64.370 264.040 66.610 264.420 ;
        RECT 31.920 263.320 34.160 263.700 ;
        RECT 64.370 263.320 66.610 263.700 ;
        RECT 62.520 262.760 62.900 263.140 ;
        RECT 94.970 262.760 95.350 263.140 ;
        RECT 25.200 261.110 25.580 261.490 ;
        RECT 29.120 261.110 29.500 261.490 ;
        RECT 31.920 261.480 34.160 261.860 ;
        RECT 31.925 259.595 34.165 259.975 ;
        RECT 31.920 258.835 34.160 259.215 ;
        RECT 25.200 258.110 25.580 258.490 ;
        RECT 29.120 258.110 29.500 258.490 ;
        RECT 31.920 256.995 34.160 257.375 ;
        RECT 25.200 255.110 25.580 255.490 ;
        RECT 29.120 255.110 29.500 255.490 ;
        RECT 31.920 255.155 34.160 255.535 ;
        RECT 31.925 253.270 34.165 253.650 ;
        RECT 31.920 252.510 34.160 252.890 ;
        RECT 25.200 252.110 25.580 252.490 ;
        RECT 29.120 252.110 29.500 252.490 ;
        RECT 31.920 250.670 34.160 251.050 ;
        RECT 25.200 249.110 25.580 249.490 ;
        RECT 29.120 249.110 29.500 249.490 ;
        RECT 31.920 248.830 34.160 249.210 ;
        RECT 25.200 246.110 25.580 246.490 ;
        RECT 29.120 246.110 29.500 246.490 ;
        RECT 35.295 246.120 37.045 249.930 ;
        RECT 39.135 246.120 40.885 251.770 ;
        RECT 42.975 246.120 44.725 254.415 ;
        RECT 46.815 246.120 48.565 256.255 ;
        RECT 50.655 246.120 52.405 258.095 ;
        RECT 54.495 246.120 56.245 260.740 ;
        RECT 58.335 246.120 60.085 262.580 ;
        RECT 64.370 261.480 66.610 261.860 ;
        RECT 62.520 260.920 62.900 261.300 ;
        RECT 64.375 259.595 66.615 259.975 ;
        RECT 64.370 258.835 66.610 259.215 ;
        RECT 62.520 258.275 62.900 258.655 ;
        RECT 64.370 256.995 66.610 257.375 ;
        RECT 62.520 256.435 62.900 256.815 ;
        RECT 64.370 255.155 66.610 255.535 ;
        RECT 62.520 254.595 62.900 254.975 ;
        RECT 64.375 253.270 66.615 253.650 ;
        RECT 64.370 252.510 66.610 252.890 ;
        RECT 62.520 251.950 62.900 252.330 ;
        RECT 64.370 250.670 66.610 251.050 ;
        RECT 62.520 250.110 62.900 250.490 ;
        RECT 64.370 248.830 66.610 249.210 ;
        RECT 62.520 248.270 62.900 248.650 ;
        RECT 67.745 246.120 69.495 249.930 ;
        RECT 71.585 246.120 73.335 251.770 ;
        RECT 75.425 246.120 77.175 254.415 ;
        RECT 79.265 246.120 81.015 256.255 ;
        RECT 83.105 246.120 84.855 258.095 ;
        RECT 86.945 246.120 88.695 260.740 ;
        RECT 90.785 246.120 92.535 262.580 ;
        RECT 94.970 260.920 95.350 261.300 ;
        RECT 97.415 259.610 97.795 259.990 ;
        RECT 99.455 259.610 99.835 259.990 ;
        RECT 101.240 259.610 101.620 259.990 ;
        RECT 94.970 258.275 95.350 258.655 ;
        RECT 94.970 256.435 95.350 256.815 ;
        RECT 97.415 256.610 97.795 256.990 ;
        RECT 99.455 256.610 99.835 256.990 ;
        RECT 101.240 256.610 101.620 256.990 ;
        RECT 94.970 254.595 95.350 254.975 ;
        RECT 97.415 253.610 97.795 253.990 ;
        RECT 99.455 253.610 99.835 253.990 ;
        RECT 101.240 253.610 101.620 253.990 ;
        RECT 94.970 251.950 95.350 252.330 ;
        RECT 97.415 250.610 97.795 250.990 ;
        RECT 99.455 250.610 99.835 250.990 ;
        RECT 101.240 250.610 101.620 250.990 ;
        RECT 94.970 250.110 95.350 250.490 ;
        RECT 94.970 248.270 95.350 248.650 ;
        RECT 97.415 247.610 97.795 247.990 ;
        RECT 99.455 247.610 99.835 247.990 ;
        RECT 101.240 247.610 101.620 247.990 ;
        RECT 34.060 245.735 34.440 245.925 ;
        RECT 37.900 245.735 38.280 245.925 ;
        RECT 41.740 245.735 42.120 245.925 ;
        RECT 45.580 245.735 45.960 245.925 ;
        RECT 49.420 245.735 49.800 245.925 ;
        RECT 53.260 245.735 53.640 245.925 ;
        RECT 57.100 245.735 57.480 245.925 ;
        RECT 60.940 245.735 61.320 245.925 ;
        RECT 66.510 245.735 66.890 245.925 ;
        RECT 70.350 245.735 70.730 245.925 ;
        RECT 74.190 245.735 74.570 245.925 ;
        RECT 78.030 245.735 78.410 245.925 ;
        RECT 81.870 245.735 82.250 245.925 ;
        RECT 85.710 245.735 86.090 245.925 ;
        RECT 89.550 245.735 89.930 245.925 ;
        RECT 93.390 245.735 93.770 245.925 ;
        RECT 28.390 244.925 101.890 245.735 ;
        RECT 25.200 243.110 25.580 243.490 ;
        RECT 28.390 243.475 29.200 244.925 ;
        RECT 96.400 244.735 96.780 244.925 ;
        RECT 98.440 244.735 98.820 244.925 ;
        RECT 100.480 244.735 100.860 244.925 ;
        RECT 96.400 243.475 96.780 243.665 ;
        RECT 98.440 243.475 98.820 243.665 ;
        RECT 100.480 243.475 100.860 243.665 ;
        RECT 28.390 242.665 101.890 243.475 ;
        RECT 32.140 242.475 32.520 242.665 ;
        RECT 35.980 242.475 36.360 242.665 ;
        RECT 39.820 242.475 40.200 242.665 ;
        RECT 43.660 242.475 44.040 242.665 ;
        RECT 47.500 242.475 47.880 242.665 ;
        RECT 51.340 242.475 51.720 242.665 ;
        RECT 55.180 242.475 55.560 242.665 ;
        RECT 59.020 242.475 59.400 242.665 ;
        RECT 64.590 242.475 64.970 242.665 ;
        RECT 68.430 242.475 68.810 242.665 ;
        RECT 72.270 242.475 72.650 242.665 ;
        RECT 76.110 242.475 76.490 242.665 ;
        RECT 79.950 242.475 80.330 242.665 ;
        RECT 83.790 242.475 84.170 242.665 ;
        RECT 87.630 242.475 88.010 242.665 ;
        RECT 91.470 242.475 91.850 242.665 ;
        RECT 25.200 240.110 25.580 240.490 ;
        RECT 27.480 237.775 27.830 241.965 ;
        RECT 25.200 237.110 25.580 237.490 ;
        RECT 28.110 236.420 28.460 240.335 ;
        RECT 29.120 240.110 29.500 240.490 ;
        RECT 31.920 239.145 34.160 239.525 ;
        RECT 37.215 238.425 38.965 242.280 ;
        RECT 29.120 237.110 29.500 237.490 ;
        RECT 31.920 237.305 34.160 237.685 ;
        RECT 41.055 236.580 42.805 242.280 ;
        RECT 27.705 236.095 28.460 236.420 ;
        RECT 28.110 236.090 28.460 236.095 ;
        RECT 31.920 235.460 34.160 235.840 ;
        RECT 31.925 234.700 34.165 235.080 ;
        RECT 25.200 234.110 25.580 234.490 ;
        RECT 29.120 234.110 29.500 234.490 ;
        RECT 44.895 233.940 46.645 242.280 ;
        RECT 31.920 232.820 34.160 233.200 ;
        RECT 48.735 232.100 50.485 242.280 ;
        RECT 25.200 231.110 25.580 231.490 ;
        RECT 29.120 231.110 29.500 231.490 ;
        RECT 31.920 230.980 34.160 231.360 ;
        RECT 52.575 230.255 54.325 242.280 ;
        RECT 31.920 229.135 34.160 229.515 ;
        RECT 25.200 228.110 25.580 228.490 ;
        RECT 29.120 228.110 29.500 228.490 ;
        RECT 31.925 228.375 34.165 228.755 ;
        RECT 56.415 227.615 58.165 242.280 ;
        RECT 31.920 226.495 34.160 226.875 ;
        RECT 60.255 225.775 62.005 242.280 ;
        RECT 62.520 239.705 62.900 240.085 ;
        RECT 64.370 239.145 66.610 239.525 ;
        RECT 69.665 238.425 71.415 242.280 ;
        RECT 62.520 237.865 62.900 238.245 ;
        RECT 64.370 237.305 66.610 237.685 ;
        RECT 73.505 236.580 75.255 242.280 ;
        RECT 62.520 236.020 62.900 236.400 ;
        RECT 64.370 235.460 66.610 235.840 ;
        RECT 64.375 234.700 66.615 235.080 ;
        RECT 77.345 233.940 79.095 242.280 ;
        RECT 62.520 233.380 62.900 233.760 ;
        RECT 64.370 232.820 66.610 233.200 ;
        RECT 81.185 232.100 82.935 242.280 ;
        RECT 62.520 231.540 62.900 231.920 ;
        RECT 64.370 230.980 66.610 231.360 ;
        RECT 85.025 230.255 86.775 242.280 ;
        RECT 62.520 229.695 62.900 230.075 ;
        RECT 64.370 229.135 66.610 229.515 ;
        RECT 64.375 228.375 66.615 228.755 ;
        RECT 88.865 227.615 90.615 242.280 ;
        RECT 62.520 227.055 62.900 227.435 ;
        RECT 64.370 226.495 66.610 226.875 ;
        RECT 92.705 225.775 94.455 242.280 ;
        RECT 97.415 241.610 97.795 241.990 ;
        RECT 99.455 241.610 99.835 241.990 ;
        RECT 101.240 241.610 101.620 241.990 ;
        RECT 94.970 239.705 95.350 240.085 ;
        RECT 97.415 238.610 97.795 238.990 ;
        RECT 99.455 238.610 99.835 238.990 ;
        RECT 101.240 238.610 101.620 238.990 ;
        RECT 94.970 237.865 95.350 238.245 ;
        RECT 94.970 236.020 95.350 236.400 ;
        RECT 97.415 235.610 97.795 235.990 ;
        RECT 99.455 235.610 99.835 235.990 ;
        RECT 101.240 235.610 101.620 235.990 ;
        RECT 94.970 233.380 95.350 233.760 ;
        RECT 97.415 232.610 97.795 232.990 ;
        RECT 99.455 232.610 99.835 232.990 ;
        RECT 101.240 232.610 101.620 232.990 ;
        RECT 94.970 231.540 95.350 231.920 ;
        RECT 94.970 229.695 95.350 230.075 ;
        RECT 97.415 229.610 97.795 229.990 ;
        RECT 99.455 229.610 99.835 229.990 ;
        RECT 101.240 229.610 101.620 229.990 ;
        RECT 94.970 227.055 95.350 227.435 ;
        RECT 97.415 226.610 97.795 226.990 ;
        RECT 99.455 226.610 99.835 226.990 ;
        RECT 101.240 226.610 101.620 226.990 ;
        RECT 25.200 225.110 25.580 225.490 ;
        RECT 29.120 225.110 29.500 225.490 ;
        RECT 62.520 225.215 62.900 225.595 ;
        RECT 94.970 225.215 95.350 225.595 ;
        RECT 31.920 224.655 34.160 225.035 ;
        RECT 64.370 224.655 66.610 225.035 ;
        RECT 31.920 223.935 34.160 224.315 ;
        RECT 64.370 223.935 66.610 224.315 ;
        RECT 62.520 223.375 62.900 223.755 ;
        RECT 94.970 223.375 95.350 223.755 ;
        RECT 25.200 221.725 25.580 222.105 ;
        RECT 29.120 221.725 29.500 222.105 ;
        RECT 31.920 222.095 34.160 222.475 ;
        RECT 31.925 220.210 34.165 220.590 ;
        RECT 31.920 219.450 34.160 219.830 ;
        RECT 25.200 218.725 25.580 219.105 ;
        RECT 29.120 218.725 29.500 219.105 ;
        RECT 31.920 217.610 34.160 217.990 ;
        RECT 25.200 215.725 25.580 216.105 ;
        RECT 29.120 215.725 29.500 216.105 ;
        RECT 31.920 215.770 34.160 216.150 ;
        RECT 31.925 213.885 34.165 214.265 ;
        RECT 31.920 213.125 34.160 213.505 ;
        RECT 25.200 212.725 25.580 213.105 ;
        RECT 29.120 212.725 29.500 213.105 ;
        RECT 31.920 211.285 34.160 211.665 ;
        RECT 25.200 209.725 25.580 210.105 ;
        RECT 29.120 209.725 29.500 210.105 ;
        RECT 31.920 209.445 34.160 209.825 ;
        RECT 25.200 206.725 25.580 207.105 ;
        RECT 29.120 206.725 29.500 207.105 ;
        RECT 35.295 206.735 37.045 210.545 ;
        RECT 39.135 206.735 40.885 212.385 ;
        RECT 42.975 206.735 44.725 215.030 ;
        RECT 46.815 206.735 48.565 216.870 ;
        RECT 50.655 206.735 52.405 218.710 ;
        RECT 54.495 206.735 56.245 221.355 ;
        RECT 58.335 206.735 60.085 223.195 ;
        RECT 64.370 222.095 66.610 222.475 ;
        RECT 62.520 221.535 62.900 221.915 ;
        RECT 64.375 220.210 66.615 220.590 ;
        RECT 64.370 219.450 66.610 219.830 ;
        RECT 62.520 218.890 62.900 219.270 ;
        RECT 64.370 217.610 66.610 217.990 ;
        RECT 62.520 217.050 62.900 217.430 ;
        RECT 64.370 215.770 66.610 216.150 ;
        RECT 62.520 215.210 62.900 215.590 ;
        RECT 64.375 213.885 66.615 214.265 ;
        RECT 64.370 213.125 66.610 213.505 ;
        RECT 62.520 212.565 62.900 212.945 ;
        RECT 64.370 211.285 66.610 211.665 ;
        RECT 62.520 210.725 62.900 211.105 ;
        RECT 64.370 209.445 66.610 209.825 ;
        RECT 62.520 208.885 62.900 209.265 ;
        RECT 67.745 206.735 69.495 210.545 ;
        RECT 71.585 206.735 73.335 212.385 ;
        RECT 75.425 206.735 77.175 215.030 ;
        RECT 79.265 206.735 81.015 216.870 ;
        RECT 83.105 206.735 84.855 218.710 ;
        RECT 86.945 206.735 88.695 221.355 ;
        RECT 90.785 206.735 92.535 223.195 ;
        RECT 94.970 221.535 95.350 221.915 ;
        RECT 97.415 220.225 97.795 220.605 ;
        RECT 99.455 220.225 99.835 220.605 ;
        RECT 101.240 220.225 101.620 220.605 ;
        RECT 94.970 218.890 95.350 219.270 ;
        RECT 94.970 217.050 95.350 217.430 ;
        RECT 97.415 217.225 97.795 217.605 ;
        RECT 99.455 217.225 99.835 217.605 ;
        RECT 101.240 217.225 101.620 217.605 ;
        RECT 94.970 215.210 95.350 215.590 ;
        RECT 97.415 214.225 97.795 214.605 ;
        RECT 99.455 214.225 99.835 214.605 ;
        RECT 101.240 214.225 101.620 214.605 ;
        RECT 94.970 212.565 95.350 212.945 ;
        RECT 97.415 211.225 97.795 211.605 ;
        RECT 99.455 211.225 99.835 211.605 ;
        RECT 101.240 211.225 101.620 211.605 ;
        RECT 94.970 210.725 95.350 211.105 ;
        RECT 94.970 208.885 95.350 209.265 ;
        RECT 97.415 208.225 97.795 208.605 ;
        RECT 99.455 208.225 99.835 208.605 ;
        RECT 101.240 208.225 101.620 208.605 ;
        RECT 34.060 206.350 34.440 206.540 ;
        RECT 37.900 206.350 38.280 206.540 ;
        RECT 41.740 206.350 42.120 206.540 ;
        RECT 45.580 206.350 45.960 206.540 ;
        RECT 49.420 206.350 49.800 206.540 ;
        RECT 53.260 206.350 53.640 206.540 ;
        RECT 57.100 206.350 57.480 206.540 ;
        RECT 60.940 206.350 61.320 206.540 ;
        RECT 66.510 206.350 66.890 206.540 ;
        RECT 70.350 206.350 70.730 206.540 ;
        RECT 74.190 206.350 74.570 206.540 ;
        RECT 78.030 206.350 78.410 206.540 ;
        RECT 81.870 206.350 82.250 206.540 ;
        RECT 85.710 206.350 86.090 206.540 ;
        RECT 89.550 206.350 89.930 206.540 ;
        RECT 93.390 206.350 93.770 206.540 ;
        RECT 28.390 205.540 101.890 206.350 ;
        RECT 25.200 203.725 25.580 204.105 ;
        RECT 28.390 204.090 29.200 205.540 ;
        RECT 96.400 205.350 96.780 205.540 ;
        RECT 98.440 205.350 98.820 205.540 ;
        RECT 100.480 205.350 100.860 205.540 ;
        RECT 96.400 204.090 96.780 204.280 ;
        RECT 98.440 204.090 98.820 204.280 ;
        RECT 100.480 204.090 100.860 204.280 ;
        RECT 28.390 203.280 101.890 204.090 ;
        RECT 32.140 203.090 32.520 203.280 ;
        RECT 35.980 203.090 36.360 203.280 ;
        RECT 39.820 203.090 40.200 203.280 ;
        RECT 43.660 203.090 44.040 203.280 ;
        RECT 47.500 203.090 47.880 203.280 ;
        RECT 51.340 203.090 51.720 203.280 ;
        RECT 55.180 203.090 55.560 203.280 ;
        RECT 59.020 203.090 59.400 203.280 ;
        RECT 64.590 203.090 64.970 203.280 ;
        RECT 68.430 203.090 68.810 203.280 ;
        RECT 72.270 203.090 72.650 203.280 ;
        RECT 76.110 203.090 76.490 203.280 ;
        RECT 79.950 203.090 80.330 203.280 ;
        RECT 83.790 203.090 84.170 203.280 ;
        RECT 87.630 203.090 88.010 203.280 ;
        RECT 91.470 203.090 91.850 203.280 ;
        RECT 25.200 200.725 25.580 201.105 ;
        RECT 27.480 198.390 27.830 202.580 ;
        RECT 25.200 197.725 25.580 198.105 ;
        RECT 28.110 197.035 28.460 200.950 ;
        RECT 29.120 200.725 29.500 201.105 ;
        RECT 31.920 199.760 34.160 200.140 ;
        RECT 37.215 199.040 38.965 202.895 ;
        RECT 29.120 197.725 29.500 198.105 ;
        RECT 31.920 197.920 34.160 198.300 ;
        RECT 41.055 197.195 42.805 202.895 ;
        RECT 27.705 196.710 28.460 197.035 ;
        RECT 28.110 196.705 28.460 196.710 ;
        RECT 31.920 196.075 34.160 196.455 ;
        RECT 31.925 195.315 34.165 195.695 ;
        RECT 25.200 194.725 25.580 195.105 ;
        RECT 29.120 194.725 29.500 195.105 ;
        RECT 44.895 194.555 46.645 202.895 ;
        RECT 31.920 193.435 34.160 193.815 ;
        RECT 48.735 192.715 50.485 202.895 ;
        RECT 25.200 191.725 25.580 192.105 ;
        RECT 29.120 191.725 29.500 192.105 ;
        RECT 31.920 191.595 34.160 191.975 ;
        RECT 52.575 190.870 54.325 202.895 ;
        RECT 31.920 189.750 34.160 190.130 ;
        RECT 25.200 188.725 25.580 189.105 ;
        RECT 29.120 188.725 29.500 189.105 ;
        RECT 31.925 188.990 34.165 189.370 ;
        RECT 56.415 188.230 58.165 202.895 ;
        RECT 31.920 187.110 34.160 187.490 ;
        RECT 60.255 186.390 62.005 202.895 ;
        RECT 62.520 200.320 62.900 200.700 ;
        RECT 64.370 199.760 66.610 200.140 ;
        RECT 69.665 199.040 71.415 202.895 ;
        RECT 62.520 198.480 62.900 198.860 ;
        RECT 64.370 197.920 66.610 198.300 ;
        RECT 73.505 197.195 75.255 202.895 ;
        RECT 62.520 196.635 62.900 197.015 ;
        RECT 64.370 196.075 66.610 196.455 ;
        RECT 64.375 195.315 66.615 195.695 ;
        RECT 77.345 194.555 79.095 202.895 ;
        RECT 62.520 193.995 62.900 194.375 ;
        RECT 64.370 193.435 66.610 193.815 ;
        RECT 81.185 192.715 82.935 202.895 ;
        RECT 62.520 192.155 62.900 192.535 ;
        RECT 64.370 191.595 66.610 191.975 ;
        RECT 85.025 190.870 86.775 202.895 ;
        RECT 62.520 190.310 62.900 190.690 ;
        RECT 64.370 189.750 66.610 190.130 ;
        RECT 64.375 188.990 66.615 189.370 ;
        RECT 88.865 188.230 90.615 202.895 ;
        RECT 62.520 187.670 62.900 188.050 ;
        RECT 64.370 187.110 66.610 187.490 ;
        RECT 92.705 186.390 94.455 202.895 ;
        RECT 97.415 202.225 97.795 202.605 ;
        RECT 99.455 202.225 99.835 202.605 ;
        RECT 101.240 202.225 101.620 202.605 ;
        RECT 94.970 200.320 95.350 200.700 ;
        RECT 97.415 199.225 97.795 199.605 ;
        RECT 99.455 199.225 99.835 199.605 ;
        RECT 101.240 199.225 101.620 199.605 ;
        RECT 94.970 198.480 95.350 198.860 ;
        RECT 94.970 196.635 95.350 197.015 ;
        RECT 97.415 196.225 97.795 196.605 ;
        RECT 99.455 196.225 99.835 196.605 ;
        RECT 101.240 196.225 101.620 196.605 ;
        RECT 94.970 193.995 95.350 194.375 ;
        RECT 97.415 193.225 97.795 193.605 ;
        RECT 99.455 193.225 99.835 193.605 ;
        RECT 101.240 193.225 101.620 193.605 ;
        RECT 94.970 192.155 95.350 192.535 ;
        RECT 94.970 190.310 95.350 190.690 ;
        RECT 97.415 190.225 97.795 190.605 ;
        RECT 99.455 190.225 99.835 190.605 ;
        RECT 101.240 190.225 101.620 190.605 ;
        RECT 94.970 187.670 95.350 188.050 ;
        RECT 97.415 187.225 97.795 187.605 ;
        RECT 99.455 187.225 99.835 187.605 ;
        RECT 101.240 187.225 101.620 187.605 ;
        RECT 25.200 185.725 25.580 186.105 ;
        RECT 29.120 185.725 29.500 186.105 ;
        RECT 62.520 185.830 62.900 186.210 ;
        RECT 94.970 185.830 95.350 186.210 ;
        RECT 31.920 185.270 34.160 185.650 ;
        RECT 64.370 185.270 66.610 185.650 ;
        RECT 31.920 184.550 34.160 184.930 ;
        RECT 64.370 184.550 66.610 184.930 ;
        RECT 62.520 183.990 62.900 184.370 ;
        RECT 94.970 183.990 95.350 184.370 ;
        RECT 25.200 182.340 25.580 182.720 ;
        RECT 29.120 182.340 29.500 182.720 ;
        RECT 31.920 182.710 34.160 183.090 ;
        RECT 31.925 180.825 34.165 181.205 ;
        RECT 31.920 180.065 34.160 180.445 ;
        RECT 25.200 179.340 25.580 179.720 ;
        RECT 29.120 179.340 29.500 179.720 ;
        RECT 31.920 178.225 34.160 178.605 ;
        RECT 25.200 176.340 25.580 176.720 ;
        RECT 29.120 176.340 29.500 176.720 ;
        RECT 31.920 176.385 34.160 176.765 ;
        RECT 31.925 174.500 34.165 174.880 ;
        RECT 31.920 173.740 34.160 174.120 ;
        RECT 25.200 173.340 25.580 173.720 ;
        RECT 29.120 173.340 29.500 173.720 ;
        RECT 31.920 171.900 34.160 172.280 ;
        RECT 25.200 170.340 25.580 170.720 ;
        RECT 29.120 170.340 29.500 170.720 ;
        RECT 31.920 170.060 34.160 170.440 ;
        RECT 25.200 167.340 25.580 167.720 ;
        RECT 29.120 167.340 29.500 167.720 ;
        RECT 35.295 167.350 37.045 171.160 ;
        RECT 39.135 167.350 40.885 173.000 ;
        RECT 42.975 167.350 44.725 175.645 ;
        RECT 46.815 167.350 48.565 177.485 ;
        RECT 50.655 167.350 52.405 179.325 ;
        RECT 54.495 167.350 56.245 181.970 ;
        RECT 58.335 167.350 60.085 183.810 ;
        RECT 64.370 182.710 66.610 183.090 ;
        RECT 62.520 182.150 62.900 182.530 ;
        RECT 64.375 180.825 66.615 181.205 ;
        RECT 64.370 180.065 66.610 180.445 ;
        RECT 62.520 179.505 62.900 179.885 ;
        RECT 64.370 178.225 66.610 178.605 ;
        RECT 62.520 177.665 62.900 178.045 ;
        RECT 64.370 176.385 66.610 176.765 ;
        RECT 62.520 175.825 62.900 176.205 ;
        RECT 64.375 174.500 66.615 174.880 ;
        RECT 64.370 173.740 66.610 174.120 ;
        RECT 62.520 173.180 62.900 173.560 ;
        RECT 64.370 171.900 66.610 172.280 ;
        RECT 62.520 171.340 62.900 171.720 ;
        RECT 64.370 170.060 66.610 170.440 ;
        RECT 62.520 169.500 62.900 169.880 ;
        RECT 67.745 167.350 69.495 171.160 ;
        RECT 71.585 167.350 73.335 173.000 ;
        RECT 75.425 167.350 77.175 175.645 ;
        RECT 79.265 167.350 81.015 177.485 ;
        RECT 83.105 167.350 84.855 179.325 ;
        RECT 86.945 167.350 88.695 181.970 ;
        RECT 90.785 167.350 92.535 183.810 ;
        RECT 94.970 182.150 95.350 182.530 ;
        RECT 97.415 180.840 97.795 181.220 ;
        RECT 99.455 180.840 99.835 181.220 ;
        RECT 101.240 180.840 101.620 181.220 ;
        RECT 94.970 179.505 95.350 179.885 ;
        RECT 94.970 177.665 95.350 178.045 ;
        RECT 97.415 177.840 97.795 178.220 ;
        RECT 99.455 177.840 99.835 178.220 ;
        RECT 101.240 177.840 101.620 178.220 ;
        RECT 94.970 175.825 95.350 176.205 ;
        RECT 97.415 174.840 97.795 175.220 ;
        RECT 99.455 174.840 99.835 175.220 ;
        RECT 101.240 174.840 101.620 175.220 ;
        RECT 94.970 173.180 95.350 173.560 ;
        RECT 97.415 171.840 97.795 172.220 ;
        RECT 99.455 171.840 99.835 172.220 ;
        RECT 101.240 171.840 101.620 172.220 ;
        RECT 94.970 171.340 95.350 171.720 ;
        RECT 94.970 169.500 95.350 169.880 ;
        RECT 97.415 168.840 97.795 169.220 ;
        RECT 99.455 168.840 99.835 169.220 ;
        RECT 101.240 168.840 101.620 169.220 ;
        RECT 34.060 166.965 34.440 167.155 ;
        RECT 37.900 166.965 38.280 167.155 ;
        RECT 41.740 166.965 42.120 167.155 ;
        RECT 45.580 166.965 45.960 167.155 ;
        RECT 49.420 166.965 49.800 167.155 ;
        RECT 53.260 166.965 53.640 167.155 ;
        RECT 57.100 166.965 57.480 167.155 ;
        RECT 60.940 166.965 61.320 167.155 ;
        RECT 66.510 166.965 66.890 167.155 ;
        RECT 70.350 166.965 70.730 167.155 ;
        RECT 74.190 166.965 74.570 167.155 ;
        RECT 78.030 166.965 78.410 167.155 ;
        RECT 81.870 166.965 82.250 167.155 ;
        RECT 85.710 166.965 86.090 167.155 ;
        RECT 89.550 166.965 89.930 167.155 ;
        RECT 93.390 166.965 93.770 167.155 ;
        RECT 28.390 166.155 101.890 166.965 ;
        RECT 25.200 164.340 25.580 164.720 ;
        RECT 28.390 164.705 29.200 166.155 ;
        RECT 96.400 165.965 96.780 166.155 ;
        RECT 98.440 165.965 98.820 166.155 ;
        RECT 100.480 165.965 100.860 166.155 ;
        RECT 96.400 164.705 96.780 164.895 ;
        RECT 98.440 164.705 98.820 164.895 ;
        RECT 100.480 164.705 100.860 164.895 ;
        RECT 28.390 163.895 101.890 164.705 ;
        RECT 32.140 163.705 32.520 163.895 ;
        RECT 35.980 163.705 36.360 163.895 ;
        RECT 39.820 163.705 40.200 163.895 ;
        RECT 43.660 163.705 44.040 163.895 ;
        RECT 47.500 163.705 47.880 163.895 ;
        RECT 51.340 163.705 51.720 163.895 ;
        RECT 55.180 163.705 55.560 163.895 ;
        RECT 59.020 163.705 59.400 163.895 ;
        RECT 64.590 163.705 64.970 163.895 ;
        RECT 68.430 163.705 68.810 163.895 ;
        RECT 72.270 163.705 72.650 163.895 ;
        RECT 76.110 163.705 76.490 163.895 ;
        RECT 79.950 163.705 80.330 163.895 ;
        RECT 83.790 163.705 84.170 163.895 ;
        RECT 87.630 163.705 88.010 163.895 ;
        RECT 91.470 163.705 91.850 163.895 ;
        RECT 25.200 161.340 25.580 161.720 ;
        RECT 27.480 159.005 27.830 163.195 ;
        RECT 25.200 158.340 25.580 158.720 ;
        RECT 28.110 157.650 28.460 161.565 ;
        RECT 29.120 161.340 29.500 161.720 ;
        RECT 31.920 160.375 34.160 160.755 ;
        RECT 37.215 159.655 38.965 163.510 ;
        RECT 29.120 158.340 29.500 158.720 ;
        RECT 31.920 158.535 34.160 158.915 ;
        RECT 41.055 157.810 42.805 163.510 ;
        RECT 27.705 157.325 28.460 157.650 ;
        RECT 28.110 157.320 28.460 157.325 ;
        RECT 31.920 156.690 34.160 157.070 ;
        RECT 31.925 155.930 34.165 156.310 ;
        RECT 25.200 155.340 25.580 155.720 ;
        RECT 29.120 155.340 29.500 155.720 ;
        RECT 44.895 155.170 46.645 163.510 ;
        RECT 31.920 154.050 34.160 154.430 ;
        RECT 48.735 153.330 50.485 163.510 ;
        RECT 25.200 152.340 25.580 152.720 ;
        RECT 29.120 152.340 29.500 152.720 ;
        RECT 31.920 152.210 34.160 152.590 ;
        RECT 52.575 151.485 54.325 163.510 ;
        RECT 31.920 150.365 34.160 150.745 ;
        RECT 25.200 149.340 25.580 149.720 ;
        RECT 29.120 149.340 29.500 149.720 ;
        RECT 31.925 149.605 34.165 149.985 ;
        RECT 56.415 148.845 58.165 163.510 ;
        RECT 31.920 147.725 34.160 148.105 ;
        RECT 60.255 147.005 62.005 163.510 ;
        RECT 62.520 160.935 62.900 161.315 ;
        RECT 64.370 160.375 66.610 160.755 ;
        RECT 69.665 159.655 71.415 163.510 ;
        RECT 62.520 159.095 62.900 159.475 ;
        RECT 64.370 158.535 66.610 158.915 ;
        RECT 73.505 157.810 75.255 163.510 ;
        RECT 62.520 157.250 62.900 157.630 ;
        RECT 64.370 156.690 66.610 157.070 ;
        RECT 64.375 155.930 66.615 156.310 ;
        RECT 77.345 155.170 79.095 163.510 ;
        RECT 62.520 154.610 62.900 154.990 ;
        RECT 64.370 154.050 66.610 154.430 ;
        RECT 81.185 153.330 82.935 163.510 ;
        RECT 62.520 152.770 62.900 153.150 ;
        RECT 64.370 152.210 66.610 152.590 ;
        RECT 85.025 151.485 86.775 163.510 ;
        RECT 62.520 150.925 62.900 151.305 ;
        RECT 64.370 150.365 66.610 150.745 ;
        RECT 64.375 149.605 66.615 149.985 ;
        RECT 88.865 148.845 90.615 163.510 ;
        RECT 62.520 148.285 62.900 148.665 ;
        RECT 64.370 147.725 66.610 148.105 ;
        RECT 92.705 147.005 94.455 163.510 ;
        RECT 97.415 162.840 97.795 163.220 ;
        RECT 99.455 162.840 99.835 163.220 ;
        RECT 101.240 162.840 101.620 163.220 ;
        RECT 94.970 160.935 95.350 161.315 ;
        RECT 97.415 159.840 97.795 160.220 ;
        RECT 99.455 159.840 99.835 160.220 ;
        RECT 101.240 159.840 101.620 160.220 ;
        RECT 94.970 159.095 95.350 159.475 ;
        RECT 94.970 157.250 95.350 157.630 ;
        RECT 97.415 156.840 97.795 157.220 ;
        RECT 99.455 156.840 99.835 157.220 ;
        RECT 101.240 156.840 101.620 157.220 ;
        RECT 94.970 154.610 95.350 154.990 ;
        RECT 97.415 153.840 97.795 154.220 ;
        RECT 99.455 153.840 99.835 154.220 ;
        RECT 101.240 153.840 101.620 154.220 ;
        RECT 94.970 152.770 95.350 153.150 ;
        RECT 94.970 150.925 95.350 151.305 ;
        RECT 97.415 150.840 97.795 151.220 ;
        RECT 99.455 150.840 99.835 151.220 ;
        RECT 101.240 150.840 101.620 151.220 ;
        RECT 94.970 148.285 95.350 148.665 ;
        RECT 97.415 147.840 97.795 148.220 ;
        RECT 99.455 147.840 99.835 148.220 ;
        RECT 101.240 147.840 101.620 148.220 ;
        RECT 25.200 146.340 25.580 146.720 ;
        RECT 29.120 146.340 29.500 146.720 ;
        RECT 62.520 146.445 62.900 146.825 ;
        RECT 94.970 146.445 95.350 146.825 ;
        RECT 31.920 145.885 34.160 146.265 ;
        RECT 64.370 145.885 66.610 146.265 ;
        RECT 31.920 145.165 34.160 145.545 ;
        RECT 64.370 145.165 66.610 145.545 ;
        RECT 62.520 144.605 62.900 144.985 ;
        RECT 94.970 144.605 95.350 144.985 ;
        RECT 25.200 142.955 25.580 143.335 ;
        RECT 29.120 142.955 29.500 143.335 ;
        RECT 31.920 143.325 34.160 143.705 ;
        RECT 31.925 141.440 34.165 141.820 ;
        RECT 31.920 140.680 34.160 141.060 ;
        RECT 25.200 139.955 25.580 140.335 ;
        RECT 29.120 139.955 29.500 140.335 ;
        RECT 31.920 138.840 34.160 139.220 ;
        RECT 25.200 136.955 25.580 137.335 ;
        RECT 29.120 136.955 29.500 137.335 ;
        RECT 31.920 137.000 34.160 137.380 ;
        RECT 31.925 135.115 34.165 135.495 ;
        RECT 31.920 134.355 34.160 134.735 ;
        RECT 25.200 133.955 25.580 134.335 ;
        RECT 29.120 133.955 29.500 134.335 ;
        RECT 31.920 132.515 34.160 132.895 ;
        RECT 25.200 130.955 25.580 131.335 ;
        RECT 29.120 130.955 29.500 131.335 ;
        RECT 31.920 130.675 34.160 131.055 ;
        RECT 25.200 127.955 25.580 128.335 ;
        RECT 29.120 127.955 29.500 128.335 ;
        RECT 35.295 127.965 37.045 131.775 ;
        RECT 39.135 127.965 40.885 133.615 ;
        RECT 42.975 127.965 44.725 136.260 ;
        RECT 46.815 127.965 48.565 138.100 ;
        RECT 50.655 127.965 52.405 139.940 ;
        RECT 54.495 127.965 56.245 142.585 ;
        RECT 58.335 127.965 60.085 144.425 ;
        RECT 64.370 143.325 66.610 143.705 ;
        RECT 62.520 142.765 62.900 143.145 ;
        RECT 64.375 141.440 66.615 141.820 ;
        RECT 64.370 140.680 66.610 141.060 ;
        RECT 62.520 140.120 62.900 140.500 ;
        RECT 64.370 138.840 66.610 139.220 ;
        RECT 62.520 138.280 62.900 138.660 ;
        RECT 64.370 137.000 66.610 137.380 ;
        RECT 62.520 136.440 62.900 136.820 ;
        RECT 64.375 135.115 66.615 135.495 ;
        RECT 64.370 134.355 66.610 134.735 ;
        RECT 62.520 133.795 62.900 134.175 ;
        RECT 64.370 132.515 66.610 132.895 ;
        RECT 62.520 131.955 62.900 132.335 ;
        RECT 64.370 130.675 66.610 131.055 ;
        RECT 62.520 130.115 62.900 130.495 ;
        RECT 67.745 127.965 69.495 131.775 ;
        RECT 71.585 127.965 73.335 133.615 ;
        RECT 75.425 127.965 77.175 136.260 ;
        RECT 79.265 127.965 81.015 138.100 ;
        RECT 83.105 127.965 84.855 139.940 ;
        RECT 86.945 127.965 88.695 142.585 ;
        RECT 90.785 127.965 92.535 144.425 ;
        RECT 94.970 142.765 95.350 143.145 ;
        RECT 97.415 141.455 97.795 141.835 ;
        RECT 99.455 141.455 99.835 141.835 ;
        RECT 101.240 141.455 101.620 141.835 ;
        RECT 94.970 140.120 95.350 140.500 ;
        RECT 94.970 138.280 95.350 138.660 ;
        RECT 97.415 138.455 97.795 138.835 ;
        RECT 99.455 138.455 99.835 138.835 ;
        RECT 101.240 138.455 101.620 138.835 ;
        RECT 94.970 136.440 95.350 136.820 ;
        RECT 97.415 135.455 97.795 135.835 ;
        RECT 99.455 135.455 99.835 135.835 ;
        RECT 101.240 135.455 101.620 135.835 ;
        RECT 94.970 133.795 95.350 134.175 ;
        RECT 97.415 132.455 97.795 132.835 ;
        RECT 99.455 132.455 99.835 132.835 ;
        RECT 101.240 132.455 101.620 132.835 ;
        RECT 94.970 131.955 95.350 132.335 ;
        RECT 94.970 130.115 95.350 130.495 ;
        RECT 97.415 129.455 97.795 129.835 ;
        RECT 99.455 129.455 99.835 129.835 ;
        RECT 101.240 129.455 101.620 129.835 ;
        RECT 34.060 127.580 34.440 127.770 ;
        RECT 37.900 127.580 38.280 127.770 ;
        RECT 41.740 127.580 42.120 127.770 ;
        RECT 45.580 127.580 45.960 127.770 ;
        RECT 49.420 127.580 49.800 127.770 ;
        RECT 53.260 127.580 53.640 127.770 ;
        RECT 57.100 127.580 57.480 127.770 ;
        RECT 60.940 127.580 61.320 127.770 ;
        RECT 66.510 127.580 66.890 127.770 ;
        RECT 70.350 127.580 70.730 127.770 ;
        RECT 74.190 127.580 74.570 127.770 ;
        RECT 78.030 127.580 78.410 127.770 ;
        RECT 81.870 127.580 82.250 127.770 ;
        RECT 85.710 127.580 86.090 127.770 ;
        RECT 89.550 127.580 89.930 127.770 ;
        RECT 93.390 127.580 93.770 127.770 ;
        RECT 28.390 126.770 101.890 127.580 ;
        RECT 25.200 124.955 25.580 125.335 ;
        RECT 28.390 125.320 29.200 126.770 ;
        RECT 96.400 126.580 96.780 126.770 ;
        RECT 98.440 126.580 98.820 126.770 ;
        RECT 100.480 126.580 100.860 126.770 ;
        RECT 96.400 125.320 96.780 125.510 ;
        RECT 98.440 125.320 98.820 125.510 ;
        RECT 100.480 125.320 100.860 125.510 ;
        RECT 28.390 124.510 101.890 125.320 ;
        RECT 32.140 124.320 32.520 124.510 ;
        RECT 35.980 124.320 36.360 124.510 ;
        RECT 39.820 124.320 40.200 124.510 ;
        RECT 43.660 124.320 44.040 124.510 ;
        RECT 47.500 124.320 47.880 124.510 ;
        RECT 51.340 124.320 51.720 124.510 ;
        RECT 55.180 124.320 55.560 124.510 ;
        RECT 59.020 124.320 59.400 124.510 ;
        RECT 64.590 124.320 64.970 124.510 ;
        RECT 68.430 124.320 68.810 124.510 ;
        RECT 72.270 124.320 72.650 124.510 ;
        RECT 76.110 124.320 76.490 124.510 ;
        RECT 79.950 124.320 80.330 124.510 ;
        RECT 83.790 124.320 84.170 124.510 ;
        RECT 87.630 124.320 88.010 124.510 ;
        RECT 91.470 124.320 91.850 124.510 ;
        RECT 25.200 121.955 25.580 122.335 ;
        RECT 27.480 119.620 27.830 123.810 ;
        RECT 25.200 118.955 25.580 119.335 ;
        RECT 28.110 118.265 28.460 122.180 ;
        RECT 29.120 121.955 29.500 122.335 ;
        RECT 31.920 120.990 34.160 121.370 ;
        RECT 37.215 120.270 38.965 124.125 ;
        RECT 29.120 118.955 29.500 119.335 ;
        RECT 31.920 119.150 34.160 119.530 ;
        RECT 41.055 118.425 42.805 124.125 ;
        RECT 27.705 117.940 28.460 118.265 ;
        RECT 28.110 117.935 28.460 117.940 ;
        RECT 31.920 117.305 34.160 117.685 ;
        RECT 31.925 116.545 34.165 116.925 ;
        RECT 25.200 115.955 25.580 116.335 ;
        RECT 29.120 115.955 29.500 116.335 ;
        RECT 44.895 115.785 46.645 124.125 ;
        RECT 31.920 114.665 34.160 115.045 ;
        RECT 48.735 113.945 50.485 124.125 ;
        RECT 25.200 112.955 25.580 113.335 ;
        RECT 29.120 112.955 29.500 113.335 ;
        RECT 31.920 112.825 34.160 113.205 ;
        RECT 52.575 112.100 54.325 124.125 ;
        RECT 31.920 110.980 34.160 111.360 ;
        RECT 25.200 109.955 25.580 110.335 ;
        RECT 29.120 109.955 29.500 110.335 ;
        RECT 31.925 110.220 34.165 110.600 ;
        RECT 56.415 109.460 58.165 124.125 ;
        RECT 31.920 108.340 34.160 108.720 ;
        RECT 60.255 107.620 62.005 124.125 ;
        RECT 62.520 121.550 62.900 121.930 ;
        RECT 64.370 120.990 66.610 121.370 ;
        RECT 69.665 120.270 71.415 124.125 ;
        RECT 62.520 119.710 62.900 120.090 ;
        RECT 64.370 119.150 66.610 119.530 ;
        RECT 73.505 118.425 75.255 124.125 ;
        RECT 62.520 117.865 62.900 118.245 ;
        RECT 64.370 117.305 66.610 117.685 ;
        RECT 64.375 116.545 66.615 116.925 ;
        RECT 77.345 115.785 79.095 124.125 ;
        RECT 62.520 115.225 62.900 115.605 ;
        RECT 64.370 114.665 66.610 115.045 ;
        RECT 81.185 113.945 82.935 124.125 ;
        RECT 62.520 113.385 62.900 113.765 ;
        RECT 64.370 112.825 66.610 113.205 ;
        RECT 85.025 112.100 86.775 124.125 ;
        RECT 62.520 111.540 62.900 111.920 ;
        RECT 64.370 110.980 66.610 111.360 ;
        RECT 64.375 110.220 66.615 110.600 ;
        RECT 88.865 109.460 90.615 124.125 ;
        RECT 62.520 108.900 62.900 109.280 ;
        RECT 64.370 108.340 66.610 108.720 ;
        RECT 92.705 107.620 94.455 124.125 ;
        RECT 97.415 123.455 97.795 123.835 ;
        RECT 99.455 123.455 99.835 123.835 ;
        RECT 101.240 123.455 101.620 123.835 ;
        RECT 94.970 121.550 95.350 121.930 ;
        RECT 97.415 120.455 97.795 120.835 ;
        RECT 99.455 120.455 99.835 120.835 ;
        RECT 101.240 120.455 101.620 120.835 ;
        RECT 94.970 119.710 95.350 120.090 ;
        RECT 94.970 117.865 95.350 118.245 ;
        RECT 97.415 117.455 97.795 117.835 ;
        RECT 99.455 117.455 99.835 117.835 ;
        RECT 101.240 117.455 101.620 117.835 ;
        RECT 94.970 115.225 95.350 115.605 ;
        RECT 97.415 114.455 97.795 114.835 ;
        RECT 99.455 114.455 99.835 114.835 ;
        RECT 101.240 114.455 101.620 114.835 ;
        RECT 94.970 113.385 95.350 113.765 ;
        RECT 94.970 111.540 95.350 111.920 ;
        RECT 97.415 111.455 97.795 111.835 ;
        RECT 99.455 111.455 99.835 111.835 ;
        RECT 101.240 111.455 101.620 111.835 ;
        RECT 94.970 108.900 95.350 109.280 ;
        RECT 97.415 108.455 97.795 108.835 ;
        RECT 99.455 108.455 99.835 108.835 ;
        RECT 101.240 108.455 101.620 108.835 ;
        RECT 25.200 106.955 25.580 107.335 ;
        RECT 29.120 106.955 29.500 107.335 ;
        RECT 62.520 107.060 62.900 107.440 ;
        RECT 94.970 107.060 95.350 107.440 ;
        RECT 31.920 106.500 34.160 106.880 ;
        RECT 64.370 106.500 66.610 106.880 ;
        RECT 31.920 105.780 34.160 106.160 ;
        RECT 64.370 105.780 66.610 106.160 ;
        RECT 62.520 105.220 62.900 105.600 ;
        RECT 94.970 105.220 95.350 105.600 ;
        RECT 25.200 103.570 25.580 103.950 ;
        RECT 29.120 103.570 29.500 103.950 ;
        RECT 31.920 103.940 34.160 104.320 ;
        RECT 31.925 102.055 34.165 102.435 ;
        RECT 31.920 101.295 34.160 101.675 ;
        RECT 25.200 100.570 25.580 100.950 ;
        RECT 29.120 100.570 29.500 100.950 ;
        RECT 31.920 99.455 34.160 99.835 ;
        RECT 25.200 97.570 25.580 97.950 ;
        RECT 29.120 97.570 29.500 97.950 ;
        RECT 31.920 97.615 34.160 97.995 ;
        RECT 31.925 95.730 34.165 96.110 ;
        RECT 31.920 94.970 34.160 95.350 ;
        RECT 25.200 94.570 25.580 94.950 ;
        RECT 29.120 94.570 29.500 94.950 ;
        RECT 31.920 93.130 34.160 93.510 ;
        RECT 25.200 91.570 25.580 91.950 ;
        RECT 29.120 91.570 29.500 91.950 ;
        RECT 31.920 91.290 34.160 91.670 ;
        RECT 25.200 88.570 25.580 88.950 ;
        RECT 29.120 88.570 29.500 88.950 ;
        RECT 35.295 88.580 37.045 92.390 ;
        RECT 39.135 88.580 40.885 94.230 ;
        RECT 42.975 88.580 44.725 96.875 ;
        RECT 46.815 88.580 48.565 98.715 ;
        RECT 50.655 88.580 52.405 100.555 ;
        RECT 54.495 88.580 56.245 103.200 ;
        RECT 58.335 88.580 60.085 105.040 ;
        RECT 64.370 103.940 66.610 104.320 ;
        RECT 62.520 103.380 62.900 103.760 ;
        RECT 64.375 102.055 66.615 102.435 ;
        RECT 64.370 101.295 66.610 101.675 ;
        RECT 62.520 100.735 62.900 101.115 ;
        RECT 64.370 99.455 66.610 99.835 ;
        RECT 62.520 98.895 62.900 99.275 ;
        RECT 64.370 97.615 66.610 97.995 ;
        RECT 62.520 97.055 62.900 97.435 ;
        RECT 64.375 95.730 66.615 96.110 ;
        RECT 64.370 94.970 66.610 95.350 ;
        RECT 62.520 94.410 62.900 94.790 ;
        RECT 64.370 93.130 66.610 93.510 ;
        RECT 62.520 92.570 62.900 92.950 ;
        RECT 64.370 91.290 66.610 91.670 ;
        RECT 62.520 90.730 62.900 91.110 ;
        RECT 67.745 88.580 69.495 92.390 ;
        RECT 71.585 88.580 73.335 94.230 ;
        RECT 75.425 88.580 77.175 96.875 ;
        RECT 79.265 88.580 81.015 98.715 ;
        RECT 83.105 88.580 84.855 100.555 ;
        RECT 86.945 88.580 88.695 103.200 ;
        RECT 90.785 88.580 92.535 105.040 ;
        RECT 94.970 103.380 95.350 103.760 ;
        RECT 97.415 102.070 97.795 102.450 ;
        RECT 99.455 102.070 99.835 102.450 ;
        RECT 101.240 102.070 101.620 102.450 ;
        RECT 94.970 100.735 95.350 101.115 ;
        RECT 94.970 98.895 95.350 99.275 ;
        RECT 97.415 99.070 97.795 99.450 ;
        RECT 99.455 99.070 99.835 99.450 ;
        RECT 101.240 99.070 101.620 99.450 ;
        RECT 94.970 97.055 95.350 97.435 ;
        RECT 97.415 96.070 97.795 96.450 ;
        RECT 99.455 96.070 99.835 96.450 ;
        RECT 101.240 96.070 101.620 96.450 ;
        RECT 94.970 94.410 95.350 94.790 ;
        RECT 97.415 93.070 97.795 93.450 ;
        RECT 99.455 93.070 99.835 93.450 ;
        RECT 101.240 93.070 101.620 93.450 ;
        RECT 94.970 92.570 95.350 92.950 ;
        RECT 94.970 90.730 95.350 91.110 ;
        RECT 97.415 90.070 97.795 90.450 ;
        RECT 99.455 90.070 99.835 90.450 ;
        RECT 101.240 90.070 101.620 90.450 ;
        RECT 34.060 88.195 34.440 88.385 ;
        RECT 37.900 88.195 38.280 88.385 ;
        RECT 41.740 88.195 42.120 88.385 ;
        RECT 45.580 88.195 45.960 88.385 ;
        RECT 49.420 88.195 49.800 88.385 ;
        RECT 53.260 88.195 53.640 88.385 ;
        RECT 57.100 88.195 57.480 88.385 ;
        RECT 60.940 88.195 61.320 88.385 ;
        RECT 66.510 88.195 66.890 88.385 ;
        RECT 70.350 88.195 70.730 88.385 ;
        RECT 74.190 88.195 74.570 88.385 ;
        RECT 78.030 88.195 78.410 88.385 ;
        RECT 81.870 88.195 82.250 88.385 ;
        RECT 85.710 88.195 86.090 88.385 ;
        RECT 89.550 88.195 89.930 88.385 ;
        RECT 93.390 88.195 93.770 88.385 ;
        RECT 28.390 87.385 101.890 88.195 ;
        RECT 25.200 85.570 25.580 85.950 ;
        RECT 28.390 85.935 29.200 87.385 ;
        RECT 96.400 87.195 96.780 87.385 ;
        RECT 98.440 87.195 98.820 87.385 ;
        RECT 100.480 87.195 100.860 87.385 ;
        RECT 96.400 85.935 96.780 86.125 ;
        RECT 98.440 85.935 98.820 86.125 ;
        RECT 100.480 85.935 100.860 86.125 ;
        RECT 28.390 85.125 101.890 85.935 ;
        RECT 32.140 84.935 32.520 85.125 ;
        RECT 35.980 84.935 36.360 85.125 ;
        RECT 39.820 84.935 40.200 85.125 ;
        RECT 43.660 84.935 44.040 85.125 ;
        RECT 47.500 84.935 47.880 85.125 ;
        RECT 51.340 84.935 51.720 85.125 ;
        RECT 55.180 84.935 55.560 85.125 ;
        RECT 59.020 84.935 59.400 85.125 ;
        RECT 64.590 84.935 64.970 85.125 ;
        RECT 68.430 84.935 68.810 85.125 ;
        RECT 72.270 84.935 72.650 85.125 ;
        RECT 76.110 84.935 76.490 85.125 ;
        RECT 79.950 84.935 80.330 85.125 ;
        RECT 83.790 84.935 84.170 85.125 ;
        RECT 87.630 84.935 88.010 85.125 ;
        RECT 91.470 84.935 91.850 85.125 ;
        RECT 25.200 82.570 25.580 82.950 ;
        RECT 27.480 80.235 27.830 84.425 ;
        RECT 25.200 79.570 25.580 79.950 ;
        RECT 28.110 78.880 28.460 82.795 ;
        RECT 29.120 82.570 29.500 82.950 ;
        RECT 31.920 81.605 34.160 81.985 ;
        RECT 37.215 80.885 38.965 84.740 ;
        RECT 29.120 79.570 29.500 79.950 ;
        RECT 31.920 79.765 34.160 80.145 ;
        RECT 41.055 79.040 42.805 84.740 ;
        RECT 27.705 78.555 28.460 78.880 ;
        RECT 28.110 78.550 28.460 78.555 ;
        RECT 31.920 77.920 34.160 78.300 ;
        RECT 31.925 77.160 34.165 77.540 ;
        RECT 25.200 76.570 25.580 76.950 ;
        RECT 29.120 76.570 29.500 76.950 ;
        RECT 44.895 76.400 46.645 84.740 ;
        RECT 31.920 75.280 34.160 75.660 ;
        RECT 48.735 74.560 50.485 84.740 ;
        RECT 25.200 73.570 25.580 73.950 ;
        RECT 29.120 73.570 29.500 73.950 ;
        RECT 31.920 73.440 34.160 73.820 ;
        RECT 52.575 72.715 54.325 84.740 ;
        RECT 31.920 71.595 34.160 71.975 ;
        RECT 25.200 70.570 25.580 70.950 ;
        RECT 29.120 70.570 29.500 70.950 ;
        RECT 31.925 70.835 34.165 71.215 ;
        RECT 56.415 70.075 58.165 84.740 ;
        RECT 31.920 68.955 34.160 69.335 ;
        RECT 60.255 68.235 62.005 84.740 ;
        RECT 62.520 82.165 62.900 82.545 ;
        RECT 64.370 81.605 66.610 81.985 ;
        RECT 69.665 80.885 71.415 84.740 ;
        RECT 62.520 80.325 62.900 80.705 ;
        RECT 64.370 79.765 66.610 80.145 ;
        RECT 73.505 79.040 75.255 84.740 ;
        RECT 62.520 78.480 62.900 78.860 ;
        RECT 64.370 77.920 66.610 78.300 ;
        RECT 64.375 77.160 66.615 77.540 ;
        RECT 77.345 76.400 79.095 84.740 ;
        RECT 62.520 75.840 62.900 76.220 ;
        RECT 64.370 75.280 66.610 75.660 ;
        RECT 81.185 74.560 82.935 84.740 ;
        RECT 62.520 74.000 62.900 74.380 ;
        RECT 64.370 73.440 66.610 73.820 ;
        RECT 85.025 72.715 86.775 84.740 ;
        RECT 62.520 72.155 62.900 72.535 ;
        RECT 64.370 71.595 66.610 71.975 ;
        RECT 64.375 70.835 66.615 71.215 ;
        RECT 88.865 70.075 90.615 84.740 ;
        RECT 62.520 69.515 62.900 69.895 ;
        RECT 64.370 68.955 66.610 69.335 ;
        RECT 92.705 68.235 94.455 84.740 ;
        RECT 97.415 84.070 97.795 84.450 ;
        RECT 99.455 84.070 99.835 84.450 ;
        RECT 101.240 84.070 101.620 84.450 ;
        RECT 94.970 82.165 95.350 82.545 ;
        RECT 97.415 81.070 97.795 81.450 ;
        RECT 99.455 81.070 99.835 81.450 ;
        RECT 101.240 81.070 101.620 81.450 ;
        RECT 94.970 80.325 95.350 80.705 ;
        RECT 94.970 78.480 95.350 78.860 ;
        RECT 97.415 78.070 97.795 78.450 ;
        RECT 99.455 78.070 99.835 78.450 ;
        RECT 101.240 78.070 101.620 78.450 ;
        RECT 94.970 75.840 95.350 76.220 ;
        RECT 97.415 75.070 97.795 75.450 ;
        RECT 99.455 75.070 99.835 75.450 ;
        RECT 101.240 75.070 101.620 75.450 ;
        RECT 94.970 74.000 95.350 74.380 ;
        RECT 94.970 72.155 95.350 72.535 ;
        RECT 97.415 72.070 97.795 72.450 ;
        RECT 99.455 72.070 99.835 72.450 ;
        RECT 101.240 72.070 101.620 72.450 ;
        RECT 94.970 69.515 95.350 69.895 ;
        RECT 97.415 69.070 97.795 69.450 ;
        RECT 99.455 69.070 99.835 69.450 ;
        RECT 101.240 69.070 101.620 69.450 ;
        RECT 25.200 67.570 25.580 67.950 ;
        RECT 29.120 67.570 29.500 67.950 ;
        RECT 62.520 67.675 62.900 68.055 ;
        RECT 94.970 67.675 95.350 68.055 ;
        RECT 31.920 67.115 34.160 67.495 ;
        RECT 64.370 67.115 66.610 67.495 ;
      LAYER Metal3 ;
        RECT 31.920 381.475 34.160 381.855 ;
        RECT 64.370 381.475 66.610 381.855 ;
        RECT 53.700 381.245 54.080 381.295 ;
        RECT 62.520 381.245 62.900 381.295 ;
        RECT 53.700 380.965 62.900 381.245 ;
        RECT 53.700 380.915 54.080 380.965 ;
        RECT 62.520 380.915 62.900 380.965 ;
        RECT 86.150 381.245 86.530 381.295 ;
        RECT 94.970 381.245 95.350 381.295 ;
        RECT 86.150 380.965 95.350 381.245 ;
        RECT 86.150 380.915 86.530 380.965 ;
        RECT 94.970 380.915 95.350 380.965 ;
        RECT 25.200 379.265 25.580 379.645 ;
        RECT 29.120 379.265 29.500 379.645 ;
        RECT 31.920 379.635 34.160 380.015 ;
        RECT 64.370 379.635 66.610 380.015 ;
        RECT 54.980 379.405 55.360 379.455 ;
        RECT 62.520 379.405 62.900 379.455 ;
        RECT 54.980 379.125 62.900 379.405 ;
        RECT 54.980 379.075 55.360 379.125 ;
        RECT 62.520 379.075 62.900 379.125 ;
        RECT 87.430 379.405 87.810 379.455 ;
        RECT 94.970 379.405 95.350 379.455 ;
        RECT 87.430 379.125 95.350 379.405 ;
        RECT 87.430 379.075 87.810 379.125 ;
        RECT 94.970 379.075 95.350 379.125 ;
        RECT 31.925 377.750 34.165 378.130 ;
        RECT 64.375 377.750 66.615 378.130 ;
        RECT 97.415 377.765 97.795 378.145 ;
        RECT 99.455 377.765 99.835 378.145 ;
        RECT 101.240 377.765 101.620 378.145 ;
        RECT 31.920 376.990 34.160 377.370 ;
        RECT 64.370 376.990 66.610 377.370 ;
        RECT 56.260 376.760 56.640 376.810 ;
        RECT 62.520 376.760 62.900 376.810 ;
        RECT 25.200 376.265 25.580 376.645 ;
        RECT 29.120 376.265 29.500 376.645 ;
        RECT 56.260 376.480 62.900 376.760 ;
        RECT 56.260 376.430 56.640 376.480 ;
        RECT 62.520 376.430 62.900 376.480 ;
        RECT 88.710 376.760 89.090 376.810 ;
        RECT 94.970 376.760 95.350 376.810 ;
        RECT 88.710 376.480 95.350 376.760 ;
        RECT 88.710 376.430 89.090 376.480 ;
        RECT 94.970 376.430 95.350 376.480 ;
        RECT 31.920 375.150 34.160 375.530 ;
        RECT 64.370 375.150 66.610 375.530 ;
        RECT 57.540 374.920 57.920 374.970 ;
        RECT 62.520 374.920 62.900 374.970 ;
        RECT 57.540 374.640 62.900 374.920 ;
        RECT 57.540 374.590 57.920 374.640 ;
        RECT 62.520 374.590 62.900 374.640 ;
        RECT 89.990 374.920 90.370 374.970 ;
        RECT 94.970 374.920 95.350 374.970 ;
        RECT 89.990 374.640 95.350 374.920 ;
        RECT 97.415 374.765 97.795 375.145 ;
        RECT 99.455 374.765 99.835 375.145 ;
        RECT 101.240 374.765 101.620 375.145 ;
        RECT 89.990 374.590 90.370 374.640 ;
        RECT 94.970 374.590 95.350 374.640 ;
        RECT 25.200 373.265 25.580 373.645 ;
        RECT 29.120 373.265 29.500 373.645 ;
        RECT 31.920 373.310 34.160 373.690 ;
        RECT 64.370 373.310 66.610 373.690 ;
        RECT 58.820 373.080 59.200 373.130 ;
        RECT 62.520 373.080 62.900 373.130 ;
        RECT 58.820 372.800 62.900 373.080 ;
        RECT 58.820 372.750 59.200 372.800 ;
        RECT 62.520 372.750 62.900 372.800 ;
        RECT 91.270 373.080 91.650 373.130 ;
        RECT 94.970 373.080 95.350 373.130 ;
        RECT 91.270 372.800 95.350 373.080 ;
        RECT 91.270 372.750 91.650 372.800 ;
        RECT 94.970 372.750 95.350 372.800 ;
        RECT 31.925 371.425 34.165 371.805 ;
        RECT 64.375 371.425 66.615 371.805 ;
        RECT 97.415 371.765 97.795 372.145 ;
        RECT 99.455 371.765 99.835 372.145 ;
        RECT 101.240 371.765 101.620 372.145 ;
        RECT 31.920 370.665 34.160 371.045 ;
        RECT 64.370 370.665 66.610 371.045 ;
        RECT 25.200 370.265 25.580 370.645 ;
        RECT 29.120 370.265 29.500 370.645 ;
        RECT 60.100 370.435 60.480 370.485 ;
        RECT 62.520 370.435 62.900 370.485 ;
        RECT 60.100 370.155 62.900 370.435 ;
        RECT 60.100 370.105 60.480 370.155 ;
        RECT 62.520 370.105 62.900 370.155 ;
        RECT 92.550 370.435 92.930 370.485 ;
        RECT 94.970 370.435 95.350 370.485 ;
        RECT 92.550 370.155 95.350 370.435 ;
        RECT 92.550 370.105 92.930 370.155 ;
        RECT 94.970 370.105 95.350 370.155 ;
        RECT 31.920 368.825 34.160 369.205 ;
        RECT 64.370 368.825 66.610 369.205 ;
        RECT 97.415 368.765 97.795 369.145 ;
        RECT 99.455 368.765 99.835 369.145 ;
        RECT 101.240 368.765 101.620 369.145 ;
        RECT 61.380 368.595 61.760 368.645 ;
        RECT 62.520 368.595 62.900 368.645 ;
        RECT 61.380 368.315 62.900 368.595 ;
        RECT 61.380 368.265 61.760 368.315 ;
        RECT 62.520 368.265 62.900 368.315 ;
        RECT 93.830 368.595 94.210 368.645 ;
        RECT 94.970 368.595 95.350 368.645 ;
        RECT 93.830 368.315 95.350 368.595 ;
        RECT 93.830 368.265 94.210 368.315 ;
        RECT 94.970 368.265 95.350 368.315 ;
        RECT 25.200 367.265 25.580 367.645 ;
        RECT 29.120 367.265 29.500 367.645 ;
        RECT 31.920 366.985 34.160 367.365 ;
        RECT 64.370 366.985 66.610 367.365 ;
        RECT 62.520 366.425 63.040 366.805 ;
        RECT 94.970 366.425 95.490 366.805 ;
        RECT 97.415 365.765 97.795 366.145 ;
        RECT 99.455 365.765 99.835 366.145 ;
        RECT 101.240 365.765 101.620 366.145 ;
        RECT 25.200 364.265 25.580 364.645 ;
        RECT 29.120 364.265 29.500 364.645 ;
        RECT 25.200 361.265 25.580 361.645 ;
        RECT 97.415 359.765 97.795 360.145 ;
        RECT 99.455 359.765 99.835 360.145 ;
        RECT 101.240 359.765 101.620 360.145 ;
        RECT 25.200 358.265 25.580 358.645 ;
        RECT 29.120 358.265 29.500 358.645 ;
        RECT 62.020 357.860 62.900 358.240 ;
        RECT 94.470 357.860 95.350 358.240 ;
        RECT 31.920 357.300 34.160 357.680 ;
        RECT 64.370 357.300 66.610 357.680 ;
        RECT 97.415 356.765 97.795 357.145 ;
        RECT 99.455 356.765 99.835 357.145 ;
        RECT 101.240 356.765 101.620 357.145 ;
        RECT 60.740 356.350 61.120 356.400 ;
        RECT 62.520 356.350 62.900 356.400 ;
        RECT 60.740 356.070 62.900 356.350 ;
        RECT 60.740 356.020 61.120 356.070 ;
        RECT 62.520 356.020 62.900 356.070 ;
        RECT 93.190 356.350 93.570 356.400 ;
        RECT 94.970 356.350 95.350 356.400 ;
        RECT 93.190 356.070 95.350 356.350 ;
        RECT 93.190 356.020 93.570 356.070 ;
        RECT 94.970 356.020 95.350 356.070 ;
        RECT 25.200 355.265 25.580 355.645 ;
        RECT 29.120 355.265 29.500 355.645 ;
        RECT 31.920 355.460 34.160 355.840 ;
        RECT 64.370 355.460 66.610 355.840 ;
        RECT 59.460 354.505 59.840 354.555 ;
        RECT 62.520 354.505 62.900 354.555 ;
        RECT 59.460 354.225 62.900 354.505 ;
        RECT 59.460 354.175 59.840 354.225 ;
        RECT 62.520 354.175 62.900 354.225 ;
        RECT 91.910 354.505 92.290 354.555 ;
        RECT 94.970 354.505 95.350 354.555 ;
        RECT 91.910 354.225 95.350 354.505 ;
        RECT 91.910 354.175 92.290 354.225 ;
        RECT 94.970 354.175 95.350 354.225 ;
        RECT 31.920 353.615 34.160 353.995 ;
        RECT 64.370 353.615 66.610 353.995 ;
        RECT 97.415 353.765 97.795 354.145 ;
        RECT 99.455 353.765 99.835 354.145 ;
        RECT 101.240 353.765 101.620 354.145 ;
        RECT 31.925 352.855 34.165 353.235 ;
        RECT 64.375 352.855 66.615 353.235 ;
        RECT 25.200 352.265 25.580 352.645 ;
        RECT 29.120 352.265 29.500 352.645 ;
        RECT 58.180 351.865 58.560 351.915 ;
        RECT 62.520 351.865 62.900 351.915 ;
        RECT 58.180 351.585 62.900 351.865 ;
        RECT 58.180 351.535 58.560 351.585 ;
        RECT 62.520 351.535 62.900 351.585 ;
        RECT 90.630 351.865 91.010 351.915 ;
        RECT 94.970 351.865 95.350 351.915 ;
        RECT 90.630 351.585 95.350 351.865 ;
        RECT 90.630 351.535 91.010 351.585 ;
        RECT 94.970 351.535 95.350 351.585 ;
        RECT 31.920 350.975 34.160 351.355 ;
        RECT 64.370 350.975 66.610 351.355 ;
        RECT 97.415 350.765 97.795 351.145 ;
        RECT 99.455 350.765 99.835 351.145 ;
        RECT 101.240 350.765 101.620 351.145 ;
        RECT 56.900 350.025 57.280 350.075 ;
        RECT 62.520 350.025 62.900 350.075 ;
        RECT 56.900 349.745 62.900 350.025 ;
        RECT 56.900 349.695 57.280 349.745 ;
        RECT 62.520 349.695 62.900 349.745 ;
        RECT 89.350 350.025 89.730 350.075 ;
        RECT 94.970 350.025 95.350 350.075 ;
        RECT 89.350 349.745 95.350 350.025 ;
        RECT 89.350 349.695 89.730 349.745 ;
        RECT 94.970 349.695 95.350 349.745 ;
        RECT 25.200 349.265 25.580 349.645 ;
        RECT 29.120 349.265 29.500 349.645 ;
        RECT 31.920 349.135 34.160 349.515 ;
        RECT 64.370 349.135 66.610 349.515 ;
        RECT 55.620 348.180 56.000 348.230 ;
        RECT 62.520 348.180 62.900 348.230 ;
        RECT 55.620 347.900 62.900 348.180 ;
        RECT 55.620 347.850 56.000 347.900 ;
        RECT 62.520 347.850 62.900 347.900 ;
        RECT 88.070 348.180 88.450 348.230 ;
        RECT 94.970 348.180 95.350 348.230 ;
        RECT 88.070 347.900 95.350 348.180 ;
        RECT 88.070 347.850 88.450 347.900 ;
        RECT 94.970 347.850 95.350 347.900 ;
        RECT 97.415 347.765 97.795 348.145 ;
        RECT 99.455 347.765 99.835 348.145 ;
        RECT 101.240 347.765 101.620 348.145 ;
        RECT 31.920 347.290 34.160 347.670 ;
        RECT 64.370 347.290 66.610 347.670 ;
        RECT 25.200 346.265 25.580 346.645 ;
        RECT 29.120 346.265 29.500 346.645 ;
        RECT 31.925 346.530 34.165 346.910 ;
        RECT 64.375 346.530 66.615 346.910 ;
        RECT 54.340 345.540 54.720 345.590 ;
        RECT 62.520 345.540 62.900 345.590 ;
        RECT 54.340 345.260 62.900 345.540 ;
        RECT 54.340 345.210 54.720 345.260 ;
        RECT 62.520 345.210 62.900 345.260 ;
        RECT 86.790 345.540 87.170 345.590 ;
        RECT 94.970 345.540 95.350 345.590 ;
        RECT 86.790 345.260 95.350 345.540 ;
        RECT 86.790 345.210 87.170 345.260 ;
        RECT 94.970 345.210 95.350 345.260 ;
        RECT 31.920 344.650 34.160 345.030 ;
        RECT 64.370 344.650 66.610 345.030 ;
        RECT 97.415 344.765 97.795 345.145 ;
        RECT 99.455 344.765 99.835 345.145 ;
        RECT 101.240 344.765 101.620 345.145 ;
        RECT 53.060 343.700 53.440 343.750 ;
        RECT 62.520 343.700 62.900 343.750 ;
        RECT 25.200 343.265 25.580 343.645 ;
        RECT 29.120 343.265 29.500 343.645 ;
        RECT 53.060 343.420 62.900 343.700 ;
        RECT 53.060 343.370 53.440 343.420 ;
        RECT 62.520 343.370 62.900 343.420 ;
        RECT 85.510 343.700 85.890 343.750 ;
        RECT 94.970 343.700 95.350 343.750 ;
        RECT 85.510 343.420 95.350 343.700 ;
        RECT 85.510 343.370 85.890 343.420 ;
        RECT 94.970 343.370 95.350 343.420 ;
        RECT 31.920 342.810 34.160 343.190 ;
        RECT 64.370 342.810 66.610 343.190 ;
        RECT 31.920 342.090 34.160 342.470 ;
        RECT 64.370 342.090 66.610 342.470 ;
        RECT 53.700 341.860 54.080 341.910 ;
        RECT 62.520 341.860 62.900 341.910 ;
        RECT 53.700 341.580 62.900 341.860 ;
        RECT 53.700 341.530 54.080 341.580 ;
        RECT 62.520 341.530 62.900 341.580 ;
        RECT 86.150 341.860 86.530 341.910 ;
        RECT 94.970 341.860 95.350 341.910 ;
        RECT 86.150 341.580 95.350 341.860 ;
        RECT 86.150 341.530 86.530 341.580 ;
        RECT 94.970 341.530 95.350 341.580 ;
        RECT 25.200 339.880 25.580 340.260 ;
        RECT 29.120 339.880 29.500 340.260 ;
        RECT 31.920 340.250 34.160 340.630 ;
        RECT 64.370 340.250 66.610 340.630 ;
        RECT 54.980 340.020 55.360 340.070 ;
        RECT 62.520 340.020 62.900 340.070 ;
        RECT 54.980 339.740 62.900 340.020 ;
        RECT 54.980 339.690 55.360 339.740 ;
        RECT 62.520 339.690 62.900 339.740 ;
        RECT 87.430 340.020 87.810 340.070 ;
        RECT 94.970 340.020 95.350 340.070 ;
        RECT 87.430 339.740 95.350 340.020 ;
        RECT 87.430 339.690 87.810 339.740 ;
        RECT 94.970 339.690 95.350 339.740 ;
        RECT 31.925 338.365 34.165 338.745 ;
        RECT 64.375 338.365 66.615 338.745 ;
        RECT 97.415 338.380 97.795 338.760 ;
        RECT 99.455 338.380 99.835 338.760 ;
        RECT 101.240 338.380 101.620 338.760 ;
        RECT 31.920 337.605 34.160 337.985 ;
        RECT 64.370 337.605 66.610 337.985 ;
        RECT 56.260 337.375 56.640 337.425 ;
        RECT 62.520 337.375 62.900 337.425 ;
        RECT 25.200 336.880 25.580 337.260 ;
        RECT 29.120 336.880 29.500 337.260 ;
        RECT 56.260 337.095 62.900 337.375 ;
        RECT 56.260 337.045 56.640 337.095 ;
        RECT 62.520 337.045 62.900 337.095 ;
        RECT 88.710 337.375 89.090 337.425 ;
        RECT 94.970 337.375 95.350 337.425 ;
        RECT 88.710 337.095 95.350 337.375 ;
        RECT 88.710 337.045 89.090 337.095 ;
        RECT 94.970 337.045 95.350 337.095 ;
        RECT 31.920 335.765 34.160 336.145 ;
        RECT 64.370 335.765 66.610 336.145 ;
        RECT 57.540 335.535 57.920 335.585 ;
        RECT 62.520 335.535 62.900 335.585 ;
        RECT 57.540 335.255 62.900 335.535 ;
        RECT 57.540 335.205 57.920 335.255 ;
        RECT 62.520 335.205 62.900 335.255 ;
        RECT 89.990 335.535 90.370 335.585 ;
        RECT 94.970 335.535 95.350 335.585 ;
        RECT 89.990 335.255 95.350 335.535 ;
        RECT 97.415 335.380 97.795 335.760 ;
        RECT 99.455 335.380 99.835 335.760 ;
        RECT 101.240 335.380 101.620 335.760 ;
        RECT 89.990 335.205 90.370 335.255 ;
        RECT 94.970 335.205 95.350 335.255 ;
        RECT 25.200 333.880 25.580 334.260 ;
        RECT 29.120 333.880 29.500 334.260 ;
        RECT 31.920 333.925 34.160 334.305 ;
        RECT 64.370 333.925 66.610 334.305 ;
        RECT 58.820 333.695 59.200 333.745 ;
        RECT 62.520 333.695 62.900 333.745 ;
        RECT 58.820 333.415 62.900 333.695 ;
        RECT 58.820 333.365 59.200 333.415 ;
        RECT 62.520 333.365 62.900 333.415 ;
        RECT 91.270 333.695 91.650 333.745 ;
        RECT 94.970 333.695 95.350 333.745 ;
        RECT 91.270 333.415 95.350 333.695 ;
        RECT 91.270 333.365 91.650 333.415 ;
        RECT 94.970 333.365 95.350 333.415 ;
        RECT 31.925 332.040 34.165 332.420 ;
        RECT 64.375 332.040 66.615 332.420 ;
        RECT 97.415 332.380 97.795 332.760 ;
        RECT 99.455 332.380 99.835 332.760 ;
        RECT 101.240 332.380 101.620 332.760 ;
        RECT 31.920 331.280 34.160 331.660 ;
        RECT 64.370 331.280 66.610 331.660 ;
        RECT 25.200 330.880 25.580 331.260 ;
        RECT 29.120 330.880 29.500 331.260 ;
        RECT 60.100 331.050 60.480 331.100 ;
        RECT 62.520 331.050 62.900 331.100 ;
        RECT 60.100 330.770 62.900 331.050 ;
        RECT 60.100 330.720 60.480 330.770 ;
        RECT 62.520 330.720 62.900 330.770 ;
        RECT 92.550 331.050 92.930 331.100 ;
        RECT 94.970 331.050 95.350 331.100 ;
        RECT 92.550 330.770 95.350 331.050 ;
        RECT 92.550 330.720 92.930 330.770 ;
        RECT 94.970 330.720 95.350 330.770 ;
        RECT 31.920 329.440 34.160 329.820 ;
        RECT 64.370 329.440 66.610 329.820 ;
        RECT 97.415 329.380 97.795 329.760 ;
        RECT 99.455 329.380 99.835 329.760 ;
        RECT 101.240 329.380 101.620 329.760 ;
        RECT 61.380 329.210 61.760 329.260 ;
        RECT 62.520 329.210 62.900 329.260 ;
        RECT 61.380 328.930 62.900 329.210 ;
        RECT 61.380 328.880 61.760 328.930 ;
        RECT 62.520 328.880 62.900 328.930 ;
        RECT 93.830 329.210 94.210 329.260 ;
        RECT 94.970 329.210 95.350 329.260 ;
        RECT 93.830 328.930 95.350 329.210 ;
        RECT 93.830 328.880 94.210 328.930 ;
        RECT 94.970 328.880 95.350 328.930 ;
        RECT 25.200 327.880 25.580 328.260 ;
        RECT 29.120 327.880 29.500 328.260 ;
        RECT 31.920 327.600 34.160 327.980 ;
        RECT 64.370 327.600 66.610 327.980 ;
        RECT 62.520 327.040 63.040 327.420 ;
        RECT 94.970 327.040 95.490 327.420 ;
        RECT 97.415 326.380 97.795 326.760 ;
        RECT 99.455 326.380 99.835 326.760 ;
        RECT 101.240 326.380 101.620 326.760 ;
        RECT 25.200 324.880 25.580 325.260 ;
        RECT 29.120 324.880 29.500 325.260 ;
        RECT 25.200 321.880 25.580 322.260 ;
        RECT 97.415 320.380 97.795 320.760 ;
        RECT 99.455 320.380 99.835 320.760 ;
        RECT 101.240 320.380 101.620 320.760 ;
        RECT 25.200 318.880 25.580 319.260 ;
        RECT 29.120 318.880 29.500 319.260 ;
        RECT 62.020 318.475 62.900 318.855 ;
        RECT 94.470 318.475 95.350 318.855 ;
        RECT 31.920 317.915 34.160 318.295 ;
        RECT 64.370 317.915 66.610 318.295 ;
        RECT 97.415 317.380 97.795 317.760 ;
        RECT 99.455 317.380 99.835 317.760 ;
        RECT 101.240 317.380 101.620 317.760 ;
        RECT 60.740 316.965 61.120 317.015 ;
        RECT 62.520 316.965 62.900 317.015 ;
        RECT 60.740 316.685 62.900 316.965 ;
        RECT 60.740 316.635 61.120 316.685 ;
        RECT 62.520 316.635 62.900 316.685 ;
        RECT 93.190 316.965 93.570 317.015 ;
        RECT 94.970 316.965 95.350 317.015 ;
        RECT 93.190 316.685 95.350 316.965 ;
        RECT 93.190 316.635 93.570 316.685 ;
        RECT 94.970 316.635 95.350 316.685 ;
        RECT 25.200 315.880 25.580 316.260 ;
        RECT 29.120 315.880 29.500 316.260 ;
        RECT 31.920 316.075 34.160 316.455 ;
        RECT 64.370 316.075 66.610 316.455 ;
        RECT 59.460 315.120 59.840 315.170 ;
        RECT 62.520 315.120 62.900 315.170 ;
        RECT 59.460 314.840 62.900 315.120 ;
        RECT 59.460 314.790 59.840 314.840 ;
        RECT 62.520 314.790 62.900 314.840 ;
        RECT 91.910 315.120 92.290 315.170 ;
        RECT 94.970 315.120 95.350 315.170 ;
        RECT 91.910 314.840 95.350 315.120 ;
        RECT 91.910 314.790 92.290 314.840 ;
        RECT 94.970 314.790 95.350 314.840 ;
        RECT 31.920 314.230 34.160 314.610 ;
        RECT 64.370 314.230 66.610 314.610 ;
        RECT 97.415 314.380 97.795 314.760 ;
        RECT 99.455 314.380 99.835 314.760 ;
        RECT 101.240 314.380 101.620 314.760 ;
        RECT 31.925 313.470 34.165 313.850 ;
        RECT 64.375 313.470 66.615 313.850 ;
        RECT 25.200 312.880 25.580 313.260 ;
        RECT 29.120 312.880 29.500 313.260 ;
        RECT 58.180 312.480 58.560 312.530 ;
        RECT 62.520 312.480 62.900 312.530 ;
        RECT 58.180 312.200 62.900 312.480 ;
        RECT 58.180 312.150 58.560 312.200 ;
        RECT 62.520 312.150 62.900 312.200 ;
        RECT 90.630 312.480 91.010 312.530 ;
        RECT 94.970 312.480 95.350 312.530 ;
        RECT 90.630 312.200 95.350 312.480 ;
        RECT 90.630 312.150 91.010 312.200 ;
        RECT 94.970 312.150 95.350 312.200 ;
        RECT 31.920 311.590 34.160 311.970 ;
        RECT 64.370 311.590 66.610 311.970 ;
        RECT 97.415 311.380 97.795 311.760 ;
        RECT 99.455 311.380 99.835 311.760 ;
        RECT 101.240 311.380 101.620 311.760 ;
        RECT 56.900 310.640 57.280 310.690 ;
        RECT 62.520 310.640 62.900 310.690 ;
        RECT 56.900 310.360 62.900 310.640 ;
        RECT 56.900 310.310 57.280 310.360 ;
        RECT 62.520 310.310 62.900 310.360 ;
        RECT 89.350 310.640 89.730 310.690 ;
        RECT 94.970 310.640 95.350 310.690 ;
        RECT 89.350 310.360 95.350 310.640 ;
        RECT 89.350 310.310 89.730 310.360 ;
        RECT 94.970 310.310 95.350 310.360 ;
        RECT 25.200 309.880 25.580 310.260 ;
        RECT 29.120 309.880 29.500 310.260 ;
        RECT 31.920 309.750 34.160 310.130 ;
        RECT 64.370 309.750 66.610 310.130 ;
        RECT 55.620 308.795 56.000 308.845 ;
        RECT 62.520 308.795 62.900 308.845 ;
        RECT 55.620 308.515 62.900 308.795 ;
        RECT 55.620 308.465 56.000 308.515 ;
        RECT 62.520 308.465 62.900 308.515 ;
        RECT 88.070 308.795 88.450 308.845 ;
        RECT 94.970 308.795 95.350 308.845 ;
        RECT 88.070 308.515 95.350 308.795 ;
        RECT 88.070 308.465 88.450 308.515 ;
        RECT 94.970 308.465 95.350 308.515 ;
        RECT 97.415 308.380 97.795 308.760 ;
        RECT 99.455 308.380 99.835 308.760 ;
        RECT 101.240 308.380 101.620 308.760 ;
        RECT 31.920 307.905 34.160 308.285 ;
        RECT 64.370 307.905 66.610 308.285 ;
        RECT 25.200 306.880 25.580 307.260 ;
        RECT 29.120 306.880 29.500 307.260 ;
        RECT 31.925 307.145 34.165 307.525 ;
        RECT 64.375 307.145 66.615 307.525 ;
        RECT 54.340 306.155 54.720 306.205 ;
        RECT 62.520 306.155 62.900 306.205 ;
        RECT 54.340 305.875 62.900 306.155 ;
        RECT 54.340 305.825 54.720 305.875 ;
        RECT 62.520 305.825 62.900 305.875 ;
        RECT 86.790 306.155 87.170 306.205 ;
        RECT 94.970 306.155 95.350 306.205 ;
        RECT 86.790 305.875 95.350 306.155 ;
        RECT 86.790 305.825 87.170 305.875 ;
        RECT 94.970 305.825 95.350 305.875 ;
        RECT 31.920 305.265 34.160 305.645 ;
        RECT 64.370 305.265 66.610 305.645 ;
        RECT 97.415 305.380 97.795 305.760 ;
        RECT 99.455 305.380 99.835 305.760 ;
        RECT 101.240 305.380 101.620 305.760 ;
        RECT 53.060 304.315 53.440 304.365 ;
        RECT 62.520 304.315 62.900 304.365 ;
        RECT 25.200 303.880 25.580 304.260 ;
        RECT 29.120 303.880 29.500 304.260 ;
        RECT 53.060 304.035 62.900 304.315 ;
        RECT 53.060 303.985 53.440 304.035 ;
        RECT 62.520 303.985 62.900 304.035 ;
        RECT 85.510 304.315 85.890 304.365 ;
        RECT 94.970 304.315 95.350 304.365 ;
        RECT 85.510 304.035 95.350 304.315 ;
        RECT 85.510 303.985 85.890 304.035 ;
        RECT 94.970 303.985 95.350 304.035 ;
        RECT 31.920 303.425 34.160 303.805 ;
        RECT 64.370 303.425 66.610 303.805 ;
        RECT 31.920 302.705 34.160 303.085 ;
        RECT 64.370 302.705 66.610 303.085 ;
        RECT 53.700 302.475 54.080 302.525 ;
        RECT 62.520 302.475 62.900 302.525 ;
        RECT 53.700 302.195 62.900 302.475 ;
        RECT 53.700 302.145 54.080 302.195 ;
        RECT 62.520 302.145 62.900 302.195 ;
        RECT 86.150 302.475 86.530 302.525 ;
        RECT 94.970 302.475 95.350 302.525 ;
        RECT 86.150 302.195 95.350 302.475 ;
        RECT 86.150 302.145 86.530 302.195 ;
        RECT 94.970 302.145 95.350 302.195 ;
        RECT 25.200 300.495 25.580 300.875 ;
        RECT 29.120 300.495 29.500 300.875 ;
        RECT 31.920 300.865 34.160 301.245 ;
        RECT 64.370 300.865 66.610 301.245 ;
        RECT 54.980 300.635 55.360 300.685 ;
        RECT 62.520 300.635 62.900 300.685 ;
        RECT 54.980 300.355 62.900 300.635 ;
        RECT 54.980 300.305 55.360 300.355 ;
        RECT 62.520 300.305 62.900 300.355 ;
        RECT 87.430 300.635 87.810 300.685 ;
        RECT 94.970 300.635 95.350 300.685 ;
        RECT 87.430 300.355 95.350 300.635 ;
        RECT 87.430 300.305 87.810 300.355 ;
        RECT 94.970 300.305 95.350 300.355 ;
        RECT 31.925 298.980 34.165 299.360 ;
        RECT 64.375 298.980 66.615 299.360 ;
        RECT 97.415 298.995 97.795 299.375 ;
        RECT 99.455 298.995 99.835 299.375 ;
        RECT 101.240 298.995 101.620 299.375 ;
        RECT 31.920 298.220 34.160 298.600 ;
        RECT 64.370 298.220 66.610 298.600 ;
        RECT 56.260 297.990 56.640 298.040 ;
        RECT 62.520 297.990 62.900 298.040 ;
        RECT 25.200 297.495 25.580 297.875 ;
        RECT 29.120 297.495 29.500 297.875 ;
        RECT 56.260 297.710 62.900 297.990 ;
        RECT 56.260 297.660 56.640 297.710 ;
        RECT 62.520 297.660 62.900 297.710 ;
        RECT 88.710 297.990 89.090 298.040 ;
        RECT 94.970 297.990 95.350 298.040 ;
        RECT 88.710 297.710 95.350 297.990 ;
        RECT 88.710 297.660 89.090 297.710 ;
        RECT 94.970 297.660 95.350 297.710 ;
        RECT 31.920 296.380 34.160 296.760 ;
        RECT 64.370 296.380 66.610 296.760 ;
        RECT 57.540 296.150 57.920 296.200 ;
        RECT 62.520 296.150 62.900 296.200 ;
        RECT 57.540 295.870 62.900 296.150 ;
        RECT 57.540 295.820 57.920 295.870 ;
        RECT 62.520 295.820 62.900 295.870 ;
        RECT 89.990 296.150 90.370 296.200 ;
        RECT 94.970 296.150 95.350 296.200 ;
        RECT 89.990 295.870 95.350 296.150 ;
        RECT 97.415 295.995 97.795 296.375 ;
        RECT 99.455 295.995 99.835 296.375 ;
        RECT 101.240 295.995 101.620 296.375 ;
        RECT 89.990 295.820 90.370 295.870 ;
        RECT 94.970 295.820 95.350 295.870 ;
        RECT 25.200 294.495 25.580 294.875 ;
        RECT 29.120 294.495 29.500 294.875 ;
        RECT 31.920 294.540 34.160 294.920 ;
        RECT 64.370 294.540 66.610 294.920 ;
        RECT 58.820 294.310 59.200 294.360 ;
        RECT 62.520 294.310 62.900 294.360 ;
        RECT 58.820 294.030 62.900 294.310 ;
        RECT 58.820 293.980 59.200 294.030 ;
        RECT 62.520 293.980 62.900 294.030 ;
        RECT 91.270 294.310 91.650 294.360 ;
        RECT 94.970 294.310 95.350 294.360 ;
        RECT 91.270 294.030 95.350 294.310 ;
        RECT 91.270 293.980 91.650 294.030 ;
        RECT 94.970 293.980 95.350 294.030 ;
        RECT 31.925 292.655 34.165 293.035 ;
        RECT 64.375 292.655 66.615 293.035 ;
        RECT 97.415 292.995 97.795 293.375 ;
        RECT 99.455 292.995 99.835 293.375 ;
        RECT 101.240 292.995 101.620 293.375 ;
        RECT 31.920 291.895 34.160 292.275 ;
        RECT 64.370 291.895 66.610 292.275 ;
        RECT 25.200 291.495 25.580 291.875 ;
        RECT 29.120 291.495 29.500 291.875 ;
        RECT 60.100 291.665 60.480 291.715 ;
        RECT 62.520 291.665 62.900 291.715 ;
        RECT 60.100 291.385 62.900 291.665 ;
        RECT 60.100 291.335 60.480 291.385 ;
        RECT 62.520 291.335 62.900 291.385 ;
        RECT 92.550 291.665 92.930 291.715 ;
        RECT 94.970 291.665 95.350 291.715 ;
        RECT 92.550 291.385 95.350 291.665 ;
        RECT 92.550 291.335 92.930 291.385 ;
        RECT 94.970 291.335 95.350 291.385 ;
        RECT 31.920 290.055 34.160 290.435 ;
        RECT 64.370 290.055 66.610 290.435 ;
        RECT 97.415 289.995 97.795 290.375 ;
        RECT 99.455 289.995 99.835 290.375 ;
        RECT 101.240 289.995 101.620 290.375 ;
        RECT 61.380 289.825 61.760 289.875 ;
        RECT 62.520 289.825 62.900 289.875 ;
        RECT 61.380 289.545 62.900 289.825 ;
        RECT 61.380 289.495 61.760 289.545 ;
        RECT 62.520 289.495 62.900 289.545 ;
        RECT 93.830 289.825 94.210 289.875 ;
        RECT 94.970 289.825 95.350 289.875 ;
        RECT 93.830 289.545 95.350 289.825 ;
        RECT 93.830 289.495 94.210 289.545 ;
        RECT 94.970 289.495 95.350 289.545 ;
        RECT 25.200 288.495 25.580 288.875 ;
        RECT 29.120 288.495 29.500 288.875 ;
        RECT 31.920 288.215 34.160 288.595 ;
        RECT 64.370 288.215 66.610 288.595 ;
        RECT 62.520 287.655 63.040 288.035 ;
        RECT 94.970 287.655 95.490 288.035 ;
        RECT 97.415 286.995 97.795 287.375 ;
        RECT 99.455 286.995 99.835 287.375 ;
        RECT 101.240 286.995 101.620 287.375 ;
        RECT 25.200 285.495 25.580 285.875 ;
        RECT 29.120 285.495 29.500 285.875 ;
        RECT 25.200 282.495 25.580 282.875 ;
        RECT 97.415 280.995 97.795 281.375 ;
        RECT 99.455 280.995 99.835 281.375 ;
        RECT 101.240 280.995 101.620 281.375 ;
        RECT 25.200 279.495 25.580 279.875 ;
        RECT 29.120 279.495 29.500 279.875 ;
        RECT 62.020 279.090 62.900 279.470 ;
        RECT 94.470 279.090 95.350 279.470 ;
        RECT 31.920 278.530 34.160 278.910 ;
        RECT 64.370 278.530 66.610 278.910 ;
        RECT 97.415 277.995 97.795 278.375 ;
        RECT 99.455 277.995 99.835 278.375 ;
        RECT 101.240 277.995 101.620 278.375 ;
        RECT 60.740 277.580 61.120 277.630 ;
        RECT 62.520 277.580 62.900 277.630 ;
        RECT 60.740 277.300 62.900 277.580 ;
        RECT 60.740 277.250 61.120 277.300 ;
        RECT 62.520 277.250 62.900 277.300 ;
        RECT 93.190 277.580 93.570 277.630 ;
        RECT 94.970 277.580 95.350 277.630 ;
        RECT 93.190 277.300 95.350 277.580 ;
        RECT 93.190 277.250 93.570 277.300 ;
        RECT 94.970 277.250 95.350 277.300 ;
        RECT 25.200 276.495 25.580 276.875 ;
        RECT 29.120 276.495 29.500 276.875 ;
        RECT 31.920 276.690 34.160 277.070 ;
        RECT 64.370 276.690 66.610 277.070 ;
        RECT 59.460 275.735 59.840 275.785 ;
        RECT 62.520 275.735 62.900 275.785 ;
        RECT 59.460 275.455 62.900 275.735 ;
        RECT 59.460 275.405 59.840 275.455 ;
        RECT 62.520 275.405 62.900 275.455 ;
        RECT 91.910 275.735 92.290 275.785 ;
        RECT 94.970 275.735 95.350 275.785 ;
        RECT 91.910 275.455 95.350 275.735 ;
        RECT 91.910 275.405 92.290 275.455 ;
        RECT 94.970 275.405 95.350 275.455 ;
        RECT 31.920 274.845 34.160 275.225 ;
        RECT 64.370 274.845 66.610 275.225 ;
        RECT 97.415 274.995 97.795 275.375 ;
        RECT 99.455 274.995 99.835 275.375 ;
        RECT 101.240 274.995 101.620 275.375 ;
        RECT 31.925 274.085 34.165 274.465 ;
        RECT 64.375 274.085 66.615 274.465 ;
        RECT 25.200 273.495 25.580 273.875 ;
        RECT 29.120 273.495 29.500 273.875 ;
        RECT 58.180 273.095 58.560 273.145 ;
        RECT 62.520 273.095 62.900 273.145 ;
        RECT 58.180 272.815 62.900 273.095 ;
        RECT 58.180 272.765 58.560 272.815 ;
        RECT 62.520 272.765 62.900 272.815 ;
        RECT 90.630 273.095 91.010 273.145 ;
        RECT 94.970 273.095 95.350 273.145 ;
        RECT 90.630 272.815 95.350 273.095 ;
        RECT 90.630 272.765 91.010 272.815 ;
        RECT 94.970 272.765 95.350 272.815 ;
        RECT 31.920 272.205 34.160 272.585 ;
        RECT 64.370 272.205 66.610 272.585 ;
        RECT 97.415 271.995 97.795 272.375 ;
        RECT 99.455 271.995 99.835 272.375 ;
        RECT 101.240 271.995 101.620 272.375 ;
        RECT 56.900 271.255 57.280 271.305 ;
        RECT 62.520 271.255 62.900 271.305 ;
        RECT 56.900 270.975 62.900 271.255 ;
        RECT 56.900 270.925 57.280 270.975 ;
        RECT 62.520 270.925 62.900 270.975 ;
        RECT 89.350 271.255 89.730 271.305 ;
        RECT 94.970 271.255 95.350 271.305 ;
        RECT 89.350 270.975 95.350 271.255 ;
        RECT 89.350 270.925 89.730 270.975 ;
        RECT 94.970 270.925 95.350 270.975 ;
        RECT 25.200 270.495 25.580 270.875 ;
        RECT 29.120 270.495 29.500 270.875 ;
        RECT 31.920 270.365 34.160 270.745 ;
        RECT 64.370 270.365 66.610 270.745 ;
        RECT 55.620 269.410 56.000 269.460 ;
        RECT 62.520 269.410 62.900 269.460 ;
        RECT 55.620 269.130 62.900 269.410 ;
        RECT 55.620 269.080 56.000 269.130 ;
        RECT 62.520 269.080 62.900 269.130 ;
        RECT 88.070 269.410 88.450 269.460 ;
        RECT 94.970 269.410 95.350 269.460 ;
        RECT 88.070 269.130 95.350 269.410 ;
        RECT 88.070 269.080 88.450 269.130 ;
        RECT 94.970 269.080 95.350 269.130 ;
        RECT 97.415 268.995 97.795 269.375 ;
        RECT 99.455 268.995 99.835 269.375 ;
        RECT 101.240 268.995 101.620 269.375 ;
        RECT 31.920 268.520 34.160 268.900 ;
        RECT 64.370 268.520 66.610 268.900 ;
        RECT 25.200 267.495 25.580 267.875 ;
        RECT 29.120 267.495 29.500 267.875 ;
        RECT 31.925 267.760 34.165 268.140 ;
        RECT 64.375 267.760 66.615 268.140 ;
        RECT 54.340 266.770 54.720 266.820 ;
        RECT 62.520 266.770 62.900 266.820 ;
        RECT 54.340 266.490 62.900 266.770 ;
        RECT 54.340 266.440 54.720 266.490 ;
        RECT 62.520 266.440 62.900 266.490 ;
        RECT 86.790 266.770 87.170 266.820 ;
        RECT 94.970 266.770 95.350 266.820 ;
        RECT 86.790 266.490 95.350 266.770 ;
        RECT 86.790 266.440 87.170 266.490 ;
        RECT 94.970 266.440 95.350 266.490 ;
        RECT 31.920 265.880 34.160 266.260 ;
        RECT 64.370 265.880 66.610 266.260 ;
        RECT 97.415 265.995 97.795 266.375 ;
        RECT 99.455 265.995 99.835 266.375 ;
        RECT 101.240 265.995 101.620 266.375 ;
        RECT 53.060 264.930 53.440 264.980 ;
        RECT 62.520 264.930 62.900 264.980 ;
        RECT 25.200 264.495 25.580 264.875 ;
        RECT 29.120 264.495 29.500 264.875 ;
        RECT 53.060 264.650 62.900 264.930 ;
        RECT 53.060 264.600 53.440 264.650 ;
        RECT 62.520 264.600 62.900 264.650 ;
        RECT 85.510 264.930 85.890 264.980 ;
        RECT 94.970 264.930 95.350 264.980 ;
        RECT 85.510 264.650 95.350 264.930 ;
        RECT 85.510 264.600 85.890 264.650 ;
        RECT 94.970 264.600 95.350 264.650 ;
        RECT 31.920 264.040 34.160 264.420 ;
        RECT 64.370 264.040 66.610 264.420 ;
        RECT 31.920 263.320 34.160 263.700 ;
        RECT 64.370 263.320 66.610 263.700 ;
        RECT 53.700 263.090 54.080 263.140 ;
        RECT 62.520 263.090 62.900 263.140 ;
        RECT 53.700 262.810 62.900 263.090 ;
        RECT 53.700 262.760 54.080 262.810 ;
        RECT 62.520 262.760 62.900 262.810 ;
        RECT 86.150 263.090 86.530 263.140 ;
        RECT 94.970 263.090 95.350 263.140 ;
        RECT 86.150 262.810 95.350 263.090 ;
        RECT 86.150 262.760 86.530 262.810 ;
        RECT 94.970 262.760 95.350 262.810 ;
        RECT 25.200 261.110 25.580 261.490 ;
        RECT 29.120 261.110 29.500 261.490 ;
        RECT 31.920 261.480 34.160 261.860 ;
        RECT 64.370 261.480 66.610 261.860 ;
        RECT 54.980 261.250 55.360 261.300 ;
        RECT 62.520 261.250 62.900 261.300 ;
        RECT 54.980 260.970 62.900 261.250 ;
        RECT 54.980 260.920 55.360 260.970 ;
        RECT 62.520 260.920 62.900 260.970 ;
        RECT 87.430 261.250 87.810 261.300 ;
        RECT 94.970 261.250 95.350 261.300 ;
        RECT 87.430 260.970 95.350 261.250 ;
        RECT 87.430 260.920 87.810 260.970 ;
        RECT 94.970 260.920 95.350 260.970 ;
        RECT 31.925 259.595 34.165 259.975 ;
        RECT 64.375 259.595 66.615 259.975 ;
        RECT 97.415 259.610 97.795 259.990 ;
        RECT 99.455 259.610 99.835 259.990 ;
        RECT 101.240 259.610 101.620 259.990 ;
        RECT 31.920 258.835 34.160 259.215 ;
        RECT 64.370 258.835 66.610 259.215 ;
        RECT 56.260 258.605 56.640 258.655 ;
        RECT 62.520 258.605 62.900 258.655 ;
        RECT 25.200 258.110 25.580 258.490 ;
        RECT 29.120 258.110 29.500 258.490 ;
        RECT 56.260 258.325 62.900 258.605 ;
        RECT 56.260 258.275 56.640 258.325 ;
        RECT 62.520 258.275 62.900 258.325 ;
        RECT 88.710 258.605 89.090 258.655 ;
        RECT 94.970 258.605 95.350 258.655 ;
        RECT 88.710 258.325 95.350 258.605 ;
        RECT 88.710 258.275 89.090 258.325 ;
        RECT 94.970 258.275 95.350 258.325 ;
        RECT 31.920 256.995 34.160 257.375 ;
        RECT 64.370 256.995 66.610 257.375 ;
        RECT 57.540 256.765 57.920 256.815 ;
        RECT 62.520 256.765 62.900 256.815 ;
        RECT 57.540 256.485 62.900 256.765 ;
        RECT 57.540 256.435 57.920 256.485 ;
        RECT 62.520 256.435 62.900 256.485 ;
        RECT 89.990 256.765 90.370 256.815 ;
        RECT 94.970 256.765 95.350 256.815 ;
        RECT 89.990 256.485 95.350 256.765 ;
        RECT 97.415 256.610 97.795 256.990 ;
        RECT 99.455 256.610 99.835 256.990 ;
        RECT 101.240 256.610 101.620 256.990 ;
        RECT 89.990 256.435 90.370 256.485 ;
        RECT 94.970 256.435 95.350 256.485 ;
        RECT 25.200 255.110 25.580 255.490 ;
        RECT 29.120 255.110 29.500 255.490 ;
        RECT 31.920 255.155 34.160 255.535 ;
        RECT 64.370 255.155 66.610 255.535 ;
        RECT 58.820 254.925 59.200 254.975 ;
        RECT 62.520 254.925 62.900 254.975 ;
        RECT 58.820 254.645 62.900 254.925 ;
        RECT 58.820 254.595 59.200 254.645 ;
        RECT 62.520 254.595 62.900 254.645 ;
        RECT 91.270 254.925 91.650 254.975 ;
        RECT 94.970 254.925 95.350 254.975 ;
        RECT 91.270 254.645 95.350 254.925 ;
        RECT 91.270 254.595 91.650 254.645 ;
        RECT 94.970 254.595 95.350 254.645 ;
        RECT 31.925 253.270 34.165 253.650 ;
        RECT 64.375 253.270 66.615 253.650 ;
        RECT 97.415 253.610 97.795 253.990 ;
        RECT 99.455 253.610 99.835 253.990 ;
        RECT 101.240 253.610 101.620 253.990 ;
        RECT 31.920 252.510 34.160 252.890 ;
        RECT 64.370 252.510 66.610 252.890 ;
        RECT 25.200 252.110 25.580 252.490 ;
        RECT 29.120 252.110 29.500 252.490 ;
        RECT 60.100 252.280 60.480 252.330 ;
        RECT 62.520 252.280 62.900 252.330 ;
        RECT 60.100 252.000 62.900 252.280 ;
        RECT 60.100 251.950 60.480 252.000 ;
        RECT 62.520 251.950 62.900 252.000 ;
        RECT 92.550 252.280 92.930 252.330 ;
        RECT 94.970 252.280 95.350 252.330 ;
        RECT 92.550 252.000 95.350 252.280 ;
        RECT 92.550 251.950 92.930 252.000 ;
        RECT 94.970 251.950 95.350 252.000 ;
        RECT 31.920 250.670 34.160 251.050 ;
        RECT 64.370 250.670 66.610 251.050 ;
        RECT 97.415 250.610 97.795 250.990 ;
        RECT 99.455 250.610 99.835 250.990 ;
        RECT 101.240 250.610 101.620 250.990 ;
        RECT 61.380 250.440 61.760 250.490 ;
        RECT 62.520 250.440 62.900 250.490 ;
        RECT 61.380 250.160 62.900 250.440 ;
        RECT 61.380 250.110 61.760 250.160 ;
        RECT 62.520 250.110 62.900 250.160 ;
        RECT 93.830 250.440 94.210 250.490 ;
        RECT 94.970 250.440 95.350 250.490 ;
        RECT 93.830 250.160 95.350 250.440 ;
        RECT 93.830 250.110 94.210 250.160 ;
        RECT 94.970 250.110 95.350 250.160 ;
        RECT 25.200 249.110 25.580 249.490 ;
        RECT 29.120 249.110 29.500 249.490 ;
        RECT 31.920 248.830 34.160 249.210 ;
        RECT 64.370 248.830 66.610 249.210 ;
        RECT 62.520 248.270 63.040 248.650 ;
        RECT 94.970 248.270 95.490 248.650 ;
        RECT 97.415 247.610 97.795 247.990 ;
        RECT 99.455 247.610 99.835 247.990 ;
        RECT 101.240 247.610 101.620 247.990 ;
        RECT 25.200 246.110 25.580 246.490 ;
        RECT 29.120 246.110 29.500 246.490 ;
        RECT 25.200 243.110 25.580 243.490 ;
        RECT 97.415 241.610 97.795 241.990 ;
        RECT 99.455 241.610 99.835 241.990 ;
        RECT 101.240 241.610 101.620 241.990 ;
        RECT 25.200 240.110 25.580 240.490 ;
        RECT 29.120 240.110 29.500 240.490 ;
        RECT 62.020 239.705 62.900 240.085 ;
        RECT 94.470 239.705 95.350 240.085 ;
        RECT 31.920 239.145 34.160 239.525 ;
        RECT 64.370 239.145 66.610 239.525 ;
        RECT 97.415 238.610 97.795 238.990 ;
        RECT 99.455 238.610 99.835 238.990 ;
        RECT 101.240 238.610 101.620 238.990 ;
        RECT 60.740 238.195 61.120 238.245 ;
        RECT 62.520 238.195 62.900 238.245 ;
        RECT 60.740 237.915 62.900 238.195 ;
        RECT 60.740 237.865 61.120 237.915 ;
        RECT 62.520 237.865 62.900 237.915 ;
        RECT 93.190 238.195 93.570 238.245 ;
        RECT 94.970 238.195 95.350 238.245 ;
        RECT 93.190 237.915 95.350 238.195 ;
        RECT 93.190 237.865 93.570 237.915 ;
        RECT 94.970 237.865 95.350 237.915 ;
        RECT 25.200 237.110 25.580 237.490 ;
        RECT 29.120 237.110 29.500 237.490 ;
        RECT 31.920 237.305 34.160 237.685 ;
        RECT 64.370 237.305 66.610 237.685 ;
        RECT 59.460 236.350 59.840 236.400 ;
        RECT 62.520 236.350 62.900 236.400 ;
        RECT 59.460 236.070 62.900 236.350 ;
        RECT 59.460 236.020 59.840 236.070 ;
        RECT 62.520 236.020 62.900 236.070 ;
        RECT 91.910 236.350 92.290 236.400 ;
        RECT 94.970 236.350 95.350 236.400 ;
        RECT 91.910 236.070 95.350 236.350 ;
        RECT 91.910 236.020 92.290 236.070 ;
        RECT 94.970 236.020 95.350 236.070 ;
        RECT 31.920 235.460 34.160 235.840 ;
        RECT 64.370 235.460 66.610 235.840 ;
        RECT 97.415 235.610 97.795 235.990 ;
        RECT 99.455 235.610 99.835 235.990 ;
        RECT 101.240 235.610 101.620 235.990 ;
        RECT 31.925 234.700 34.165 235.080 ;
        RECT 64.375 234.700 66.615 235.080 ;
        RECT 25.200 234.110 25.580 234.490 ;
        RECT 29.120 234.110 29.500 234.490 ;
        RECT 58.180 233.710 58.560 233.760 ;
        RECT 62.520 233.710 62.900 233.760 ;
        RECT 58.180 233.430 62.900 233.710 ;
        RECT 58.180 233.380 58.560 233.430 ;
        RECT 62.520 233.380 62.900 233.430 ;
        RECT 90.630 233.710 91.010 233.760 ;
        RECT 94.970 233.710 95.350 233.760 ;
        RECT 90.630 233.430 95.350 233.710 ;
        RECT 90.630 233.380 91.010 233.430 ;
        RECT 94.970 233.380 95.350 233.430 ;
        RECT 31.920 232.820 34.160 233.200 ;
        RECT 64.370 232.820 66.610 233.200 ;
        RECT 97.415 232.610 97.795 232.990 ;
        RECT 99.455 232.610 99.835 232.990 ;
        RECT 101.240 232.610 101.620 232.990 ;
        RECT 56.900 231.870 57.280 231.920 ;
        RECT 62.520 231.870 62.900 231.920 ;
        RECT 56.900 231.590 62.900 231.870 ;
        RECT 56.900 231.540 57.280 231.590 ;
        RECT 62.520 231.540 62.900 231.590 ;
        RECT 89.350 231.870 89.730 231.920 ;
        RECT 94.970 231.870 95.350 231.920 ;
        RECT 89.350 231.590 95.350 231.870 ;
        RECT 89.350 231.540 89.730 231.590 ;
        RECT 94.970 231.540 95.350 231.590 ;
        RECT 25.200 231.110 25.580 231.490 ;
        RECT 29.120 231.110 29.500 231.490 ;
        RECT 31.920 230.980 34.160 231.360 ;
        RECT 64.370 230.980 66.610 231.360 ;
        RECT 55.620 230.025 56.000 230.075 ;
        RECT 62.520 230.025 62.900 230.075 ;
        RECT 55.620 229.745 62.900 230.025 ;
        RECT 55.620 229.695 56.000 229.745 ;
        RECT 62.520 229.695 62.900 229.745 ;
        RECT 88.070 230.025 88.450 230.075 ;
        RECT 94.970 230.025 95.350 230.075 ;
        RECT 88.070 229.745 95.350 230.025 ;
        RECT 88.070 229.695 88.450 229.745 ;
        RECT 94.970 229.695 95.350 229.745 ;
        RECT 97.415 229.610 97.795 229.990 ;
        RECT 99.455 229.610 99.835 229.990 ;
        RECT 101.240 229.610 101.620 229.990 ;
        RECT 31.920 229.135 34.160 229.515 ;
        RECT 64.370 229.135 66.610 229.515 ;
        RECT 25.200 228.110 25.580 228.490 ;
        RECT 29.120 228.110 29.500 228.490 ;
        RECT 31.925 228.375 34.165 228.755 ;
        RECT 64.375 228.375 66.615 228.755 ;
        RECT 54.340 227.385 54.720 227.435 ;
        RECT 62.520 227.385 62.900 227.435 ;
        RECT 54.340 227.105 62.900 227.385 ;
        RECT 54.340 227.055 54.720 227.105 ;
        RECT 62.520 227.055 62.900 227.105 ;
        RECT 86.790 227.385 87.170 227.435 ;
        RECT 94.970 227.385 95.350 227.435 ;
        RECT 86.790 227.105 95.350 227.385 ;
        RECT 86.790 227.055 87.170 227.105 ;
        RECT 94.970 227.055 95.350 227.105 ;
        RECT 31.920 226.495 34.160 226.875 ;
        RECT 64.370 226.495 66.610 226.875 ;
        RECT 97.415 226.610 97.795 226.990 ;
        RECT 99.455 226.610 99.835 226.990 ;
        RECT 101.240 226.610 101.620 226.990 ;
        RECT 53.060 225.545 53.440 225.595 ;
        RECT 62.520 225.545 62.900 225.595 ;
        RECT 25.200 225.110 25.580 225.490 ;
        RECT 29.120 225.110 29.500 225.490 ;
        RECT 53.060 225.265 62.900 225.545 ;
        RECT 53.060 225.215 53.440 225.265 ;
        RECT 62.520 225.215 62.900 225.265 ;
        RECT 85.510 225.545 85.890 225.595 ;
        RECT 94.970 225.545 95.350 225.595 ;
        RECT 85.510 225.265 95.350 225.545 ;
        RECT 85.510 225.215 85.890 225.265 ;
        RECT 94.970 225.215 95.350 225.265 ;
        RECT 31.920 224.655 34.160 225.035 ;
        RECT 64.370 224.655 66.610 225.035 ;
        RECT 31.920 223.935 34.160 224.315 ;
        RECT 64.370 223.935 66.610 224.315 ;
        RECT 53.700 223.705 54.080 223.755 ;
        RECT 62.520 223.705 62.900 223.755 ;
        RECT 53.700 223.425 62.900 223.705 ;
        RECT 53.700 223.375 54.080 223.425 ;
        RECT 62.520 223.375 62.900 223.425 ;
        RECT 86.150 223.705 86.530 223.755 ;
        RECT 94.970 223.705 95.350 223.755 ;
        RECT 86.150 223.425 95.350 223.705 ;
        RECT 86.150 223.375 86.530 223.425 ;
        RECT 94.970 223.375 95.350 223.425 ;
        RECT 25.200 221.725 25.580 222.105 ;
        RECT 29.120 221.725 29.500 222.105 ;
        RECT 31.920 222.095 34.160 222.475 ;
        RECT 64.370 222.095 66.610 222.475 ;
        RECT 54.980 221.865 55.360 221.915 ;
        RECT 62.520 221.865 62.900 221.915 ;
        RECT 54.980 221.585 62.900 221.865 ;
        RECT 54.980 221.535 55.360 221.585 ;
        RECT 62.520 221.535 62.900 221.585 ;
        RECT 87.430 221.865 87.810 221.915 ;
        RECT 94.970 221.865 95.350 221.915 ;
        RECT 87.430 221.585 95.350 221.865 ;
        RECT 87.430 221.535 87.810 221.585 ;
        RECT 94.970 221.535 95.350 221.585 ;
        RECT 31.925 220.210 34.165 220.590 ;
        RECT 64.375 220.210 66.615 220.590 ;
        RECT 97.415 220.225 97.795 220.605 ;
        RECT 99.455 220.225 99.835 220.605 ;
        RECT 101.240 220.225 101.620 220.605 ;
        RECT 31.920 219.450 34.160 219.830 ;
        RECT 64.370 219.450 66.610 219.830 ;
        RECT 56.260 219.220 56.640 219.270 ;
        RECT 62.520 219.220 62.900 219.270 ;
        RECT 25.200 218.725 25.580 219.105 ;
        RECT 29.120 218.725 29.500 219.105 ;
        RECT 56.260 218.940 62.900 219.220 ;
        RECT 56.260 218.890 56.640 218.940 ;
        RECT 62.520 218.890 62.900 218.940 ;
        RECT 88.710 219.220 89.090 219.270 ;
        RECT 94.970 219.220 95.350 219.270 ;
        RECT 88.710 218.940 95.350 219.220 ;
        RECT 88.710 218.890 89.090 218.940 ;
        RECT 94.970 218.890 95.350 218.940 ;
        RECT 31.920 217.610 34.160 217.990 ;
        RECT 64.370 217.610 66.610 217.990 ;
        RECT 57.540 217.380 57.920 217.430 ;
        RECT 62.520 217.380 62.900 217.430 ;
        RECT 57.540 217.100 62.900 217.380 ;
        RECT 57.540 217.050 57.920 217.100 ;
        RECT 62.520 217.050 62.900 217.100 ;
        RECT 89.990 217.380 90.370 217.430 ;
        RECT 94.970 217.380 95.350 217.430 ;
        RECT 89.990 217.100 95.350 217.380 ;
        RECT 97.415 217.225 97.795 217.605 ;
        RECT 99.455 217.225 99.835 217.605 ;
        RECT 101.240 217.225 101.620 217.605 ;
        RECT 89.990 217.050 90.370 217.100 ;
        RECT 94.970 217.050 95.350 217.100 ;
        RECT 25.200 215.725 25.580 216.105 ;
        RECT 29.120 215.725 29.500 216.105 ;
        RECT 31.920 215.770 34.160 216.150 ;
        RECT 64.370 215.770 66.610 216.150 ;
        RECT 58.820 215.540 59.200 215.590 ;
        RECT 62.520 215.540 62.900 215.590 ;
        RECT 58.820 215.260 62.900 215.540 ;
        RECT 58.820 215.210 59.200 215.260 ;
        RECT 62.520 215.210 62.900 215.260 ;
        RECT 91.270 215.540 91.650 215.590 ;
        RECT 94.970 215.540 95.350 215.590 ;
        RECT 91.270 215.260 95.350 215.540 ;
        RECT 91.270 215.210 91.650 215.260 ;
        RECT 94.970 215.210 95.350 215.260 ;
        RECT 31.925 213.885 34.165 214.265 ;
        RECT 64.375 213.885 66.615 214.265 ;
        RECT 97.415 214.225 97.795 214.605 ;
        RECT 99.455 214.225 99.835 214.605 ;
        RECT 101.240 214.225 101.620 214.605 ;
        RECT 31.920 213.125 34.160 213.505 ;
        RECT 64.370 213.125 66.610 213.505 ;
        RECT 25.200 212.725 25.580 213.105 ;
        RECT 29.120 212.725 29.500 213.105 ;
        RECT 60.100 212.895 60.480 212.945 ;
        RECT 62.520 212.895 62.900 212.945 ;
        RECT 60.100 212.615 62.900 212.895 ;
        RECT 60.100 212.565 60.480 212.615 ;
        RECT 62.520 212.565 62.900 212.615 ;
        RECT 92.550 212.895 92.930 212.945 ;
        RECT 94.970 212.895 95.350 212.945 ;
        RECT 92.550 212.615 95.350 212.895 ;
        RECT 92.550 212.565 92.930 212.615 ;
        RECT 94.970 212.565 95.350 212.615 ;
        RECT 31.920 211.285 34.160 211.665 ;
        RECT 64.370 211.285 66.610 211.665 ;
        RECT 97.415 211.225 97.795 211.605 ;
        RECT 99.455 211.225 99.835 211.605 ;
        RECT 101.240 211.225 101.620 211.605 ;
        RECT 61.380 211.055 61.760 211.105 ;
        RECT 62.520 211.055 62.900 211.105 ;
        RECT 61.380 210.775 62.900 211.055 ;
        RECT 61.380 210.725 61.760 210.775 ;
        RECT 62.520 210.725 62.900 210.775 ;
        RECT 93.830 211.055 94.210 211.105 ;
        RECT 94.970 211.055 95.350 211.105 ;
        RECT 93.830 210.775 95.350 211.055 ;
        RECT 93.830 210.725 94.210 210.775 ;
        RECT 94.970 210.725 95.350 210.775 ;
        RECT 25.200 209.725 25.580 210.105 ;
        RECT 29.120 209.725 29.500 210.105 ;
        RECT 31.920 209.445 34.160 209.825 ;
        RECT 64.370 209.445 66.610 209.825 ;
        RECT 62.520 208.885 63.040 209.265 ;
        RECT 94.970 208.885 95.490 209.265 ;
        RECT 97.415 208.225 97.795 208.605 ;
        RECT 99.455 208.225 99.835 208.605 ;
        RECT 101.240 208.225 101.620 208.605 ;
        RECT 25.200 206.725 25.580 207.105 ;
        RECT 29.120 206.725 29.500 207.105 ;
        RECT 25.200 203.725 25.580 204.105 ;
        RECT 97.415 202.225 97.795 202.605 ;
        RECT 99.455 202.225 99.835 202.605 ;
        RECT 101.240 202.225 101.620 202.605 ;
        RECT 25.200 200.725 25.580 201.105 ;
        RECT 29.120 200.725 29.500 201.105 ;
        RECT 62.020 200.320 62.900 200.700 ;
        RECT 94.470 200.320 95.350 200.700 ;
        RECT 31.920 199.760 34.160 200.140 ;
        RECT 64.370 199.760 66.610 200.140 ;
        RECT 97.415 199.225 97.795 199.605 ;
        RECT 99.455 199.225 99.835 199.605 ;
        RECT 101.240 199.225 101.620 199.605 ;
        RECT 60.740 198.810 61.120 198.860 ;
        RECT 62.520 198.810 62.900 198.860 ;
        RECT 60.740 198.530 62.900 198.810 ;
        RECT 60.740 198.480 61.120 198.530 ;
        RECT 62.520 198.480 62.900 198.530 ;
        RECT 93.190 198.810 93.570 198.860 ;
        RECT 94.970 198.810 95.350 198.860 ;
        RECT 93.190 198.530 95.350 198.810 ;
        RECT 93.190 198.480 93.570 198.530 ;
        RECT 94.970 198.480 95.350 198.530 ;
        RECT 25.200 197.725 25.580 198.105 ;
        RECT 29.120 197.725 29.500 198.105 ;
        RECT 31.920 197.920 34.160 198.300 ;
        RECT 64.370 197.920 66.610 198.300 ;
        RECT 59.460 196.965 59.840 197.015 ;
        RECT 62.520 196.965 62.900 197.015 ;
        RECT 59.460 196.685 62.900 196.965 ;
        RECT 59.460 196.635 59.840 196.685 ;
        RECT 62.520 196.635 62.900 196.685 ;
        RECT 91.910 196.965 92.290 197.015 ;
        RECT 94.970 196.965 95.350 197.015 ;
        RECT 91.910 196.685 95.350 196.965 ;
        RECT 91.910 196.635 92.290 196.685 ;
        RECT 94.970 196.635 95.350 196.685 ;
        RECT 31.920 196.075 34.160 196.455 ;
        RECT 64.370 196.075 66.610 196.455 ;
        RECT 97.415 196.225 97.795 196.605 ;
        RECT 99.455 196.225 99.835 196.605 ;
        RECT 101.240 196.225 101.620 196.605 ;
        RECT 31.925 195.315 34.165 195.695 ;
        RECT 64.375 195.315 66.615 195.695 ;
        RECT 25.200 194.725 25.580 195.105 ;
        RECT 29.120 194.725 29.500 195.105 ;
        RECT 58.180 194.325 58.560 194.375 ;
        RECT 62.520 194.325 62.900 194.375 ;
        RECT 58.180 194.045 62.900 194.325 ;
        RECT 58.180 193.995 58.560 194.045 ;
        RECT 62.520 193.995 62.900 194.045 ;
        RECT 90.630 194.325 91.010 194.375 ;
        RECT 94.970 194.325 95.350 194.375 ;
        RECT 90.630 194.045 95.350 194.325 ;
        RECT 90.630 193.995 91.010 194.045 ;
        RECT 94.970 193.995 95.350 194.045 ;
        RECT 31.920 193.435 34.160 193.815 ;
        RECT 64.370 193.435 66.610 193.815 ;
        RECT 97.415 193.225 97.795 193.605 ;
        RECT 99.455 193.225 99.835 193.605 ;
        RECT 101.240 193.225 101.620 193.605 ;
        RECT 56.900 192.485 57.280 192.535 ;
        RECT 62.520 192.485 62.900 192.535 ;
        RECT 56.900 192.205 62.900 192.485 ;
        RECT 56.900 192.155 57.280 192.205 ;
        RECT 62.520 192.155 62.900 192.205 ;
        RECT 89.350 192.485 89.730 192.535 ;
        RECT 94.970 192.485 95.350 192.535 ;
        RECT 89.350 192.205 95.350 192.485 ;
        RECT 89.350 192.155 89.730 192.205 ;
        RECT 94.970 192.155 95.350 192.205 ;
        RECT 25.200 191.725 25.580 192.105 ;
        RECT 29.120 191.725 29.500 192.105 ;
        RECT 31.920 191.595 34.160 191.975 ;
        RECT 64.370 191.595 66.610 191.975 ;
        RECT 55.620 190.640 56.000 190.690 ;
        RECT 62.520 190.640 62.900 190.690 ;
        RECT 55.620 190.360 62.900 190.640 ;
        RECT 55.620 190.310 56.000 190.360 ;
        RECT 62.520 190.310 62.900 190.360 ;
        RECT 88.070 190.640 88.450 190.690 ;
        RECT 94.970 190.640 95.350 190.690 ;
        RECT 88.070 190.360 95.350 190.640 ;
        RECT 88.070 190.310 88.450 190.360 ;
        RECT 94.970 190.310 95.350 190.360 ;
        RECT 97.415 190.225 97.795 190.605 ;
        RECT 99.455 190.225 99.835 190.605 ;
        RECT 101.240 190.225 101.620 190.605 ;
        RECT 31.920 189.750 34.160 190.130 ;
        RECT 64.370 189.750 66.610 190.130 ;
        RECT 25.200 188.725 25.580 189.105 ;
        RECT 29.120 188.725 29.500 189.105 ;
        RECT 31.925 188.990 34.165 189.370 ;
        RECT 64.375 188.990 66.615 189.370 ;
        RECT 54.340 188.000 54.720 188.050 ;
        RECT 62.520 188.000 62.900 188.050 ;
        RECT 54.340 187.720 62.900 188.000 ;
        RECT 54.340 187.670 54.720 187.720 ;
        RECT 62.520 187.670 62.900 187.720 ;
        RECT 86.790 188.000 87.170 188.050 ;
        RECT 94.970 188.000 95.350 188.050 ;
        RECT 86.790 187.720 95.350 188.000 ;
        RECT 86.790 187.670 87.170 187.720 ;
        RECT 94.970 187.670 95.350 187.720 ;
        RECT 31.920 187.110 34.160 187.490 ;
        RECT 64.370 187.110 66.610 187.490 ;
        RECT 97.415 187.225 97.795 187.605 ;
        RECT 99.455 187.225 99.835 187.605 ;
        RECT 101.240 187.225 101.620 187.605 ;
        RECT 53.060 186.160 53.440 186.210 ;
        RECT 62.520 186.160 62.900 186.210 ;
        RECT 25.200 185.725 25.580 186.105 ;
        RECT 29.120 185.725 29.500 186.105 ;
        RECT 53.060 185.880 62.900 186.160 ;
        RECT 53.060 185.830 53.440 185.880 ;
        RECT 62.520 185.830 62.900 185.880 ;
        RECT 85.510 186.160 85.890 186.210 ;
        RECT 94.970 186.160 95.350 186.210 ;
        RECT 85.510 185.880 95.350 186.160 ;
        RECT 85.510 185.830 85.890 185.880 ;
        RECT 94.970 185.830 95.350 185.880 ;
        RECT 31.920 185.270 34.160 185.650 ;
        RECT 64.370 185.270 66.610 185.650 ;
        RECT 31.920 184.550 34.160 184.930 ;
        RECT 64.370 184.550 66.610 184.930 ;
        RECT 53.700 184.320 54.080 184.370 ;
        RECT 62.520 184.320 62.900 184.370 ;
        RECT 53.700 184.040 62.900 184.320 ;
        RECT 53.700 183.990 54.080 184.040 ;
        RECT 62.520 183.990 62.900 184.040 ;
        RECT 86.150 184.320 86.530 184.370 ;
        RECT 94.970 184.320 95.350 184.370 ;
        RECT 86.150 184.040 95.350 184.320 ;
        RECT 86.150 183.990 86.530 184.040 ;
        RECT 94.970 183.990 95.350 184.040 ;
        RECT 25.200 182.340 25.580 182.720 ;
        RECT 29.120 182.340 29.500 182.720 ;
        RECT 31.920 182.710 34.160 183.090 ;
        RECT 64.370 182.710 66.610 183.090 ;
        RECT 54.980 182.480 55.360 182.530 ;
        RECT 62.520 182.480 62.900 182.530 ;
        RECT 54.980 182.200 62.900 182.480 ;
        RECT 54.980 182.150 55.360 182.200 ;
        RECT 62.520 182.150 62.900 182.200 ;
        RECT 87.430 182.480 87.810 182.530 ;
        RECT 94.970 182.480 95.350 182.530 ;
        RECT 87.430 182.200 95.350 182.480 ;
        RECT 87.430 182.150 87.810 182.200 ;
        RECT 94.970 182.150 95.350 182.200 ;
        RECT 31.925 180.825 34.165 181.205 ;
        RECT 64.375 180.825 66.615 181.205 ;
        RECT 97.415 180.840 97.795 181.220 ;
        RECT 99.455 180.840 99.835 181.220 ;
        RECT 101.240 180.840 101.620 181.220 ;
        RECT 31.920 180.065 34.160 180.445 ;
        RECT 64.370 180.065 66.610 180.445 ;
        RECT 56.260 179.835 56.640 179.885 ;
        RECT 62.520 179.835 62.900 179.885 ;
        RECT 25.200 179.340 25.580 179.720 ;
        RECT 29.120 179.340 29.500 179.720 ;
        RECT 56.260 179.555 62.900 179.835 ;
        RECT 56.260 179.505 56.640 179.555 ;
        RECT 62.520 179.505 62.900 179.555 ;
        RECT 88.710 179.835 89.090 179.885 ;
        RECT 94.970 179.835 95.350 179.885 ;
        RECT 88.710 179.555 95.350 179.835 ;
        RECT 88.710 179.505 89.090 179.555 ;
        RECT 94.970 179.505 95.350 179.555 ;
        RECT 31.920 178.225 34.160 178.605 ;
        RECT 64.370 178.225 66.610 178.605 ;
        RECT 57.540 177.995 57.920 178.045 ;
        RECT 62.520 177.995 62.900 178.045 ;
        RECT 57.540 177.715 62.900 177.995 ;
        RECT 57.540 177.665 57.920 177.715 ;
        RECT 62.520 177.665 62.900 177.715 ;
        RECT 89.990 177.995 90.370 178.045 ;
        RECT 94.970 177.995 95.350 178.045 ;
        RECT 89.990 177.715 95.350 177.995 ;
        RECT 97.415 177.840 97.795 178.220 ;
        RECT 99.455 177.840 99.835 178.220 ;
        RECT 101.240 177.840 101.620 178.220 ;
        RECT 89.990 177.665 90.370 177.715 ;
        RECT 94.970 177.665 95.350 177.715 ;
        RECT 25.200 176.340 25.580 176.720 ;
        RECT 29.120 176.340 29.500 176.720 ;
        RECT 31.920 176.385 34.160 176.765 ;
        RECT 64.370 176.385 66.610 176.765 ;
        RECT 58.820 176.155 59.200 176.205 ;
        RECT 62.520 176.155 62.900 176.205 ;
        RECT 58.820 175.875 62.900 176.155 ;
        RECT 58.820 175.825 59.200 175.875 ;
        RECT 62.520 175.825 62.900 175.875 ;
        RECT 91.270 176.155 91.650 176.205 ;
        RECT 94.970 176.155 95.350 176.205 ;
        RECT 91.270 175.875 95.350 176.155 ;
        RECT 91.270 175.825 91.650 175.875 ;
        RECT 94.970 175.825 95.350 175.875 ;
        RECT 31.925 174.500 34.165 174.880 ;
        RECT 64.375 174.500 66.615 174.880 ;
        RECT 97.415 174.840 97.795 175.220 ;
        RECT 99.455 174.840 99.835 175.220 ;
        RECT 101.240 174.840 101.620 175.220 ;
        RECT 31.920 173.740 34.160 174.120 ;
        RECT 64.370 173.740 66.610 174.120 ;
        RECT 25.200 173.340 25.580 173.720 ;
        RECT 29.120 173.340 29.500 173.720 ;
        RECT 60.100 173.510 60.480 173.560 ;
        RECT 62.520 173.510 62.900 173.560 ;
        RECT 60.100 173.230 62.900 173.510 ;
        RECT 60.100 173.180 60.480 173.230 ;
        RECT 62.520 173.180 62.900 173.230 ;
        RECT 92.550 173.510 92.930 173.560 ;
        RECT 94.970 173.510 95.350 173.560 ;
        RECT 92.550 173.230 95.350 173.510 ;
        RECT 92.550 173.180 92.930 173.230 ;
        RECT 94.970 173.180 95.350 173.230 ;
        RECT 31.920 171.900 34.160 172.280 ;
        RECT 64.370 171.900 66.610 172.280 ;
        RECT 97.415 171.840 97.795 172.220 ;
        RECT 99.455 171.840 99.835 172.220 ;
        RECT 101.240 171.840 101.620 172.220 ;
        RECT 61.380 171.670 61.760 171.720 ;
        RECT 62.520 171.670 62.900 171.720 ;
        RECT 61.380 171.390 62.900 171.670 ;
        RECT 61.380 171.340 61.760 171.390 ;
        RECT 62.520 171.340 62.900 171.390 ;
        RECT 93.830 171.670 94.210 171.720 ;
        RECT 94.970 171.670 95.350 171.720 ;
        RECT 93.830 171.390 95.350 171.670 ;
        RECT 93.830 171.340 94.210 171.390 ;
        RECT 94.970 171.340 95.350 171.390 ;
        RECT 25.200 170.340 25.580 170.720 ;
        RECT 29.120 170.340 29.500 170.720 ;
        RECT 31.920 170.060 34.160 170.440 ;
        RECT 64.370 170.060 66.610 170.440 ;
        RECT 62.520 169.500 63.040 169.880 ;
        RECT 94.970 169.500 95.490 169.880 ;
        RECT 97.415 168.840 97.795 169.220 ;
        RECT 99.455 168.840 99.835 169.220 ;
        RECT 101.240 168.840 101.620 169.220 ;
        RECT 25.200 167.340 25.580 167.720 ;
        RECT 29.120 167.340 29.500 167.720 ;
        RECT 25.200 164.340 25.580 164.720 ;
        RECT 97.415 162.840 97.795 163.220 ;
        RECT 99.455 162.840 99.835 163.220 ;
        RECT 101.240 162.840 101.620 163.220 ;
        RECT 25.200 161.340 25.580 161.720 ;
        RECT 29.120 161.340 29.500 161.720 ;
        RECT 62.020 160.935 62.900 161.315 ;
        RECT 94.470 160.935 95.350 161.315 ;
        RECT 31.920 160.375 34.160 160.755 ;
        RECT 64.370 160.375 66.610 160.755 ;
        RECT 97.415 159.840 97.795 160.220 ;
        RECT 99.455 159.840 99.835 160.220 ;
        RECT 101.240 159.840 101.620 160.220 ;
        RECT 60.740 159.425 61.120 159.475 ;
        RECT 62.520 159.425 62.900 159.475 ;
        RECT 60.740 159.145 62.900 159.425 ;
        RECT 60.740 159.095 61.120 159.145 ;
        RECT 62.520 159.095 62.900 159.145 ;
        RECT 93.190 159.425 93.570 159.475 ;
        RECT 94.970 159.425 95.350 159.475 ;
        RECT 93.190 159.145 95.350 159.425 ;
        RECT 93.190 159.095 93.570 159.145 ;
        RECT 94.970 159.095 95.350 159.145 ;
        RECT 25.200 158.340 25.580 158.720 ;
        RECT 29.120 158.340 29.500 158.720 ;
        RECT 31.920 158.535 34.160 158.915 ;
        RECT 64.370 158.535 66.610 158.915 ;
        RECT 59.460 157.580 59.840 157.630 ;
        RECT 62.520 157.580 62.900 157.630 ;
        RECT 59.460 157.300 62.900 157.580 ;
        RECT 59.460 157.250 59.840 157.300 ;
        RECT 62.520 157.250 62.900 157.300 ;
        RECT 91.910 157.580 92.290 157.630 ;
        RECT 94.970 157.580 95.350 157.630 ;
        RECT 91.910 157.300 95.350 157.580 ;
        RECT 91.910 157.250 92.290 157.300 ;
        RECT 94.970 157.250 95.350 157.300 ;
        RECT 31.920 156.690 34.160 157.070 ;
        RECT 64.370 156.690 66.610 157.070 ;
        RECT 97.415 156.840 97.795 157.220 ;
        RECT 99.455 156.840 99.835 157.220 ;
        RECT 101.240 156.840 101.620 157.220 ;
        RECT 31.925 155.930 34.165 156.310 ;
        RECT 64.375 155.930 66.615 156.310 ;
        RECT 25.200 155.340 25.580 155.720 ;
        RECT 29.120 155.340 29.500 155.720 ;
        RECT 58.180 154.940 58.560 154.990 ;
        RECT 62.520 154.940 62.900 154.990 ;
        RECT 58.180 154.660 62.900 154.940 ;
        RECT 58.180 154.610 58.560 154.660 ;
        RECT 62.520 154.610 62.900 154.660 ;
        RECT 90.630 154.940 91.010 154.990 ;
        RECT 94.970 154.940 95.350 154.990 ;
        RECT 90.630 154.660 95.350 154.940 ;
        RECT 90.630 154.610 91.010 154.660 ;
        RECT 94.970 154.610 95.350 154.660 ;
        RECT 31.920 154.050 34.160 154.430 ;
        RECT 64.370 154.050 66.610 154.430 ;
        RECT 97.415 153.840 97.795 154.220 ;
        RECT 99.455 153.840 99.835 154.220 ;
        RECT 101.240 153.840 101.620 154.220 ;
        RECT 56.900 153.100 57.280 153.150 ;
        RECT 62.520 153.100 62.900 153.150 ;
        RECT 56.900 152.820 62.900 153.100 ;
        RECT 56.900 152.770 57.280 152.820 ;
        RECT 62.520 152.770 62.900 152.820 ;
        RECT 89.350 153.100 89.730 153.150 ;
        RECT 94.970 153.100 95.350 153.150 ;
        RECT 89.350 152.820 95.350 153.100 ;
        RECT 89.350 152.770 89.730 152.820 ;
        RECT 94.970 152.770 95.350 152.820 ;
        RECT 25.200 152.340 25.580 152.720 ;
        RECT 29.120 152.340 29.500 152.720 ;
        RECT 31.920 152.210 34.160 152.590 ;
        RECT 64.370 152.210 66.610 152.590 ;
        RECT 55.620 151.255 56.000 151.305 ;
        RECT 62.520 151.255 62.900 151.305 ;
        RECT 55.620 150.975 62.900 151.255 ;
        RECT 55.620 150.925 56.000 150.975 ;
        RECT 62.520 150.925 62.900 150.975 ;
        RECT 88.070 151.255 88.450 151.305 ;
        RECT 94.970 151.255 95.350 151.305 ;
        RECT 88.070 150.975 95.350 151.255 ;
        RECT 88.070 150.925 88.450 150.975 ;
        RECT 94.970 150.925 95.350 150.975 ;
        RECT 97.415 150.840 97.795 151.220 ;
        RECT 99.455 150.840 99.835 151.220 ;
        RECT 101.240 150.840 101.620 151.220 ;
        RECT 31.920 150.365 34.160 150.745 ;
        RECT 64.370 150.365 66.610 150.745 ;
        RECT 25.200 149.340 25.580 149.720 ;
        RECT 29.120 149.340 29.500 149.720 ;
        RECT 31.925 149.605 34.165 149.985 ;
        RECT 64.375 149.605 66.615 149.985 ;
        RECT 54.340 148.615 54.720 148.665 ;
        RECT 62.520 148.615 62.900 148.665 ;
        RECT 54.340 148.335 62.900 148.615 ;
        RECT 54.340 148.285 54.720 148.335 ;
        RECT 62.520 148.285 62.900 148.335 ;
        RECT 86.790 148.615 87.170 148.665 ;
        RECT 94.970 148.615 95.350 148.665 ;
        RECT 86.790 148.335 95.350 148.615 ;
        RECT 86.790 148.285 87.170 148.335 ;
        RECT 94.970 148.285 95.350 148.335 ;
        RECT 31.920 147.725 34.160 148.105 ;
        RECT 64.370 147.725 66.610 148.105 ;
        RECT 97.415 147.840 97.795 148.220 ;
        RECT 99.455 147.840 99.835 148.220 ;
        RECT 101.240 147.840 101.620 148.220 ;
        RECT 53.060 146.775 53.440 146.825 ;
        RECT 62.520 146.775 62.900 146.825 ;
        RECT 25.200 146.340 25.580 146.720 ;
        RECT 29.120 146.340 29.500 146.720 ;
        RECT 53.060 146.495 62.900 146.775 ;
        RECT 53.060 146.445 53.440 146.495 ;
        RECT 62.520 146.445 62.900 146.495 ;
        RECT 85.510 146.775 85.890 146.825 ;
        RECT 94.970 146.775 95.350 146.825 ;
        RECT 85.510 146.495 95.350 146.775 ;
        RECT 85.510 146.445 85.890 146.495 ;
        RECT 94.970 146.445 95.350 146.495 ;
        RECT 31.920 145.885 34.160 146.265 ;
        RECT 64.370 145.885 66.610 146.265 ;
        RECT 31.920 145.165 34.160 145.545 ;
        RECT 64.370 145.165 66.610 145.545 ;
        RECT 53.700 144.935 54.080 144.985 ;
        RECT 62.520 144.935 62.900 144.985 ;
        RECT 53.700 144.655 62.900 144.935 ;
        RECT 53.700 144.605 54.080 144.655 ;
        RECT 62.520 144.605 62.900 144.655 ;
        RECT 86.150 144.935 86.530 144.985 ;
        RECT 94.970 144.935 95.350 144.985 ;
        RECT 86.150 144.655 95.350 144.935 ;
        RECT 86.150 144.605 86.530 144.655 ;
        RECT 94.970 144.605 95.350 144.655 ;
        RECT 25.200 142.955 25.580 143.335 ;
        RECT 29.120 142.955 29.500 143.335 ;
        RECT 31.920 143.325 34.160 143.705 ;
        RECT 64.370 143.325 66.610 143.705 ;
        RECT 54.980 143.095 55.360 143.145 ;
        RECT 62.520 143.095 62.900 143.145 ;
        RECT 54.980 142.815 62.900 143.095 ;
        RECT 54.980 142.765 55.360 142.815 ;
        RECT 62.520 142.765 62.900 142.815 ;
        RECT 87.430 143.095 87.810 143.145 ;
        RECT 94.970 143.095 95.350 143.145 ;
        RECT 87.430 142.815 95.350 143.095 ;
        RECT 87.430 142.765 87.810 142.815 ;
        RECT 94.970 142.765 95.350 142.815 ;
        RECT 31.925 141.440 34.165 141.820 ;
        RECT 64.375 141.440 66.615 141.820 ;
        RECT 97.415 141.455 97.795 141.835 ;
        RECT 99.455 141.455 99.835 141.835 ;
        RECT 101.240 141.455 101.620 141.835 ;
        RECT 31.920 140.680 34.160 141.060 ;
        RECT 64.370 140.680 66.610 141.060 ;
        RECT 56.260 140.450 56.640 140.500 ;
        RECT 62.520 140.450 62.900 140.500 ;
        RECT 25.200 139.955 25.580 140.335 ;
        RECT 29.120 139.955 29.500 140.335 ;
        RECT 56.260 140.170 62.900 140.450 ;
        RECT 56.260 140.120 56.640 140.170 ;
        RECT 62.520 140.120 62.900 140.170 ;
        RECT 88.710 140.450 89.090 140.500 ;
        RECT 94.970 140.450 95.350 140.500 ;
        RECT 88.710 140.170 95.350 140.450 ;
        RECT 88.710 140.120 89.090 140.170 ;
        RECT 94.970 140.120 95.350 140.170 ;
        RECT 31.920 138.840 34.160 139.220 ;
        RECT 64.370 138.840 66.610 139.220 ;
        RECT 57.540 138.610 57.920 138.660 ;
        RECT 62.520 138.610 62.900 138.660 ;
        RECT 57.540 138.330 62.900 138.610 ;
        RECT 57.540 138.280 57.920 138.330 ;
        RECT 62.520 138.280 62.900 138.330 ;
        RECT 89.990 138.610 90.370 138.660 ;
        RECT 94.970 138.610 95.350 138.660 ;
        RECT 89.990 138.330 95.350 138.610 ;
        RECT 97.415 138.455 97.795 138.835 ;
        RECT 99.455 138.455 99.835 138.835 ;
        RECT 101.240 138.455 101.620 138.835 ;
        RECT 89.990 138.280 90.370 138.330 ;
        RECT 94.970 138.280 95.350 138.330 ;
        RECT 25.200 136.955 25.580 137.335 ;
        RECT 29.120 136.955 29.500 137.335 ;
        RECT 31.920 137.000 34.160 137.380 ;
        RECT 64.370 137.000 66.610 137.380 ;
        RECT 58.820 136.770 59.200 136.820 ;
        RECT 62.520 136.770 62.900 136.820 ;
        RECT 58.820 136.490 62.900 136.770 ;
        RECT 58.820 136.440 59.200 136.490 ;
        RECT 62.520 136.440 62.900 136.490 ;
        RECT 91.270 136.770 91.650 136.820 ;
        RECT 94.970 136.770 95.350 136.820 ;
        RECT 91.270 136.490 95.350 136.770 ;
        RECT 91.270 136.440 91.650 136.490 ;
        RECT 94.970 136.440 95.350 136.490 ;
        RECT 31.925 135.115 34.165 135.495 ;
        RECT 64.375 135.115 66.615 135.495 ;
        RECT 97.415 135.455 97.795 135.835 ;
        RECT 99.455 135.455 99.835 135.835 ;
        RECT 101.240 135.455 101.620 135.835 ;
        RECT 31.920 134.355 34.160 134.735 ;
        RECT 64.370 134.355 66.610 134.735 ;
        RECT 25.200 133.955 25.580 134.335 ;
        RECT 29.120 133.955 29.500 134.335 ;
        RECT 60.100 134.125 60.480 134.175 ;
        RECT 62.520 134.125 62.900 134.175 ;
        RECT 60.100 133.845 62.900 134.125 ;
        RECT 60.100 133.795 60.480 133.845 ;
        RECT 62.520 133.795 62.900 133.845 ;
        RECT 92.550 134.125 92.930 134.175 ;
        RECT 94.970 134.125 95.350 134.175 ;
        RECT 92.550 133.845 95.350 134.125 ;
        RECT 92.550 133.795 92.930 133.845 ;
        RECT 94.970 133.795 95.350 133.845 ;
        RECT 31.920 132.515 34.160 132.895 ;
        RECT 64.370 132.515 66.610 132.895 ;
        RECT 97.415 132.455 97.795 132.835 ;
        RECT 99.455 132.455 99.835 132.835 ;
        RECT 101.240 132.455 101.620 132.835 ;
        RECT 61.380 132.285 61.760 132.335 ;
        RECT 62.520 132.285 62.900 132.335 ;
        RECT 61.380 132.005 62.900 132.285 ;
        RECT 61.380 131.955 61.760 132.005 ;
        RECT 62.520 131.955 62.900 132.005 ;
        RECT 93.830 132.285 94.210 132.335 ;
        RECT 94.970 132.285 95.350 132.335 ;
        RECT 93.830 132.005 95.350 132.285 ;
        RECT 93.830 131.955 94.210 132.005 ;
        RECT 94.970 131.955 95.350 132.005 ;
        RECT 25.200 130.955 25.580 131.335 ;
        RECT 29.120 130.955 29.500 131.335 ;
        RECT 31.920 130.675 34.160 131.055 ;
        RECT 64.370 130.675 66.610 131.055 ;
        RECT 62.520 130.115 63.040 130.495 ;
        RECT 94.970 130.115 95.490 130.495 ;
        RECT 97.415 129.455 97.795 129.835 ;
        RECT 99.455 129.455 99.835 129.835 ;
        RECT 101.240 129.455 101.620 129.835 ;
        RECT 25.200 127.955 25.580 128.335 ;
        RECT 29.120 127.955 29.500 128.335 ;
        RECT 25.200 124.955 25.580 125.335 ;
        RECT 97.415 123.455 97.795 123.835 ;
        RECT 99.455 123.455 99.835 123.835 ;
        RECT 101.240 123.455 101.620 123.835 ;
        RECT 25.200 121.955 25.580 122.335 ;
        RECT 29.120 121.955 29.500 122.335 ;
        RECT 62.020 121.550 62.900 121.930 ;
        RECT 94.470 121.550 95.350 121.930 ;
        RECT 31.920 120.990 34.160 121.370 ;
        RECT 64.370 120.990 66.610 121.370 ;
        RECT 97.415 120.455 97.795 120.835 ;
        RECT 99.455 120.455 99.835 120.835 ;
        RECT 101.240 120.455 101.620 120.835 ;
        RECT 60.740 120.040 61.120 120.090 ;
        RECT 62.520 120.040 62.900 120.090 ;
        RECT 60.740 119.760 62.900 120.040 ;
        RECT 60.740 119.710 61.120 119.760 ;
        RECT 62.520 119.710 62.900 119.760 ;
        RECT 93.190 120.040 93.570 120.090 ;
        RECT 94.970 120.040 95.350 120.090 ;
        RECT 93.190 119.760 95.350 120.040 ;
        RECT 93.190 119.710 93.570 119.760 ;
        RECT 94.970 119.710 95.350 119.760 ;
        RECT 25.200 118.955 25.580 119.335 ;
        RECT 29.120 118.955 29.500 119.335 ;
        RECT 31.920 119.150 34.160 119.530 ;
        RECT 64.370 119.150 66.610 119.530 ;
        RECT 59.460 118.195 59.840 118.245 ;
        RECT 62.520 118.195 62.900 118.245 ;
        RECT 59.460 117.915 62.900 118.195 ;
        RECT 59.460 117.865 59.840 117.915 ;
        RECT 62.520 117.865 62.900 117.915 ;
        RECT 91.910 118.195 92.290 118.245 ;
        RECT 94.970 118.195 95.350 118.245 ;
        RECT 91.910 117.915 95.350 118.195 ;
        RECT 91.910 117.865 92.290 117.915 ;
        RECT 94.970 117.865 95.350 117.915 ;
        RECT 31.920 117.305 34.160 117.685 ;
        RECT 64.370 117.305 66.610 117.685 ;
        RECT 97.415 117.455 97.795 117.835 ;
        RECT 99.455 117.455 99.835 117.835 ;
        RECT 101.240 117.455 101.620 117.835 ;
        RECT 31.925 116.545 34.165 116.925 ;
        RECT 64.375 116.545 66.615 116.925 ;
        RECT 25.200 115.955 25.580 116.335 ;
        RECT 29.120 115.955 29.500 116.335 ;
        RECT 58.180 115.555 58.560 115.605 ;
        RECT 62.520 115.555 62.900 115.605 ;
        RECT 58.180 115.275 62.900 115.555 ;
        RECT 58.180 115.225 58.560 115.275 ;
        RECT 62.520 115.225 62.900 115.275 ;
        RECT 90.630 115.555 91.010 115.605 ;
        RECT 94.970 115.555 95.350 115.605 ;
        RECT 90.630 115.275 95.350 115.555 ;
        RECT 90.630 115.225 91.010 115.275 ;
        RECT 94.970 115.225 95.350 115.275 ;
        RECT 31.920 114.665 34.160 115.045 ;
        RECT 64.370 114.665 66.610 115.045 ;
        RECT 97.415 114.455 97.795 114.835 ;
        RECT 99.455 114.455 99.835 114.835 ;
        RECT 101.240 114.455 101.620 114.835 ;
        RECT 56.900 113.715 57.280 113.765 ;
        RECT 62.520 113.715 62.900 113.765 ;
        RECT 56.900 113.435 62.900 113.715 ;
        RECT 56.900 113.385 57.280 113.435 ;
        RECT 62.520 113.385 62.900 113.435 ;
        RECT 89.350 113.715 89.730 113.765 ;
        RECT 94.970 113.715 95.350 113.765 ;
        RECT 89.350 113.435 95.350 113.715 ;
        RECT 89.350 113.385 89.730 113.435 ;
        RECT 94.970 113.385 95.350 113.435 ;
        RECT 25.200 112.955 25.580 113.335 ;
        RECT 29.120 112.955 29.500 113.335 ;
        RECT 31.920 112.825 34.160 113.205 ;
        RECT 64.370 112.825 66.610 113.205 ;
        RECT 55.620 111.870 56.000 111.920 ;
        RECT 62.520 111.870 62.900 111.920 ;
        RECT 55.620 111.590 62.900 111.870 ;
        RECT 55.620 111.540 56.000 111.590 ;
        RECT 62.520 111.540 62.900 111.590 ;
        RECT 88.070 111.870 88.450 111.920 ;
        RECT 94.970 111.870 95.350 111.920 ;
        RECT 88.070 111.590 95.350 111.870 ;
        RECT 88.070 111.540 88.450 111.590 ;
        RECT 94.970 111.540 95.350 111.590 ;
        RECT 97.415 111.455 97.795 111.835 ;
        RECT 99.455 111.455 99.835 111.835 ;
        RECT 101.240 111.455 101.620 111.835 ;
        RECT 31.920 110.980 34.160 111.360 ;
        RECT 64.370 110.980 66.610 111.360 ;
        RECT 25.200 109.955 25.580 110.335 ;
        RECT 29.120 109.955 29.500 110.335 ;
        RECT 31.925 110.220 34.165 110.600 ;
        RECT 64.375 110.220 66.615 110.600 ;
        RECT 54.340 109.230 54.720 109.280 ;
        RECT 62.520 109.230 62.900 109.280 ;
        RECT 54.340 108.950 62.900 109.230 ;
        RECT 54.340 108.900 54.720 108.950 ;
        RECT 62.520 108.900 62.900 108.950 ;
        RECT 86.790 109.230 87.170 109.280 ;
        RECT 94.970 109.230 95.350 109.280 ;
        RECT 86.790 108.950 95.350 109.230 ;
        RECT 86.790 108.900 87.170 108.950 ;
        RECT 94.970 108.900 95.350 108.950 ;
        RECT 31.920 108.340 34.160 108.720 ;
        RECT 64.370 108.340 66.610 108.720 ;
        RECT 97.415 108.455 97.795 108.835 ;
        RECT 99.455 108.455 99.835 108.835 ;
        RECT 101.240 108.455 101.620 108.835 ;
        RECT 53.060 107.390 53.440 107.440 ;
        RECT 62.520 107.390 62.900 107.440 ;
        RECT 25.200 106.955 25.580 107.335 ;
        RECT 29.120 106.955 29.500 107.335 ;
        RECT 53.060 107.110 62.900 107.390 ;
        RECT 53.060 107.060 53.440 107.110 ;
        RECT 62.520 107.060 62.900 107.110 ;
        RECT 85.510 107.390 85.890 107.440 ;
        RECT 94.970 107.390 95.350 107.440 ;
        RECT 85.510 107.110 95.350 107.390 ;
        RECT 85.510 107.060 85.890 107.110 ;
        RECT 94.970 107.060 95.350 107.110 ;
        RECT 31.920 106.500 34.160 106.880 ;
        RECT 64.370 106.500 66.610 106.880 ;
        RECT 31.920 105.780 34.160 106.160 ;
        RECT 64.370 105.780 66.610 106.160 ;
        RECT 53.700 105.550 54.080 105.600 ;
        RECT 62.520 105.550 62.900 105.600 ;
        RECT 53.700 105.270 62.900 105.550 ;
        RECT 53.700 105.220 54.080 105.270 ;
        RECT 62.520 105.220 62.900 105.270 ;
        RECT 86.150 105.550 86.530 105.600 ;
        RECT 94.970 105.550 95.350 105.600 ;
        RECT 86.150 105.270 95.350 105.550 ;
        RECT 86.150 105.220 86.530 105.270 ;
        RECT 94.970 105.220 95.350 105.270 ;
        RECT 25.200 103.570 25.580 103.950 ;
        RECT 29.120 103.570 29.500 103.950 ;
        RECT 31.920 103.940 34.160 104.320 ;
        RECT 64.370 103.940 66.610 104.320 ;
        RECT 54.980 103.710 55.360 103.760 ;
        RECT 62.520 103.710 62.900 103.760 ;
        RECT 54.980 103.430 62.900 103.710 ;
        RECT 54.980 103.380 55.360 103.430 ;
        RECT 62.520 103.380 62.900 103.430 ;
        RECT 87.430 103.710 87.810 103.760 ;
        RECT 94.970 103.710 95.350 103.760 ;
        RECT 87.430 103.430 95.350 103.710 ;
        RECT 87.430 103.380 87.810 103.430 ;
        RECT 94.970 103.380 95.350 103.430 ;
        RECT 31.925 102.055 34.165 102.435 ;
        RECT 64.375 102.055 66.615 102.435 ;
        RECT 97.415 102.070 97.795 102.450 ;
        RECT 99.455 102.070 99.835 102.450 ;
        RECT 101.240 102.070 101.620 102.450 ;
        RECT 31.920 101.295 34.160 101.675 ;
        RECT 64.370 101.295 66.610 101.675 ;
        RECT 56.260 101.065 56.640 101.115 ;
        RECT 62.520 101.065 62.900 101.115 ;
        RECT 25.200 100.570 25.580 100.950 ;
        RECT 29.120 100.570 29.500 100.950 ;
        RECT 56.260 100.785 62.900 101.065 ;
        RECT 56.260 100.735 56.640 100.785 ;
        RECT 62.520 100.735 62.900 100.785 ;
        RECT 88.710 101.065 89.090 101.115 ;
        RECT 94.970 101.065 95.350 101.115 ;
        RECT 88.710 100.785 95.350 101.065 ;
        RECT 88.710 100.735 89.090 100.785 ;
        RECT 94.970 100.735 95.350 100.785 ;
        RECT 31.920 99.455 34.160 99.835 ;
        RECT 64.370 99.455 66.610 99.835 ;
        RECT 57.540 99.225 57.920 99.275 ;
        RECT 62.520 99.225 62.900 99.275 ;
        RECT 57.540 98.945 62.900 99.225 ;
        RECT 57.540 98.895 57.920 98.945 ;
        RECT 62.520 98.895 62.900 98.945 ;
        RECT 89.990 99.225 90.370 99.275 ;
        RECT 94.970 99.225 95.350 99.275 ;
        RECT 89.990 98.945 95.350 99.225 ;
        RECT 97.415 99.070 97.795 99.450 ;
        RECT 99.455 99.070 99.835 99.450 ;
        RECT 101.240 99.070 101.620 99.450 ;
        RECT 89.990 98.895 90.370 98.945 ;
        RECT 94.970 98.895 95.350 98.945 ;
        RECT 25.200 97.570 25.580 97.950 ;
        RECT 29.120 97.570 29.500 97.950 ;
        RECT 31.920 97.615 34.160 97.995 ;
        RECT 64.370 97.615 66.610 97.995 ;
        RECT 58.820 97.385 59.200 97.435 ;
        RECT 62.520 97.385 62.900 97.435 ;
        RECT 58.820 97.105 62.900 97.385 ;
        RECT 58.820 97.055 59.200 97.105 ;
        RECT 62.520 97.055 62.900 97.105 ;
        RECT 91.270 97.385 91.650 97.435 ;
        RECT 94.970 97.385 95.350 97.435 ;
        RECT 91.270 97.105 95.350 97.385 ;
        RECT 91.270 97.055 91.650 97.105 ;
        RECT 94.970 97.055 95.350 97.105 ;
        RECT 31.925 95.730 34.165 96.110 ;
        RECT 64.375 95.730 66.615 96.110 ;
        RECT 97.415 96.070 97.795 96.450 ;
        RECT 99.455 96.070 99.835 96.450 ;
        RECT 101.240 96.070 101.620 96.450 ;
        RECT 31.920 94.970 34.160 95.350 ;
        RECT 64.370 94.970 66.610 95.350 ;
        RECT 25.200 94.570 25.580 94.950 ;
        RECT 29.120 94.570 29.500 94.950 ;
        RECT 60.100 94.740 60.480 94.790 ;
        RECT 62.520 94.740 62.900 94.790 ;
        RECT 60.100 94.460 62.900 94.740 ;
        RECT 60.100 94.410 60.480 94.460 ;
        RECT 62.520 94.410 62.900 94.460 ;
        RECT 92.550 94.740 92.930 94.790 ;
        RECT 94.970 94.740 95.350 94.790 ;
        RECT 92.550 94.460 95.350 94.740 ;
        RECT 92.550 94.410 92.930 94.460 ;
        RECT 94.970 94.410 95.350 94.460 ;
        RECT 31.920 93.130 34.160 93.510 ;
        RECT 64.370 93.130 66.610 93.510 ;
        RECT 97.415 93.070 97.795 93.450 ;
        RECT 99.455 93.070 99.835 93.450 ;
        RECT 101.240 93.070 101.620 93.450 ;
        RECT 61.380 92.900 61.760 92.950 ;
        RECT 62.520 92.900 62.900 92.950 ;
        RECT 61.380 92.620 62.900 92.900 ;
        RECT 61.380 92.570 61.760 92.620 ;
        RECT 62.520 92.570 62.900 92.620 ;
        RECT 93.830 92.900 94.210 92.950 ;
        RECT 94.970 92.900 95.350 92.950 ;
        RECT 93.830 92.620 95.350 92.900 ;
        RECT 93.830 92.570 94.210 92.620 ;
        RECT 94.970 92.570 95.350 92.620 ;
        RECT 25.200 91.570 25.580 91.950 ;
        RECT 29.120 91.570 29.500 91.950 ;
        RECT 31.920 91.290 34.160 91.670 ;
        RECT 64.370 91.290 66.610 91.670 ;
        RECT 62.520 90.730 63.040 91.110 ;
        RECT 94.970 90.730 95.490 91.110 ;
        RECT 97.415 90.070 97.795 90.450 ;
        RECT 99.455 90.070 99.835 90.450 ;
        RECT 101.240 90.070 101.620 90.450 ;
        RECT 25.200 88.570 25.580 88.950 ;
        RECT 29.120 88.570 29.500 88.950 ;
        RECT 25.200 85.570 25.580 85.950 ;
        RECT 97.415 84.070 97.795 84.450 ;
        RECT 99.455 84.070 99.835 84.450 ;
        RECT 101.240 84.070 101.620 84.450 ;
        RECT 25.200 82.570 25.580 82.950 ;
        RECT 29.120 82.570 29.500 82.950 ;
        RECT 62.020 82.165 62.900 82.545 ;
        RECT 94.470 82.165 95.350 82.545 ;
        RECT 31.920 81.605 34.160 81.985 ;
        RECT 64.370 81.605 66.610 81.985 ;
        RECT 97.415 81.070 97.795 81.450 ;
        RECT 99.455 81.070 99.835 81.450 ;
        RECT 101.240 81.070 101.620 81.450 ;
        RECT 60.740 80.655 61.120 80.705 ;
        RECT 62.520 80.655 62.900 80.705 ;
        RECT 60.740 80.375 62.900 80.655 ;
        RECT 60.740 80.325 61.120 80.375 ;
        RECT 62.520 80.325 62.900 80.375 ;
        RECT 93.190 80.655 93.570 80.705 ;
        RECT 94.970 80.655 95.350 80.705 ;
        RECT 93.190 80.375 95.350 80.655 ;
        RECT 93.190 80.325 93.570 80.375 ;
        RECT 94.970 80.325 95.350 80.375 ;
        RECT 25.200 79.570 25.580 79.950 ;
        RECT 29.120 79.570 29.500 79.950 ;
        RECT 31.920 79.765 34.160 80.145 ;
        RECT 64.370 79.765 66.610 80.145 ;
        RECT 59.460 78.810 59.840 78.860 ;
        RECT 62.520 78.810 62.900 78.860 ;
        RECT 59.460 78.530 62.900 78.810 ;
        RECT 59.460 78.480 59.840 78.530 ;
        RECT 62.520 78.480 62.900 78.530 ;
        RECT 91.910 78.810 92.290 78.860 ;
        RECT 94.970 78.810 95.350 78.860 ;
        RECT 91.910 78.530 95.350 78.810 ;
        RECT 91.910 78.480 92.290 78.530 ;
        RECT 94.970 78.480 95.350 78.530 ;
        RECT 31.920 77.920 34.160 78.300 ;
        RECT 64.370 77.920 66.610 78.300 ;
        RECT 97.415 78.070 97.795 78.450 ;
        RECT 99.455 78.070 99.835 78.450 ;
        RECT 101.240 78.070 101.620 78.450 ;
        RECT 31.925 77.160 34.165 77.540 ;
        RECT 64.375 77.160 66.615 77.540 ;
        RECT 25.200 76.570 25.580 76.950 ;
        RECT 29.120 76.570 29.500 76.950 ;
        RECT 58.180 76.170 58.560 76.220 ;
        RECT 62.520 76.170 62.900 76.220 ;
        RECT 58.180 75.890 62.900 76.170 ;
        RECT 58.180 75.840 58.560 75.890 ;
        RECT 62.520 75.840 62.900 75.890 ;
        RECT 90.630 76.170 91.010 76.220 ;
        RECT 94.970 76.170 95.350 76.220 ;
        RECT 90.630 75.890 95.350 76.170 ;
        RECT 90.630 75.840 91.010 75.890 ;
        RECT 94.970 75.840 95.350 75.890 ;
        RECT 31.920 75.280 34.160 75.660 ;
        RECT 64.370 75.280 66.610 75.660 ;
        RECT 97.415 75.070 97.795 75.450 ;
        RECT 99.455 75.070 99.835 75.450 ;
        RECT 101.240 75.070 101.620 75.450 ;
        RECT 56.900 74.330 57.280 74.380 ;
        RECT 62.520 74.330 62.900 74.380 ;
        RECT 56.900 74.050 62.900 74.330 ;
        RECT 56.900 74.000 57.280 74.050 ;
        RECT 62.520 74.000 62.900 74.050 ;
        RECT 89.350 74.330 89.730 74.380 ;
        RECT 94.970 74.330 95.350 74.380 ;
        RECT 89.350 74.050 95.350 74.330 ;
        RECT 89.350 74.000 89.730 74.050 ;
        RECT 94.970 74.000 95.350 74.050 ;
        RECT 25.200 73.570 25.580 73.950 ;
        RECT 29.120 73.570 29.500 73.950 ;
        RECT 31.920 73.440 34.160 73.820 ;
        RECT 64.370 73.440 66.610 73.820 ;
        RECT 55.620 72.485 56.000 72.535 ;
        RECT 62.520 72.485 62.900 72.535 ;
        RECT 55.620 72.205 62.900 72.485 ;
        RECT 55.620 72.155 56.000 72.205 ;
        RECT 62.520 72.155 62.900 72.205 ;
        RECT 88.070 72.485 88.450 72.535 ;
        RECT 94.970 72.485 95.350 72.535 ;
        RECT 88.070 72.205 95.350 72.485 ;
        RECT 88.070 72.155 88.450 72.205 ;
        RECT 94.970 72.155 95.350 72.205 ;
        RECT 97.415 72.070 97.795 72.450 ;
        RECT 99.455 72.070 99.835 72.450 ;
        RECT 101.240 72.070 101.620 72.450 ;
        RECT 31.920 71.595 34.160 71.975 ;
        RECT 64.370 71.595 66.610 71.975 ;
        RECT 25.200 70.570 25.580 70.950 ;
        RECT 29.120 70.570 29.500 70.950 ;
        RECT 31.925 70.835 34.165 71.215 ;
        RECT 64.375 70.835 66.615 71.215 ;
        RECT 54.340 69.845 54.720 69.895 ;
        RECT 62.520 69.845 62.900 69.895 ;
        RECT 54.340 69.565 62.900 69.845 ;
        RECT 54.340 69.515 54.720 69.565 ;
        RECT 62.520 69.515 62.900 69.565 ;
        RECT 86.790 69.845 87.170 69.895 ;
        RECT 94.970 69.845 95.350 69.895 ;
        RECT 86.790 69.565 95.350 69.845 ;
        RECT 86.790 69.515 87.170 69.565 ;
        RECT 94.970 69.515 95.350 69.565 ;
        RECT 31.920 68.955 34.160 69.335 ;
        RECT 64.370 68.955 66.610 69.335 ;
        RECT 97.415 69.070 97.795 69.450 ;
        RECT 99.455 69.070 99.835 69.450 ;
        RECT 101.240 69.070 101.620 69.450 ;
        RECT 53.060 68.005 53.440 68.055 ;
        RECT 62.520 68.005 62.900 68.055 ;
        RECT 25.200 67.570 25.580 67.950 ;
        RECT 29.120 67.570 29.500 67.950 ;
        RECT 53.060 67.725 62.900 68.005 ;
        RECT 53.060 67.675 53.440 67.725 ;
        RECT 62.520 67.675 62.900 67.725 ;
        RECT 85.510 68.005 85.890 68.055 ;
        RECT 94.970 68.005 95.350 68.055 ;
        RECT 85.510 67.725 95.350 68.005 ;
        RECT 85.510 67.675 85.890 67.725 ;
        RECT 94.970 67.675 95.350 67.725 ;
        RECT 31.920 67.115 34.160 67.495 ;
        RECT 64.370 67.115 66.610 67.495 ;
  END
END efuse_array_32x8
END LIBRARY

