VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_array_16x1
  CLASS BLOCK ;
  FOREIGN efuse_array_16x1 ;
  ORIGIN -24.960 -66.885 ;
  SIZE 44.480 BY 40.130 ;
  PIN COL_PROG_N[0]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 64.400 106.315 67.960 106.615 ;
    END
  END COL_PROG_N[0]
  PIN OUT[0]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 77.995 28.780 78.325 ;
    END
  END OUT[0]
  PIN PRESET_N
    ANTENNAGATEAREA 1.220000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.970 86.725 26.250 107.015 ;
        RECT 25.970 86.345 26.330 86.725 ;
        RECT 25.970 66.885 26.250 86.345 ;
    END
  END PRESET_N
  PIN SENSE
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.615 85.540 26.895 107.015 ;
        RECT 26.615 85.160 28.040 85.540 ;
        RECT 26.615 66.885 26.895 85.160 ;
    END
  END SENSE
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 31.430 66.885 34.430 107.015 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 28.670 66.885 29.670 107.015 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 25.030 66.885 26.030 107.015 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 64.950 66.885 69.200 107.015 ;
    END
  END VDD
  PIN BIT_SEL[0]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 62.700 91.110 62.980 106.390 ;
        RECT 62.660 90.730 63.040 91.110 ;
        RECT 62.700 66.885 62.980 90.730 ;
    END
  END BIT_SEL[0]
  PIN BIT_SEL[1]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 62.060 82.545 62.340 106.390 ;
        RECT 62.020 82.165 62.400 82.545 ;
        RECT 62.060 66.885 62.340 82.165 ;
    END
  END BIT_SEL[1]
  PIN BIT_SEL[2]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 61.420 92.950 61.700 106.390 ;
        RECT 61.380 92.570 61.760 92.950 ;
        RECT 61.420 66.885 61.700 92.570 ;
    END
  END BIT_SEL[2]
  PIN BIT_SEL[3]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 60.780 80.705 61.060 106.390 ;
        RECT 60.740 80.325 61.120 80.705 ;
        RECT 60.780 66.885 61.060 80.325 ;
    END
  END BIT_SEL[3]
  PIN BIT_SEL[4]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 60.140 94.790 60.420 106.390 ;
        RECT 60.100 94.410 60.480 94.790 ;
        RECT 60.140 66.885 60.420 94.410 ;
    END
  END BIT_SEL[4]
  PIN BIT_SEL[5]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 59.500 78.860 59.780 106.390 ;
        RECT 59.460 78.480 59.840 78.860 ;
        RECT 59.500 66.885 59.780 78.480 ;
    END
  END BIT_SEL[5]
  PIN BIT_SEL[6]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 58.860 97.435 59.140 106.390 ;
        RECT 58.820 97.055 59.200 97.435 ;
        RECT 58.860 66.885 59.140 97.055 ;
    END
  END BIT_SEL[6]
  PIN BIT_SEL[7]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 58.220 76.220 58.500 106.390 ;
        RECT 58.180 75.840 58.560 76.220 ;
        RECT 58.220 66.885 58.500 75.840 ;
    END
  END BIT_SEL[7]
  PIN BIT_SEL[8]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 57.580 99.275 57.860 106.390 ;
        RECT 57.540 98.895 57.920 99.275 ;
        RECT 57.580 66.885 57.860 98.895 ;
    END
  END BIT_SEL[8]
  PIN BIT_SEL[9]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 56.940 74.380 57.220 106.390 ;
        RECT 56.900 74.000 57.280 74.380 ;
        RECT 56.940 66.885 57.220 74.000 ;
    END
  END BIT_SEL[9]
  PIN BIT_SEL[10]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 56.300 101.115 56.580 106.390 ;
        RECT 56.260 100.735 56.640 101.115 ;
        RECT 56.300 66.885 56.580 100.735 ;
    END
  END BIT_SEL[10]
  PIN BIT_SEL[11]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 55.660 72.535 55.940 106.390 ;
        RECT 55.620 72.155 56.000 72.535 ;
        RECT 55.660 66.885 55.940 72.155 ;
    END
  END BIT_SEL[11]
  PIN BIT_SEL[12]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 55.020 103.760 55.300 106.390 ;
        RECT 54.980 103.380 55.360 103.760 ;
        RECT 55.020 66.885 55.300 103.380 ;
    END
  END BIT_SEL[12]
  PIN BIT_SEL[13]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 54.380 69.895 54.660 106.390 ;
        RECT 54.340 69.515 54.720 69.895 ;
        RECT 54.380 66.885 54.660 69.515 ;
    END
  END BIT_SEL[13]
  PIN BIT_SEL[14]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 53.740 105.600 54.020 106.390 ;
        RECT 53.700 105.220 54.080 105.600 ;
        RECT 53.740 66.885 54.020 105.220 ;
    END
  END BIT_SEL[14]
  PIN BIT_SEL[15]
    ANTENNAGATEAREA 18.299999 ;
    PORT
      LAYER Metal4 ;
        RECT 53.100 68.055 53.380 106.390 ;
        RECT 53.060 67.675 53.440 68.055 ;
        RECT 53.100 66.885 53.380 67.675 ;
    END
  END BIT_SEL[15]
  OBS
      LAYER Metal1 ;
        RECT 25.090 88.160 25.690 107.015 ;
        RECT 29.010 88.160 29.610 107.015 ;
        RECT 31.650 105.780 62.170 106.160 ;
        RECT 30.800 105.525 31.420 105.710 ;
        RECT 62.400 105.525 63.020 105.710 ;
        RECT 30.800 105.295 63.020 105.525 ;
        RECT 30.800 105.110 31.420 105.295 ;
        RECT 62.400 105.110 63.020 105.295 ;
        RECT 58.400 105.030 60.020 105.040 ;
        RECT 31.650 104.660 62.170 105.030 ;
        RECT 31.650 103.940 62.170 104.320 ;
        RECT 30.800 103.685 31.420 103.870 ;
        RECT 62.400 103.685 63.020 103.870 ;
        RECT 30.800 103.455 63.020 103.685 ;
        RECT 30.800 103.270 31.420 103.455 ;
        RECT 62.400 103.270 63.020 103.455 ;
        RECT 54.560 103.190 56.180 103.200 ;
        RECT 31.650 102.820 62.170 103.190 ;
        RECT 31.660 102.025 62.160 102.465 ;
        RECT 31.650 101.295 62.170 101.675 ;
        RECT 30.800 101.040 31.420 101.225 ;
        RECT 62.400 101.040 63.020 101.225 ;
        RECT 30.800 100.810 63.020 101.040 ;
        RECT 30.800 100.625 31.420 100.810 ;
        RECT 62.400 100.625 63.020 100.810 ;
        RECT 50.720 100.545 52.340 100.555 ;
        RECT 31.650 100.175 62.170 100.545 ;
        RECT 31.650 99.455 62.170 99.835 ;
        RECT 30.800 99.200 31.420 99.385 ;
        RECT 62.400 99.200 63.020 99.385 ;
        RECT 30.800 98.970 63.020 99.200 ;
        RECT 30.800 98.785 31.420 98.970 ;
        RECT 62.400 98.785 63.020 98.970 ;
        RECT 46.880 98.705 48.500 98.715 ;
        RECT 31.650 98.335 62.170 98.705 ;
        RECT 31.650 97.615 62.170 97.995 ;
        RECT 30.800 97.360 31.420 97.545 ;
        RECT 62.400 97.360 63.020 97.545 ;
        RECT 30.800 97.130 63.020 97.360 ;
        RECT 30.800 96.945 31.420 97.130 ;
        RECT 62.400 96.945 63.020 97.130 ;
        RECT 43.040 96.865 44.660 96.875 ;
        RECT 31.650 96.495 62.170 96.865 ;
        RECT 31.660 95.700 62.160 96.140 ;
        RECT 31.650 94.970 62.170 95.350 ;
        RECT 30.800 94.715 31.420 94.900 ;
        RECT 62.400 94.715 63.020 94.900 ;
        RECT 30.800 94.485 63.020 94.715 ;
        RECT 30.800 94.300 31.420 94.485 ;
        RECT 62.400 94.300 63.020 94.485 ;
        RECT 39.200 94.220 40.820 94.230 ;
        RECT 31.650 93.850 62.170 94.220 ;
        RECT 31.650 93.130 62.170 93.510 ;
        RECT 30.800 92.875 31.420 93.060 ;
        RECT 62.400 92.875 63.020 93.060 ;
        RECT 30.800 92.645 63.020 92.875 ;
        RECT 30.800 92.460 31.420 92.645 ;
        RECT 62.400 92.460 63.020 92.645 ;
        RECT 35.360 92.380 36.980 92.390 ;
        RECT 31.650 92.010 62.170 92.380 ;
        RECT 31.650 91.290 62.170 91.670 ;
        RECT 30.800 91.035 31.420 91.220 ;
        RECT 62.400 91.035 63.020 91.220 ;
        RECT 30.800 90.805 63.020 91.035 ;
        RECT 30.800 90.620 31.420 90.805 ;
        RECT 62.400 90.620 63.020 90.805 ;
        RECT 31.650 90.170 62.170 90.540 ;
        RECT 25.090 87.820 27.380 88.160 ;
        RECT 28.125 87.820 29.610 88.160 ;
        RECT 25.090 87.185 25.690 87.820 ;
        RECT 25.090 86.955 26.670 87.185 ;
        RECT 25.090 84.915 25.690 86.955 ;
        RECT 27.100 86.725 27.460 86.810 ;
        RECT 25.970 86.495 27.460 86.725 ;
        RECT 25.970 86.345 26.330 86.495 ;
        RECT 25.920 85.710 26.870 86.115 ;
        RECT 25.090 84.685 26.380 84.915 ;
        RECT 25.090 83.725 25.690 84.685 ;
        RECT 26.610 84.365 26.870 85.710 ;
        RECT 27.100 85.060 27.460 86.495 ;
        RECT 27.690 85.160 28.040 86.360 ;
        RECT 28.400 85.750 28.780 87.395 ;
        RECT 27.480 84.365 27.830 84.425 ;
        RECT 28.400 84.365 28.740 84.970 ;
        RECT 26.610 84.105 28.740 84.365 ;
        RECT 27.480 84.045 27.830 84.105 ;
        RECT 29.010 83.825 29.610 87.820 ;
        RECT 31.455 87.385 33.205 90.170 ;
        RECT 33.845 87.385 34.655 88.385 ;
        RECT 35.295 87.385 37.045 89.680 ;
        RECT 37.685 87.385 38.495 88.385 ;
        RECT 39.135 87.385 40.885 89.680 ;
        RECT 41.525 87.385 42.335 88.385 ;
        RECT 42.975 87.385 44.725 89.680 ;
        RECT 45.365 87.385 46.175 88.385 ;
        RECT 46.815 87.385 48.565 89.680 ;
        RECT 49.205 87.385 50.015 88.385 ;
        RECT 50.655 87.385 52.405 89.680 ;
        RECT 53.045 87.385 53.855 88.385 ;
        RECT 54.495 87.385 56.245 89.680 ;
        RECT 56.885 87.385 57.695 88.385 ;
        RECT 58.335 87.385 60.085 89.680 ;
        RECT 60.725 87.385 61.535 88.385 ;
        RECT 63.950 87.575 64.320 106.085 ;
        RECT 64.970 102.450 65.340 106.085 ;
        RECT 64.965 102.070 65.345 102.450 ;
        RECT 64.970 99.450 65.340 102.070 ;
        RECT 64.965 99.070 65.345 99.450 ;
        RECT 64.970 96.450 65.340 99.070 ;
        RECT 64.965 96.070 65.345 96.450 ;
        RECT 64.970 93.450 65.340 96.070 ;
        RECT 64.965 93.070 65.345 93.450 ;
        RECT 64.970 90.450 65.340 93.070 ;
        RECT 64.965 90.070 65.345 90.450 ;
        RECT 63.950 87.195 64.330 87.575 ;
        RECT 63.950 86.125 64.320 87.195 ;
        RECT 31.925 84.935 32.735 85.935 ;
        RECT 25.090 83.495 26.780 83.725 ;
        RECT 28.150 83.595 29.610 83.825 ;
        RECT 25.090 81.485 25.690 83.495 ;
        RECT 27.110 83.035 28.110 83.360 ;
        RECT 25.920 82.475 28.780 82.805 ;
        RECT 25.090 81.255 26.780 81.485 ;
        RECT 25.090 79.245 25.690 81.255 ;
        RECT 27.495 81.120 27.760 82.475 ;
        RECT 29.010 81.585 29.610 83.595 ;
        RECT 33.375 83.105 35.125 85.935 ;
        RECT 35.765 84.935 36.575 85.935 ;
        RECT 37.215 83.640 38.965 85.935 ;
        RECT 39.605 84.935 40.415 85.935 ;
        RECT 41.055 83.640 42.805 85.935 ;
        RECT 43.445 84.935 44.255 85.935 ;
        RECT 44.895 83.640 46.645 85.935 ;
        RECT 47.285 84.935 48.095 85.935 ;
        RECT 48.735 83.640 50.485 85.935 ;
        RECT 51.125 84.935 51.935 85.935 ;
        RECT 52.575 83.640 54.325 85.935 ;
        RECT 54.965 84.935 55.775 85.935 ;
        RECT 56.415 83.640 58.165 85.935 ;
        RECT 58.805 84.935 59.615 85.935 ;
        RECT 60.255 83.640 62.005 85.935 ;
        RECT 63.950 85.745 64.330 86.125 ;
        RECT 31.650 82.735 62.170 83.105 ;
        RECT 30.800 82.470 31.420 82.655 ;
        RECT 62.400 82.470 63.020 82.655 ;
        RECT 30.800 82.240 63.020 82.470 ;
        RECT 30.800 82.055 31.420 82.240 ;
        RECT 62.400 82.055 63.020 82.240 ;
        RECT 31.650 81.605 62.170 81.985 ;
        RECT 28.150 81.355 29.610 81.585 ;
        RECT 27.110 80.795 28.110 81.120 ;
        RECT 25.920 80.235 28.780 80.565 ;
        RECT 29.010 79.345 29.610 81.355 ;
        RECT 31.650 80.895 62.170 81.265 ;
        RECT 37.280 80.885 38.900 80.895 ;
        RECT 30.800 80.630 31.420 80.815 ;
        RECT 62.400 80.630 63.020 80.815 ;
        RECT 30.800 80.400 63.020 80.630 ;
        RECT 30.800 80.215 31.420 80.400 ;
        RECT 62.400 80.215 63.020 80.400 ;
        RECT 31.650 79.765 62.170 80.145 ;
        RECT 25.090 79.015 26.780 79.245 ;
        RECT 28.150 79.115 29.610 79.345 ;
        RECT 25.090 76.960 25.690 79.015 ;
        RECT 27.110 78.555 28.110 78.880 ;
        RECT 29.010 76.960 29.610 79.115 ;
        RECT 31.650 79.050 62.170 79.420 ;
        RECT 41.120 79.040 42.740 79.050 ;
        RECT 30.800 78.785 31.420 78.970 ;
        RECT 62.400 78.785 63.020 78.970 ;
        RECT 30.800 78.555 63.020 78.785 ;
        RECT 30.800 78.370 31.420 78.555 ;
        RECT 62.400 78.370 63.020 78.555 ;
        RECT 31.650 77.920 62.170 78.300 ;
        RECT 31.660 77.130 62.160 77.570 ;
        RECT 25.090 76.620 27.380 76.960 ;
        RECT 28.125 76.620 29.610 76.960 ;
        RECT 25.090 66.885 25.690 76.620 ;
        RECT 29.010 66.885 29.610 76.620 ;
        RECT 31.650 76.410 62.170 76.780 ;
        RECT 44.960 76.400 46.580 76.410 ;
        RECT 30.800 76.145 31.420 76.330 ;
        RECT 62.400 76.145 63.020 76.330 ;
        RECT 30.800 75.915 63.020 76.145 ;
        RECT 30.800 75.730 31.420 75.915 ;
        RECT 62.400 75.730 63.020 75.915 ;
        RECT 31.650 75.280 62.170 75.660 ;
        RECT 31.650 74.570 62.170 74.940 ;
        RECT 48.800 74.560 50.420 74.570 ;
        RECT 30.800 74.305 31.420 74.490 ;
        RECT 62.400 74.305 63.020 74.490 ;
        RECT 30.800 74.075 63.020 74.305 ;
        RECT 30.800 73.890 31.420 74.075 ;
        RECT 62.400 73.890 63.020 74.075 ;
        RECT 31.650 73.440 62.170 73.820 ;
        RECT 31.650 72.725 62.170 73.095 ;
        RECT 52.640 72.715 54.260 72.725 ;
        RECT 30.800 72.460 31.420 72.645 ;
        RECT 62.400 72.460 63.020 72.645 ;
        RECT 30.800 72.230 63.020 72.460 ;
        RECT 30.800 72.045 31.420 72.230 ;
        RECT 62.400 72.045 63.020 72.230 ;
        RECT 31.650 71.595 62.170 71.975 ;
        RECT 31.660 70.805 62.160 71.245 ;
        RECT 31.650 70.085 62.170 70.455 ;
        RECT 56.480 70.075 58.100 70.085 ;
        RECT 30.800 69.820 31.420 70.005 ;
        RECT 62.400 69.820 63.020 70.005 ;
        RECT 30.800 69.590 63.020 69.820 ;
        RECT 30.800 69.405 31.420 69.590 ;
        RECT 62.400 69.405 63.020 69.590 ;
        RECT 31.650 68.955 62.170 69.335 ;
        RECT 31.650 68.245 62.170 68.615 ;
        RECT 60.320 68.235 61.940 68.245 ;
        RECT 30.800 67.980 31.420 68.165 ;
        RECT 62.400 67.980 63.020 68.165 ;
        RECT 30.800 67.750 63.020 67.980 ;
        RECT 63.950 67.815 64.320 85.745 ;
        RECT 64.970 84.450 65.340 90.070 ;
        RECT 65.990 87.575 66.360 106.085 ;
        RECT 67.010 102.450 67.380 106.085 ;
        RECT 67.005 102.070 67.385 102.450 ;
        RECT 67.010 99.450 67.380 102.070 ;
        RECT 67.005 99.070 67.385 99.450 ;
        RECT 67.010 96.450 67.380 99.070 ;
        RECT 67.005 96.070 67.385 96.450 ;
        RECT 67.010 93.450 67.380 96.070 ;
        RECT 67.005 93.070 67.385 93.450 ;
        RECT 67.010 90.450 67.380 93.070 ;
        RECT 67.005 90.070 67.385 90.450 ;
        RECT 65.990 87.195 66.370 87.575 ;
        RECT 65.990 86.125 66.360 87.195 ;
        RECT 65.990 85.745 66.370 86.125 ;
        RECT 64.965 84.070 65.345 84.450 ;
        RECT 64.970 81.450 65.340 84.070 ;
        RECT 64.965 81.070 65.345 81.450 ;
        RECT 64.970 78.450 65.340 81.070 ;
        RECT 64.965 78.070 65.345 78.450 ;
        RECT 64.970 75.450 65.340 78.070 ;
        RECT 64.965 75.070 65.345 75.450 ;
        RECT 64.970 72.450 65.340 75.070 ;
        RECT 64.965 72.070 65.345 72.450 ;
        RECT 64.970 69.450 65.340 72.070 ;
        RECT 64.965 69.070 65.345 69.450 ;
        RECT 64.970 67.815 65.340 69.070 ;
        RECT 65.990 67.815 66.360 85.745 ;
        RECT 67.010 84.450 67.380 90.070 ;
        RECT 67.005 84.070 67.385 84.450 ;
        RECT 67.010 81.450 67.380 84.070 ;
        RECT 67.005 81.070 67.385 81.450 ;
        RECT 67.010 78.450 67.380 81.070 ;
        RECT 67.005 78.070 67.385 78.450 ;
        RECT 67.010 75.450 67.380 78.070 ;
        RECT 67.005 75.070 67.385 75.450 ;
        RECT 67.010 72.450 67.380 75.070 ;
        RECT 67.005 72.070 67.385 72.450 ;
        RECT 67.010 69.450 67.380 72.070 ;
        RECT 67.005 69.070 67.385 69.450 ;
        RECT 67.010 67.815 67.380 69.070 ;
        RECT 68.030 67.815 68.410 106.085 ;
        RECT 68.760 67.825 69.200 106.075 ;
        RECT 30.800 67.565 31.420 67.750 ;
        RECT 62.400 67.565 63.020 67.750 ;
        RECT 31.650 67.115 62.170 67.495 ;
      LAYER Metal2 ;
        RECT 31.920 105.780 34.160 106.160 ;
        RECT 62.520 105.220 62.900 105.600 ;
        RECT 25.200 103.570 25.580 103.950 ;
        RECT 29.120 103.570 29.500 103.950 ;
        RECT 31.920 103.940 34.160 104.320 ;
        RECT 31.925 102.055 34.165 102.435 ;
        RECT 31.920 101.295 34.160 101.675 ;
        RECT 25.200 100.570 25.580 100.950 ;
        RECT 29.120 100.570 29.500 100.950 ;
        RECT 31.920 99.455 34.160 99.835 ;
        RECT 25.200 97.570 25.580 97.950 ;
        RECT 29.120 97.570 29.500 97.950 ;
        RECT 31.920 97.615 34.160 97.995 ;
        RECT 31.925 95.730 34.165 96.110 ;
        RECT 31.920 94.970 34.160 95.350 ;
        RECT 25.200 94.570 25.580 94.950 ;
        RECT 29.120 94.570 29.500 94.950 ;
        RECT 31.920 93.130 34.160 93.510 ;
        RECT 25.200 91.570 25.580 91.950 ;
        RECT 29.120 91.570 29.500 91.950 ;
        RECT 31.920 91.290 34.160 91.670 ;
        RECT 25.200 88.570 25.580 88.950 ;
        RECT 29.120 88.570 29.500 88.950 ;
        RECT 35.295 88.580 37.045 92.390 ;
        RECT 39.135 88.580 40.885 94.230 ;
        RECT 42.975 88.580 44.725 96.875 ;
        RECT 46.815 88.580 48.565 98.715 ;
        RECT 50.655 88.580 52.405 100.555 ;
        RECT 54.495 88.580 56.245 103.200 ;
        RECT 58.335 88.580 60.085 105.040 ;
        RECT 62.520 103.380 62.900 103.760 ;
        RECT 64.965 102.070 65.345 102.450 ;
        RECT 67.005 102.070 67.385 102.450 ;
        RECT 68.790 102.070 69.170 102.450 ;
        RECT 62.520 100.735 62.900 101.115 ;
        RECT 62.520 98.895 62.900 99.275 ;
        RECT 64.965 99.070 65.345 99.450 ;
        RECT 67.005 99.070 67.385 99.450 ;
        RECT 68.790 99.070 69.170 99.450 ;
        RECT 62.520 97.055 62.900 97.435 ;
        RECT 64.965 96.070 65.345 96.450 ;
        RECT 67.005 96.070 67.385 96.450 ;
        RECT 68.790 96.070 69.170 96.450 ;
        RECT 62.520 94.410 62.900 94.790 ;
        RECT 64.965 93.070 65.345 93.450 ;
        RECT 67.005 93.070 67.385 93.450 ;
        RECT 68.790 93.070 69.170 93.450 ;
        RECT 62.520 92.570 62.900 92.950 ;
        RECT 62.520 90.730 62.900 91.110 ;
        RECT 64.965 90.070 65.345 90.450 ;
        RECT 67.005 90.070 67.385 90.450 ;
        RECT 68.790 90.070 69.170 90.450 ;
        RECT 34.060 88.195 34.440 88.385 ;
        RECT 37.900 88.195 38.280 88.385 ;
        RECT 41.740 88.195 42.120 88.385 ;
        RECT 45.580 88.195 45.960 88.385 ;
        RECT 49.420 88.195 49.800 88.385 ;
        RECT 53.260 88.195 53.640 88.385 ;
        RECT 57.100 88.195 57.480 88.385 ;
        RECT 60.940 88.195 61.320 88.385 ;
        RECT 28.390 87.385 69.440 88.195 ;
        RECT 25.200 85.570 25.580 85.950 ;
        RECT 28.390 85.935 29.200 87.385 ;
        RECT 63.950 87.195 64.330 87.385 ;
        RECT 65.990 87.195 66.370 87.385 ;
        RECT 68.030 87.195 68.410 87.385 ;
        RECT 63.950 85.935 64.330 86.125 ;
        RECT 65.990 85.935 66.370 86.125 ;
        RECT 68.030 85.935 68.410 86.125 ;
        RECT 28.390 85.125 69.440 85.935 ;
        RECT 32.140 84.935 32.520 85.125 ;
        RECT 35.980 84.935 36.360 85.125 ;
        RECT 39.820 84.935 40.200 85.125 ;
        RECT 43.660 84.935 44.040 85.125 ;
        RECT 47.500 84.935 47.880 85.125 ;
        RECT 51.340 84.935 51.720 85.125 ;
        RECT 55.180 84.935 55.560 85.125 ;
        RECT 59.020 84.935 59.400 85.125 ;
        RECT 25.200 82.570 25.580 82.950 ;
        RECT 27.480 80.235 27.830 84.425 ;
        RECT 25.200 79.570 25.580 79.950 ;
        RECT 28.110 78.880 28.460 82.795 ;
        RECT 29.120 82.570 29.500 82.950 ;
        RECT 31.920 81.605 34.160 81.985 ;
        RECT 37.215 80.885 38.965 84.740 ;
        RECT 29.120 79.570 29.500 79.950 ;
        RECT 31.920 79.765 34.160 80.145 ;
        RECT 41.055 79.040 42.805 84.740 ;
        RECT 27.705 78.555 28.460 78.880 ;
        RECT 28.110 78.550 28.460 78.555 ;
        RECT 31.920 77.920 34.160 78.300 ;
        RECT 31.925 77.160 34.165 77.540 ;
        RECT 25.200 76.570 25.580 76.950 ;
        RECT 29.120 76.570 29.500 76.950 ;
        RECT 44.895 76.400 46.645 84.740 ;
        RECT 31.920 75.280 34.160 75.660 ;
        RECT 48.735 74.560 50.485 84.740 ;
        RECT 25.200 73.570 25.580 73.950 ;
        RECT 29.120 73.570 29.500 73.950 ;
        RECT 31.920 73.440 34.160 73.820 ;
        RECT 52.575 72.715 54.325 84.740 ;
        RECT 31.920 71.595 34.160 71.975 ;
        RECT 25.200 70.570 25.580 70.950 ;
        RECT 29.120 70.570 29.500 70.950 ;
        RECT 31.925 70.835 34.165 71.215 ;
        RECT 56.415 70.075 58.165 84.740 ;
        RECT 31.920 68.955 34.160 69.335 ;
        RECT 60.255 68.235 62.005 84.740 ;
        RECT 64.965 84.070 65.345 84.450 ;
        RECT 67.005 84.070 67.385 84.450 ;
        RECT 68.790 84.070 69.170 84.450 ;
        RECT 62.520 82.165 62.900 82.545 ;
        RECT 64.965 81.070 65.345 81.450 ;
        RECT 67.005 81.070 67.385 81.450 ;
        RECT 68.790 81.070 69.170 81.450 ;
        RECT 62.520 80.325 62.900 80.705 ;
        RECT 62.520 78.480 62.900 78.860 ;
        RECT 64.965 78.070 65.345 78.450 ;
        RECT 67.005 78.070 67.385 78.450 ;
        RECT 68.790 78.070 69.170 78.450 ;
        RECT 62.520 75.840 62.900 76.220 ;
        RECT 64.965 75.070 65.345 75.450 ;
        RECT 67.005 75.070 67.385 75.450 ;
        RECT 68.790 75.070 69.170 75.450 ;
        RECT 62.520 74.000 62.900 74.380 ;
        RECT 62.520 72.155 62.900 72.535 ;
        RECT 64.965 72.070 65.345 72.450 ;
        RECT 67.005 72.070 67.385 72.450 ;
        RECT 68.790 72.070 69.170 72.450 ;
        RECT 62.520 69.515 62.900 69.895 ;
        RECT 64.965 69.070 65.345 69.450 ;
        RECT 67.005 69.070 67.385 69.450 ;
        RECT 68.790 69.070 69.170 69.450 ;
        RECT 25.200 67.570 25.580 67.950 ;
        RECT 29.120 67.570 29.500 67.950 ;
        RECT 62.520 67.675 62.900 68.055 ;
        RECT 31.920 67.115 34.160 67.495 ;
      LAYER Metal3 ;
        RECT 31.920 105.780 34.160 106.160 ;
        RECT 53.700 105.550 54.080 105.600 ;
        RECT 62.520 105.550 62.900 105.600 ;
        RECT 53.700 105.270 62.900 105.550 ;
        RECT 53.700 105.220 54.080 105.270 ;
        RECT 62.520 105.220 62.900 105.270 ;
        RECT 25.200 103.570 25.580 103.950 ;
        RECT 29.120 103.570 29.500 103.950 ;
        RECT 31.920 103.940 34.160 104.320 ;
        RECT 54.980 103.710 55.360 103.760 ;
        RECT 62.520 103.710 62.900 103.760 ;
        RECT 54.980 103.430 62.900 103.710 ;
        RECT 54.980 103.380 55.360 103.430 ;
        RECT 62.520 103.380 62.900 103.430 ;
        RECT 31.925 102.055 34.165 102.435 ;
        RECT 64.965 102.070 65.345 102.450 ;
        RECT 67.005 102.070 67.385 102.450 ;
        RECT 68.790 102.070 69.170 102.450 ;
        RECT 31.920 101.295 34.160 101.675 ;
        RECT 56.260 101.065 56.640 101.115 ;
        RECT 62.520 101.065 62.900 101.115 ;
        RECT 25.200 100.570 25.580 100.950 ;
        RECT 29.120 100.570 29.500 100.950 ;
        RECT 56.260 100.785 62.900 101.065 ;
        RECT 56.260 100.735 56.640 100.785 ;
        RECT 62.520 100.735 62.900 100.785 ;
        RECT 31.920 99.455 34.160 99.835 ;
        RECT 57.540 99.225 57.920 99.275 ;
        RECT 62.520 99.225 62.900 99.275 ;
        RECT 57.540 98.945 62.900 99.225 ;
        RECT 64.965 99.070 65.345 99.450 ;
        RECT 67.005 99.070 67.385 99.450 ;
        RECT 68.790 99.070 69.170 99.450 ;
        RECT 57.540 98.895 57.920 98.945 ;
        RECT 62.520 98.895 62.900 98.945 ;
        RECT 25.200 97.570 25.580 97.950 ;
        RECT 29.120 97.570 29.500 97.950 ;
        RECT 31.920 97.615 34.160 97.995 ;
        RECT 58.820 97.385 59.200 97.435 ;
        RECT 62.520 97.385 62.900 97.435 ;
        RECT 58.820 97.105 62.900 97.385 ;
        RECT 58.820 97.055 59.200 97.105 ;
        RECT 62.520 97.055 62.900 97.105 ;
        RECT 31.925 95.730 34.165 96.110 ;
        RECT 64.965 96.070 65.345 96.450 ;
        RECT 67.005 96.070 67.385 96.450 ;
        RECT 68.790 96.070 69.170 96.450 ;
        RECT 31.920 94.970 34.160 95.350 ;
        RECT 25.200 94.570 25.580 94.950 ;
        RECT 29.120 94.570 29.500 94.950 ;
        RECT 60.100 94.740 60.480 94.790 ;
        RECT 62.520 94.740 62.900 94.790 ;
        RECT 60.100 94.460 62.900 94.740 ;
        RECT 60.100 94.410 60.480 94.460 ;
        RECT 62.520 94.410 62.900 94.460 ;
        RECT 31.920 93.130 34.160 93.510 ;
        RECT 64.965 93.070 65.345 93.450 ;
        RECT 67.005 93.070 67.385 93.450 ;
        RECT 68.790 93.070 69.170 93.450 ;
        RECT 61.380 92.900 61.760 92.950 ;
        RECT 62.520 92.900 62.900 92.950 ;
        RECT 61.380 92.620 62.900 92.900 ;
        RECT 61.380 92.570 61.760 92.620 ;
        RECT 62.520 92.570 62.900 92.620 ;
        RECT 25.200 91.570 25.580 91.950 ;
        RECT 29.120 91.570 29.500 91.950 ;
        RECT 31.920 91.290 34.160 91.670 ;
        RECT 62.520 90.730 63.040 91.110 ;
        RECT 64.965 90.070 65.345 90.450 ;
        RECT 67.005 90.070 67.385 90.450 ;
        RECT 68.790 90.070 69.170 90.450 ;
        RECT 25.200 88.570 25.580 88.950 ;
        RECT 29.120 88.570 29.500 88.950 ;
        RECT 25.200 85.570 25.580 85.950 ;
        RECT 64.965 84.070 65.345 84.450 ;
        RECT 67.005 84.070 67.385 84.450 ;
        RECT 68.790 84.070 69.170 84.450 ;
        RECT 25.200 82.570 25.580 82.950 ;
        RECT 29.120 82.570 29.500 82.950 ;
        RECT 62.020 82.165 62.900 82.545 ;
        RECT 31.920 81.605 34.160 81.985 ;
        RECT 64.965 81.070 65.345 81.450 ;
        RECT 67.005 81.070 67.385 81.450 ;
        RECT 68.790 81.070 69.170 81.450 ;
        RECT 60.740 80.655 61.120 80.705 ;
        RECT 62.520 80.655 62.900 80.705 ;
        RECT 60.740 80.375 62.900 80.655 ;
        RECT 60.740 80.325 61.120 80.375 ;
        RECT 62.520 80.325 62.900 80.375 ;
        RECT 25.200 79.570 25.580 79.950 ;
        RECT 29.120 79.570 29.500 79.950 ;
        RECT 31.920 79.765 34.160 80.145 ;
        RECT 59.460 78.810 59.840 78.860 ;
        RECT 62.520 78.810 62.900 78.860 ;
        RECT 59.460 78.530 62.900 78.810 ;
        RECT 59.460 78.480 59.840 78.530 ;
        RECT 62.520 78.480 62.900 78.530 ;
        RECT 31.920 77.920 34.160 78.300 ;
        RECT 64.965 78.070 65.345 78.450 ;
        RECT 67.005 78.070 67.385 78.450 ;
        RECT 68.790 78.070 69.170 78.450 ;
        RECT 31.925 77.160 34.165 77.540 ;
        RECT 25.200 76.570 25.580 76.950 ;
        RECT 29.120 76.570 29.500 76.950 ;
        RECT 58.180 76.170 58.560 76.220 ;
        RECT 62.520 76.170 62.900 76.220 ;
        RECT 58.180 75.890 62.900 76.170 ;
        RECT 58.180 75.840 58.560 75.890 ;
        RECT 62.520 75.840 62.900 75.890 ;
        RECT 31.920 75.280 34.160 75.660 ;
        RECT 64.965 75.070 65.345 75.450 ;
        RECT 67.005 75.070 67.385 75.450 ;
        RECT 68.790 75.070 69.170 75.450 ;
        RECT 56.900 74.330 57.280 74.380 ;
        RECT 62.520 74.330 62.900 74.380 ;
        RECT 56.900 74.050 62.900 74.330 ;
        RECT 56.900 74.000 57.280 74.050 ;
        RECT 62.520 74.000 62.900 74.050 ;
        RECT 25.200 73.570 25.580 73.950 ;
        RECT 29.120 73.570 29.500 73.950 ;
        RECT 31.920 73.440 34.160 73.820 ;
        RECT 55.620 72.485 56.000 72.535 ;
        RECT 62.520 72.485 62.900 72.535 ;
        RECT 55.620 72.205 62.900 72.485 ;
        RECT 55.620 72.155 56.000 72.205 ;
        RECT 62.520 72.155 62.900 72.205 ;
        RECT 64.965 72.070 65.345 72.450 ;
        RECT 67.005 72.070 67.385 72.450 ;
        RECT 68.790 72.070 69.170 72.450 ;
        RECT 31.920 71.595 34.160 71.975 ;
        RECT 25.200 70.570 25.580 70.950 ;
        RECT 29.120 70.570 29.500 70.950 ;
        RECT 31.925 70.835 34.165 71.215 ;
        RECT 54.340 69.845 54.720 69.895 ;
        RECT 62.520 69.845 62.900 69.895 ;
        RECT 54.340 69.565 62.900 69.845 ;
        RECT 54.340 69.515 54.720 69.565 ;
        RECT 62.520 69.515 62.900 69.565 ;
        RECT 31.920 68.955 34.160 69.335 ;
        RECT 64.965 69.070 65.345 69.450 ;
        RECT 67.005 69.070 67.385 69.450 ;
        RECT 68.790 69.070 69.170 69.450 ;
        RECT 53.060 68.005 53.440 68.055 ;
        RECT 62.520 68.005 62.900 68.055 ;
        RECT 25.200 67.570 25.580 67.950 ;
        RECT 29.120 67.570 29.500 67.950 ;
        RECT 53.060 67.725 62.900 68.005 ;
        RECT 53.060 67.675 53.440 67.725 ;
        RECT 62.520 67.675 62.900 67.725 ;
        RECT 31.920 67.115 34.160 67.495 ;
  END
END efuse_array_16x1
END LIBRARY

