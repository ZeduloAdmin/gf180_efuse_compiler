VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO efuse_array_64x8
  CLASS BLOCK ;
  FOREIGN efuse_array_64x8 ;
  ORIGIN -24.960 -66.885 ;
  SIZE 141.830 BY 315.825 ;
  PIN COL_PROG_N[0]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 161.750 106.315 165.310 106.615 ;
    END
  END COL_PROG_N[0]
  PIN OUT[0]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 77.995 28.780 78.325 ;
    END
  END OUT[0]
  PIN COL_PROG_N[1]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 161.750 145.700 165.310 146.000 ;
    END
  END COL_PROG_N[1]
  PIN OUT[1]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 117.380 28.780 117.710 ;
    END
  END OUT[1]
  PIN COL_PROG_N[2]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 161.750 185.085 165.310 185.385 ;
    END
  END COL_PROG_N[2]
  PIN OUT[2]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 156.765 28.780 157.095 ;
    END
  END OUT[2]
  PIN COL_PROG_N[3]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 161.750 224.470 165.310 224.770 ;
    END
  END COL_PROG_N[3]
  PIN OUT[3]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 196.150 28.780 196.480 ;
    END
  END OUT[3]
  PIN COL_PROG_N[4]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 161.750 263.855 165.310 264.155 ;
    END
  END COL_PROG_N[4]
  PIN OUT[4]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 235.535 28.780 235.865 ;
    END
  END OUT[4]
  PIN COL_PROG_N[5]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 161.750 303.240 165.310 303.540 ;
    END
  END COL_PROG_N[5]
  PIN OUT[5]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 274.920 28.780 275.250 ;
    END
  END OUT[5]
  PIN COL_PROG_N[6]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 161.750 342.625 165.310 342.925 ;
    END
  END COL_PROG_N[6]
  PIN OUT[6]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 314.305 28.780 314.635 ;
    END
  END OUT[6]
  PIN COL_PROG_N[7]
    ANTENNAGATEAREA 76.500000 ;
    PORT
      LAYER Metal1 ;
        RECT 161.750 382.010 165.310 382.310 ;
    END
  END COL_PROG_N[7]
  PIN OUT[7]
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 25.920 353.690 28.780 354.020 ;
    END
  END OUT[7]
  PIN PRESET_N
    ANTENNAGATEAREA 9.760000 ;
    PORT
      LAYER Metal2 ;
        RECT 25.970 362.420 26.250 382.710 ;
        RECT 25.970 362.040 26.330 362.420 ;
        RECT 25.970 323.035 26.250 362.040 ;
        RECT 25.970 322.655 26.330 323.035 ;
        RECT 25.970 283.650 26.250 322.655 ;
        RECT 25.970 283.270 26.330 283.650 ;
        RECT 25.970 244.265 26.250 283.270 ;
        RECT 25.970 243.885 26.330 244.265 ;
        RECT 25.970 204.880 26.250 243.885 ;
        RECT 25.970 204.500 26.330 204.880 ;
        RECT 25.970 165.495 26.250 204.500 ;
        RECT 25.970 165.115 26.330 165.495 ;
        RECT 25.970 126.110 26.250 165.115 ;
        RECT 25.970 125.730 26.330 126.110 ;
        RECT 25.970 86.725 26.250 125.730 ;
        RECT 25.970 86.345 26.330 86.725 ;
        RECT 25.970 66.885 26.250 86.345 ;
    END
  END PRESET_N
  PIN SENSE
    ANTENNAGATEAREA 3.936000 ;
    PORT
      LAYER Metal2 ;
        RECT 26.615 361.235 26.895 382.710 ;
        RECT 26.615 360.855 28.040 361.235 ;
        RECT 26.615 321.850 26.895 360.855 ;
        RECT 26.615 321.470 28.040 321.850 ;
        RECT 26.615 282.465 26.895 321.470 ;
        RECT 26.615 282.085 28.040 282.465 ;
        RECT 26.615 243.080 26.895 282.085 ;
        RECT 26.615 242.700 28.040 243.080 ;
        RECT 26.615 203.695 26.895 242.700 ;
        RECT 26.615 203.315 28.040 203.695 ;
        RECT 26.615 164.310 26.895 203.315 ;
        RECT 26.615 163.930 28.040 164.310 ;
        RECT 26.615 124.925 26.895 163.930 ;
        RECT 26.615 124.545 28.040 124.925 ;
        RECT 26.615 85.540 26.895 124.545 ;
        RECT 26.615 85.160 28.040 85.540 ;
        RECT 26.615 66.885 26.895 85.160 ;
    END
  END SENSE
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 128.780 66.885 131.780 382.710 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 96.330 66.885 99.330 382.710 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 63.880 66.885 66.880 382.710 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 28.670 66.885 29.670 382.710 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 31.430 66.885 34.430 382.710 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 162.300 66.885 166.550 382.710 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 25.030 66.885 26.030 382.710 ;
    END
  END VDD
  PIN BIT_SEL[48]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 160.050 366.805 160.330 382.085 ;
        RECT 160.010 366.425 160.390 366.805 ;
        RECT 160.050 327.420 160.330 366.425 ;
        RECT 160.010 327.040 160.390 327.420 ;
        RECT 160.050 288.035 160.330 327.040 ;
        RECT 160.010 287.655 160.390 288.035 ;
        RECT 160.050 248.650 160.330 287.655 ;
        RECT 160.010 248.270 160.390 248.650 ;
        RECT 160.050 209.265 160.330 248.270 ;
        RECT 160.010 208.885 160.390 209.265 ;
        RECT 160.050 169.880 160.330 208.885 ;
        RECT 160.010 169.500 160.390 169.880 ;
        RECT 160.050 130.495 160.330 169.500 ;
        RECT 160.010 130.115 160.390 130.495 ;
        RECT 160.050 91.110 160.330 130.115 ;
        RECT 160.010 90.730 160.390 91.110 ;
        RECT 160.050 66.885 160.330 90.730 ;
    END
  END BIT_SEL[48]
  PIN BIT_SEL[49]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 159.410 358.240 159.690 382.085 ;
        RECT 159.370 357.860 159.750 358.240 ;
        RECT 159.410 318.855 159.690 357.860 ;
        RECT 159.370 318.475 159.750 318.855 ;
        RECT 159.410 279.470 159.690 318.475 ;
        RECT 159.370 279.090 159.750 279.470 ;
        RECT 159.410 240.085 159.690 279.090 ;
        RECT 159.370 239.705 159.750 240.085 ;
        RECT 159.410 200.700 159.690 239.705 ;
        RECT 159.370 200.320 159.750 200.700 ;
        RECT 159.410 161.315 159.690 200.320 ;
        RECT 159.370 160.935 159.750 161.315 ;
        RECT 159.410 121.930 159.690 160.935 ;
        RECT 159.370 121.550 159.750 121.930 ;
        RECT 159.410 82.545 159.690 121.550 ;
        RECT 159.370 82.165 159.750 82.545 ;
        RECT 159.410 66.885 159.690 82.165 ;
    END
  END BIT_SEL[49]
  PIN BIT_SEL[50]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 158.770 368.645 159.050 382.085 ;
        RECT 158.730 368.265 159.110 368.645 ;
        RECT 158.770 329.260 159.050 368.265 ;
        RECT 158.730 328.880 159.110 329.260 ;
        RECT 158.770 289.875 159.050 328.880 ;
        RECT 158.730 289.495 159.110 289.875 ;
        RECT 158.770 250.490 159.050 289.495 ;
        RECT 158.730 250.110 159.110 250.490 ;
        RECT 158.770 211.105 159.050 250.110 ;
        RECT 158.730 210.725 159.110 211.105 ;
        RECT 158.770 171.720 159.050 210.725 ;
        RECT 158.730 171.340 159.110 171.720 ;
        RECT 158.770 132.335 159.050 171.340 ;
        RECT 158.730 131.955 159.110 132.335 ;
        RECT 158.770 92.950 159.050 131.955 ;
        RECT 158.730 92.570 159.110 92.950 ;
        RECT 158.770 66.885 159.050 92.570 ;
    END
  END BIT_SEL[50]
  PIN BIT_SEL[51]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 158.130 356.400 158.410 382.085 ;
        RECT 158.090 356.020 158.470 356.400 ;
        RECT 158.130 317.015 158.410 356.020 ;
        RECT 158.090 316.635 158.470 317.015 ;
        RECT 158.130 277.630 158.410 316.635 ;
        RECT 158.090 277.250 158.470 277.630 ;
        RECT 158.130 238.245 158.410 277.250 ;
        RECT 158.090 237.865 158.470 238.245 ;
        RECT 158.130 198.860 158.410 237.865 ;
        RECT 158.090 198.480 158.470 198.860 ;
        RECT 158.130 159.475 158.410 198.480 ;
        RECT 158.090 159.095 158.470 159.475 ;
        RECT 158.130 120.090 158.410 159.095 ;
        RECT 158.090 119.710 158.470 120.090 ;
        RECT 158.130 80.705 158.410 119.710 ;
        RECT 158.090 80.325 158.470 80.705 ;
        RECT 158.130 66.885 158.410 80.325 ;
    END
  END BIT_SEL[51]
  PIN BIT_SEL[52]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 157.490 370.485 157.770 382.085 ;
        RECT 157.450 370.105 157.830 370.485 ;
        RECT 157.490 331.100 157.770 370.105 ;
        RECT 157.450 330.720 157.830 331.100 ;
        RECT 157.490 291.715 157.770 330.720 ;
        RECT 157.450 291.335 157.830 291.715 ;
        RECT 157.490 252.330 157.770 291.335 ;
        RECT 157.450 251.950 157.830 252.330 ;
        RECT 157.490 212.945 157.770 251.950 ;
        RECT 157.450 212.565 157.830 212.945 ;
        RECT 157.490 173.560 157.770 212.565 ;
        RECT 157.450 173.180 157.830 173.560 ;
        RECT 157.490 134.175 157.770 173.180 ;
        RECT 157.450 133.795 157.830 134.175 ;
        RECT 157.490 94.790 157.770 133.795 ;
        RECT 157.450 94.410 157.830 94.790 ;
        RECT 157.490 66.885 157.770 94.410 ;
    END
  END BIT_SEL[52]
  PIN BIT_SEL[53]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 156.850 354.555 157.130 382.085 ;
        RECT 156.810 354.175 157.190 354.555 ;
        RECT 156.850 315.170 157.130 354.175 ;
        RECT 156.810 314.790 157.190 315.170 ;
        RECT 156.850 275.785 157.130 314.790 ;
        RECT 156.810 275.405 157.190 275.785 ;
        RECT 156.850 236.400 157.130 275.405 ;
        RECT 156.810 236.020 157.190 236.400 ;
        RECT 156.850 197.015 157.130 236.020 ;
        RECT 156.810 196.635 157.190 197.015 ;
        RECT 156.850 157.630 157.130 196.635 ;
        RECT 156.810 157.250 157.190 157.630 ;
        RECT 156.850 118.245 157.130 157.250 ;
        RECT 156.810 117.865 157.190 118.245 ;
        RECT 156.850 78.860 157.130 117.865 ;
        RECT 156.810 78.480 157.190 78.860 ;
        RECT 156.850 66.885 157.130 78.480 ;
    END
  END BIT_SEL[53]
  PIN BIT_SEL[54]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 156.210 373.130 156.490 382.085 ;
        RECT 156.170 372.750 156.550 373.130 ;
        RECT 156.210 333.745 156.490 372.750 ;
        RECT 156.170 333.365 156.550 333.745 ;
        RECT 156.210 294.360 156.490 333.365 ;
        RECT 156.170 293.980 156.550 294.360 ;
        RECT 156.210 254.975 156.490 293.980 ;
        RECT 156.170 254.595 156.550 254.975 ;
        RECT 156.210 215.590 156.490 254.595 ;
        RECT 156.170 215.210 156.550 215.590 ;
        RECT 156.210 176.205 156.490 215.210 ;
        RECT 156.170 175.825 156.550 176.205 ;
        RECT 156.210 136.820 156.490 175.825 ;
        RECT 156.170 136.440 156.550 136.820 ;
        RECT 156.210 97.435 156.490 136.440 ;
        RECT 156.170 97.055 156.550 97.435 ;
        RECT 156.210 66.885 156.490 97.055 ;
    END
  END BIT_SEL[54]
  PIN BIT_SEL[55]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 155.570 351.915 155.850 382.085 ;
        RECT 155.530 351.535 155.910 351.915 ;
        RECT 155.570 312.530 155.850 351.535 ;
        RECT 155.530 312.150 155.910 312.530 ;
        RECT 155.570 273.145 155.850 312.150 ;
        RECT 155.530 272.765 155.910 273.145 ;
        RECT 155.570 233.760 155.850 272.765 ;
        RECT 155.530 233.380 155.910 233.760 ;
        RECT 155.570 194.375 155.850 233.380 ;
        RECT 155.530 193.995 155.910 194.375 ;
        RECT 155.570 154.990 155.850 193.995 ;
        RECT 155.530 154.610 155.910 154.990 ;
        RECT 155.570 115.605 155.850 154.610 ;
        RECT 155.530 115.225 155.910 115.605 ;
        RECT 155.570 76.220 155.850 115.225 ;
        RECT 155.530 75.840 155.910 76.220 ;
        RECT 155.570 66.885 155.850 75.840 ;
    END
  END BIT_SEL[55]
  PIN BIT_SEL[56]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 154.930 374.970 155.210 382.085 ;
        RECT 154.890 374.590 155.270 374.970 ;
        RECT 154.930 335.585 155.210 374.590 ;
        RECT 154.890 335.205 155.270 335.585 ;
        RECT 154.930 296.200 155.210 335.205 ;
        RECT 154.890 295.820 155.270 296.200 ;
        RECT 154.930 256.815 155.210 295.820 ;
        RECT 154.890 256.435 155.270 256.815 ;
        RECT 154.930 217.430 155.210 256.435 ;
        RECT 154.890 217.050 155.270 217.430 ;
        RECT 154.930 178.045 155.210 217.050 ;
        RECT 154.890 177.665 155.270 178.045 ;
        RECT 154.930 138.660 155.210 177.665 ;
        RECT 154.890 138.280 155.270 138.660 ;
        RECT 154.930 99.275 155.210 138.280 ;
        RECT 154.890 98.895 155.270 99.275 ;
        RECT 154.930 66.885 155.210 98.895 ;
    END
  END BIT_SEL[56]
  PIN BIT_SEL[57]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 154.290 350.075 154.570 382.085 ;
        RECT 154.250 349.695 154.630 350.075 ;
        RECT 154.290 310.690 154.570 349.695 ;
        RECT 154.250 310.310 154.630 310.690 ;
        RECT 154.290 271.305 154.570 310.310 ;
        RECT 154.250 270.925 154.630 271.305 ;
        RECT 154.290 231.920 154.570 270.925 ;
        RECT 154.250 231.540 154.630 231.920 ;
        RECT 154.290 192.535 154.570 231.540 ;
        RECT 154.250 192.155 154.630 192.535 ;
        RECT 154.290 153.150 154.570 192.155 ;
        RECT 154.250 152.770 154.630 153.150 ;
        RECT 154.290 113.765 154.570 152.770 ;
        RECT 154.250 113.385 154.630 113.765 ;
        RECT 154.290 74.380 154.570 113.385 ;
        RECT 154.250 74.000 154.630 74.380 ;
        RECT 154.290 66.885 154.570 74.000 ;
    END
  END BIT_SEL[57]
  PIN BIT_SEL[58]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 153.650 376.810 153.930 382.085 ;
        RECT 153.610 376.430 153.990 376.810 ;
        RECT 153.650 337.425 153.930 376.430 ;
        RECT 153.610 337.045 153.990 337.425 ;
        RECT 153.650 298.040 153.930 337.045 ;
        RECT 153.610 297.660 153.990 298.040 ;
        RECT 153.650 258.655 153.930 297.660 ;
        RECT 153.610 258.275 153.990 258.655 ;
        RECT 153.650 219.270 153.930 258.275 ;
        RECT 153.610 218.890 153.990 219.270 ;
        RECT 153.650 179.885 153.930 218.890 ;
        RECT 153.610 179.505 153.990 179.885 ;
        RECT 153.650 140.500 153.930 179.505 ;
        RECT 153.610 140.120 153.990 140.500 ;
        RECT 153.650 101.115 153.930 140.120 ;
        RECT 153.610 100.735 153.990 101.115 ;
        RECT 153.650 66.885 153.930 100.735 ;
    END
  END BIT_SEL[58]
  PIN BIT_SEL[59]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 153.010 348.230 153.290 382.085 ;
        RECT 152.970 347.850 153.350 348.230 ;
        RECT 153.010 308.845 153.290 347.850 ;
        RECT 152.970 308.465 153.350 308.845 ;
        RECT 153.010 269.460 153.290 308.465 ;
        RECT 152.970 269.080 153.350 269.460 ;
        RECT 153.010 230.075 153.290 269.080 ;
        RECT 152.970 229.695 153.350 230.075 ;
        RECT 153.010 190.690 153.290 229.695 ;
        RECT 152.970 190.310 153.350 190.690 ;
        RECT 153.010 151.305 153.290 190.310 ;
        RECT 152.970 150.925 153.350 151.305 ;
        RECT 153.010 111.920 153.290 150.925 ;
        RECT 152.970 111.540 153.350 111.920 ;
        RECT 153.010 72.535 153.290 111.540 ;
        RECT 152.970 72.155 153.350 72.535 ;
        RECT 153.010 66.885 153.290 72.155 ;
    END
  END BIT_SEL[59]
  PIN BIT_SEL[60]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 152.370 379.455 152.650 382.085 ;
        RECT 152.330 379.075 152.710 379.455 ;
        RECT 152.370 340.070 152.650 379.075 ;
        RECT 152.330 339.690 152.710 340.070 ;
        RECT 152.370 300.685 152.650 339.690 ;
        RECT 152.330 300.305 152.710 300.685 ;
        RECT 152.370 261.300 152.650 300.305 ;
        RECT 152.330 260.920 152.710 261.300 ;
        RECT 152.370 221.915 152.650 260.920 ;
        RECT 152.330 221.535 152.710 221.915 ;
        RECT 152.370 182.530 152.650 221.535 ;
        RECT 152.330 182.150 152.710 182.530 ;
        RECT 152.370 143.145 152.650 182.150 ;
        RECT 152.330 142.765 152.710 143.145 ;
        RECT 152.370 103.760 152.650 142.765 ;
        RECT 152.330 103.380 152.710 103.760 ;
        RECT 152.370 66.885 152.650 103.380 ;
    END
  END BIT_SEL[60]
  PIN BIT_SEL[61]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 151.730 345.590 152.010 382.085 ;
        RECT 151.690 345.210 152.070 345.590 ;
        RECT 151.730 306.205 152.010 345.210 ;
        RECT 151.690 305.825 152.070 306.205 ;
        RECT 151.730 266.820 152.010 305.825 ;
        RECT 151.690 266.440 152.070 266.820 ;
        RECT 151.730 227.435 152.010 266.440 ;
        RECT 151.690 227.055 152.070 227.435 ;
        RECT 151.730 188.050 152.010 227.055 ;
        RECT 151.690 187.670 152.070 188.050 ;
        RECT 151.730 148.665 152.010 187.670 ;
        RECT 151.690 148.285 152.070 148.665 ;
        RECT 151.730 109.280 152.010 148.285 ;
        RECT 151.690 108.900 152.070 109.280 ;
        RECT 151.730 69.895 152.010 108.900 ;
        RECT 151.690 69.515 152.070 69.895 ;
        RECT 151.730 66.885 152.010 69.515 ;
    END
  END BIT_SEL[61]
  PIN BIT_SEL[62]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 151.090 381.295 151.370 382.085 ;
        RECT 151.050 380.915 151.430 381.295 ;
        RECT 151.090 341.910 151.370 380.915 ;
        RECT 151.050 341.530 151.430 341.910 ;
        RECT 151.090 302.525 151.370 341.530 ;
        RECT 151.050 302.145 151.430 302.525 ;
        RECT 151.090 263.140 151.370 302.145 ;
        RECT 151.050 262.760 151.430 263.140 ;
        RECT 151.090 223.755 151.370 262.760 ;
        RECT 151.050 223.375 151.430 223.755 ;
        RECT 151.090 184.370 151.370 223.375 ;
        RECT 151.050 183.990 151.430 184.370 ;
        RECT 151.090 144.985 151.370 183.990 ;
        RECT 151.050 144.605 151.430 144.985 ;
        RECT 151.090 105.600 151.370 144.605 ;
        RECT 151.050 105.220 151.430 105.600 ;
        RECT 151.090 66.885 151.370 105.220 ;
    END
  END BIT_SEL[62]
  PIN BIT_SEL[63]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 150.450 343.750 150.730 382.085 ;
        RECT 150.410 343.370 150.790 343.750 ;
        RECT 150.450 304.365 150.730 343.370 ;
        RECT 150.410 303.985 150.790 304.365 ;
        RECT 150.450 264.980 150.730 303.985 ;
        RECT 150.410 264.600 150.790 264.980 ;
        RECT 150.450 225.595 150.730 264.600 ;
        RECT 150.410 225.215 150.790 225.595 ;
        RECT 150.450 186.210 150.730 225.215 ;
        RECT 150.410 185.830 150.790 186.210 ;
        RECT 150.450 146.825 150.730 185.830 ;
        RECT 150.410 146.445 150.790 146.825 ;
        RECT 150.450 107.440 150.730 146.445 ;
        RECT 150.410 107.060 150.790 107.440 ;
        RECT 150.450 68.055 150.730 107.060 ;
        RECT 150.410 67.675 150.790 68.055 ;
        RECT 150.450 66.885 150.730 67.675 ;
    END
  END BIT_SEL[63]
  PIN BIT_SEL[46]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 118.640 381.295 118.920 382.085 ;
        RECT 118.600 380.915 118.980 381.295 ;
        RECT 118.640 341.910 118.920 380.915 ;
        RECT 118.600 341.530 118.980 341.910 ;
        RECT 118.640 302.525 118.920 341.530 ;
        RECT 118.600 302.145 118.980 302.525 ;
        RECT 118.640 263.140 118.920 302.145 ;
        RECT 118.600 262.760 118.980 263.140 ;
        RECT 118.640 223.755 118.920 262.760 ;
        RECT 118.600 223.375 118.980 223.755 ;
        RECT 118.640 184.370 118.920 223.375 ;
        RECT 118.600 183.990 118.980 184.370 ;
        RECT 118.640 144.985 118.920 183.990 ;
        RECT 118.600 144.605 118.980 144.985 ;
        RECT 118.640 105.600 118.920 144.605 ;
        RECT 118.600 105.220 118.980 105.600 ;
        RECT 118.640 66.885 118.920 105.220 ;
    END
  END BIT_SEL[46]
  PIN BIT_SEL[47]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 118.000 343.750 118.280 382.085 ;
        RECT 117.960 343.370 118.340 343.750 ;
        RECT 118.000 304.365 118.280 343.370 ;
        RECT 117.960 303.985 118.340 304.365 ;
        RECT 118.000 264.980 118.280 303.985 ;
        RECT 117.960 264.600 118.340 264.980 ;
        RECT 118.000 225.595 118.280 264.600 ;
        RECT 117.960 225.215 118.340 225.595 ;
        RECT 118.000 186.210 118.280 225.215 ;
        RECT 117.960 185.830 118.340 186.210 ;
        RECT 118.000 146.825 118.280 185.830 ;
        RECT 117.960 146.445 118.340 146.825 ;
        RECT 118.000 107.440 118.280 146.445 ;
        RECT 117.960 107.060 118.340 107.440 ;
        RECT 118.000 68.055 118.280 107.060 ;
        RECT 117.960 67.675 118.340 68.055 ;
        RECT 118.000 66.885 118.280 67.675 ;
    END
  END BIT_SEL[47]
  PIN BIT_SEL[16]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 95.150 366.805 95.430 382.085 ;
        RECT 95.110 366.425 95.490 366.805 ;
        RECT 95.150 327.420 95.430 366.425 ;
        RECT 95.110 327.040 95.490 327.420 ;
        RECT 95.150 288.035 95.430 327.040 ;
        RECT 95.110 287.655 95.490 288.035 ;
        RECT 95.150 248.650 95.430 287.655 ;
        RECT 95.110 248.270 95.490 248.650 ;
        RECT 95.150 209.265 95.430 248.270 ;
        RECT 95.110 208.885 95.490 209.265 ;
        RECT 95.150 169.880 95.430 208.885 ;
        RECT 95.110 169.500 95.490 169.880 ;
        RECT 95.150 130.495 95.430 169.500 ;
        RECT 95.110 130.115 95.490 130.495 ;
        RECT 95.150 91.110 95.430 130.115 ;
        RECT 95.110 90.730 95.490 91.110 ;
        RECT 95.150 66.885 95.430 90.730 ;
    END
  END BIT_SEL[16]
  PIN BIT_SEL[32]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 127.600 366.805 127.880 382.085 ;
        RECT 127.560 366.425 127.940 366.805 ;
        RECT 127.600 327.420 127.880 366.425 ;
        RECT 127.560 327.040 127.940 327.420 ;
        RECT 127.600 288.035 127.880 327.040 ;
        RECT 127.560 287.655 127.940 288.035 ;
        RECT 127.600 248.650 127.880 287.655 ;
        RECT 127.560 248.270 127.940 248.650 ;
        RECT 127.600 209.265 127.880 248.270 ;
        RECT 127.560 208.885 127.940 209.265 ;
        RECT 127.600 169.880 127.880 208.885 ;
        RECT 127.560 169.500 127.940 169.880 ;
        RECT 127.600 130.495 127.880 169.500 ;
        RECT 127.560 130.115 127.940 130.495 ;
        RECT 127.600 91.110 127.880 130.115 ;
        RECT 127.560 90.730 127.940 91.110 ;
        RECT 127.600 66.885 127.880 90.730 ;
    END
  END BIT_SEL[32]
  PIN BIT_SEL[33]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 126.960 358.240 127.240 382.085 ;
        RECT 126.920 357.860 127.300 358.240 ;
        RECT 126.960 318.855 127.240 357.860 ;
        RECT 126.920 318.475 127.300 318.855 ;
        RECT 126.960 279.470 127.240 318.475 ;
        RECT 126.920 279.090 127.300 279.470 ;
        RECT 126.960 240.085 127.240 279.090 ;
        RECT 126.920 239.705 127.300 240.085 ;
        RECT 126.960 200.700 127.240 239.705 ;
        RECT 126.920 200.320 127.300 200.700 ;
        RECT 126.960 161.315 127.240 200.320 ;
        RECT 126.920 160.935 127.300 161.315 ;
        RECT 126.960 121.930 127.240 160.935 ;
        RECT 126.920 121.550 127.300 121.930 ;
        RECT 126.960 82.545 127.240 121.550 ;
        RECT 126.920 82.165 127.300 82.545 ;
        RECT 126.960 66.885 127.240 82.165 ;
    END
  END BIT_SEL[33]
  PIN BIT_SEL[34]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 126.320 368.645 126.600 382.085 ;
        RECT 126.280 368.265 126.660 368.645 ;
        RECT 126.320 329.260 126.600 368.265 ;
        RECT 126.280 328.880 126.660 329.260 ;
        RECT 126.320 289.875 126.600 328.880 ;
        RECT 126.280 289.495 126.660 289.875 ;
        RECT 126.320 250.490 126.600 289.495 ;
        RECT 126.280 250.110 126.660 250.490 ;
        RECT 126.320 211.105 126.600 250.110 ;
        RECT 126.280 210.725 126.660 211.105 ;
        RECT 126.320 171.720 126.600 210.725 ;
        RECT 126.280 171.340 126.660 171.720 ;
        RECT 126.320 132.335 126.600 171.340 ;
        RECT 126.280 131.955 126.660 132.335 ;
        RECT 126.320 92.950 126.600 131.955 ;
        RECT 126.280 92.570 126.660 92.950 ;
        RECT 126.320 66.885 126.600 92.570 ;
    END
  END BIT_SEL[34]
  PIN BIT_SEL[35]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 125.680 356.400 125.960 382.085 ;
        RECT 125.640 356.020 126.020 356.400 ;
        RECT 125.680 317.015 125.960 356.020 ;
        RECT 125.640 316.635 126.020 317.015 ;
        RECT 125.680 277.630 125.960 316.635 ;
        RECT 125.640 277.250 126.020 277.630 ;
        RECT 125.680 238.245 125.960 277.250 ;
        RECT 125.640 237.865 126.020 238.245 ;
        RECT 125.680 198.860 125.960 237.865 ;
        RECT 125.640 198.480 126.020 198.860 ;
        RECT 125.680 159.475 125.960 198.480 ;
        RECT 125.640 159.095 126.020 159.475 ;
        RECT 125.680 120.090 125.960 159.095 ;
        RECT 125.640 119.710 126.020 120.090 ;
        RECT 125.680 80.705 125.960 119.710 ;
        RECT 125.640 80.325 126.020 80.705 ;
        RECT 125.680 66.885 125.960 80.325 ;
    END
  END BIT_SEL[35]
  PIN BIT_SEL[36]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 125.040 370.485 125.320 382.085 ;
        RECT 125.000 370.105 125.380 370.485 ;
        RECT 125.040 331.100 125.320 370.105 ;
        RECT 125.000 330.720 125.380 331.100 ;
        RECT 125.040 291.715 125.320 330.720 ;
        RECT 125.000 291.335 125.380 291.715 ;
        RECT 125.040 252.330 125.320 291.335 ;
        RECT 125.000 251.950 125.380 252.330 ;
        RECT 125.040 212.945 125.320 251.950 ;
        RECT 125.000 212.565 125.380 212.945 ;
        RECT 125.040 173.560 125.320 212.565 ;
        RECT 125.000 173.180 125.380 173.560 ;
        RECT 125.040 134.175 125.320 173.180 ;
        RECT 125.000 133.795 125.380 134.175 ;
        RECT 125.040 94.790 125.320 133.795 ;
        RECT 125.000 94.410 125.380 94.790 ;
        RECT 125.040 66.885 125.320 94.410 ;
    END
  END BIT_SEL[36]
  PIN BIT_SEL[37]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 124.400 354.555 124.680 382.085 ;
        RECT 124.360 354.175 124.740 354.555 ;
        RECT 124.400 315.170 124.680 354.175 ;
        RECT 124.360 314.790 124.740 315.170 ;
        RECT 124.400 275.785 124.680 314.790 ;
        RECT 124.360 275.405 124.740 275.785 ;
        RECT 124.400 236.400 124.680 275.405 ;
        RECT 124.360 236.020 124.740 236.400 ;
        RECT 124.400 197.015 124.680 236.020 ;
        RECT 124.360 196.635 124.740 197.015 ;
        RECT 124.400 157.630 124.680 196.635 ;
        RECT 124.360 157.250 124.740 157.630 ;
        RECT 124.400 118.245 124.680 157.250 ;
        RECT 124.360 117.865 124.740 118.245 ;
        RECT 124.400 78.860 124.680 117.865 ;
        RECT 124.360 78.480 124.740 78.860 ;
        RECT 124.400 66.885 124.680 78.480 ;
    END
  END BIT_SEL[37]
  PIN BIT_SEL[38]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 123.760 373.130 124.040 382.085 ;
        RECT 123.720 372.750 124.100 373.130 ;
        RECT 123.760 333.745 124.040 372.750 ;
        RECT 123.720 333.365 124.100 333.745 ;
        RECT 123.760 294.360 124.040 333.365 ;
        RECT 123.720 293.980 124.100 294.360 ;
        RECT 123.760 254.975 124.040 293.980 ;
        RECT 123.720 254.595 124.100 254.975 ;
        RECT 123.760 215.590 124.040 254.595 ;
        RECT 123.720 215.210 124.100 215.590 ;
        RECT 123.760 176.205 124.040 215.210 ;
        RECT 123.720 175.825 124.100 176.205 ;
        RECT 123.760 136.820 124.040 175.825 ;
        RECT 123.720 136.440 124.100 136.820 ;
        RECT 123.760 97.435 124.040 136.440 ;
        RECT 123.720 97.055 124.100 97.435 ;
        RECT 123.760 66.885 124.040 97.055 ;
    END
  END BIT_SEL[38]
  PIN BIT_SEL[39]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 123.120 351.915 123.400 382.085 ;
        RECT 123.080 351.535 123.460 351.915 ;
        RECT 123.120 312.530 123.400 351.535 ;
        RECT 123.080 312.150 123.460 312.530 ;
        RECT 123.120 273.145 123.400 312.150 ;
        RECT 123.080 272.765 123.460 273.145 ;
        RECT 123.120 233.760 123.400 272.765 ;
        RECT 123.080 233.380 123.460 233.760 ;
        RECT 123.120 194.375 123.400 233.380 ;
        RECT 123.080 193.995 123.460 194.375 ;
        RECT 123.120 154.990 123.400 193.995 ;
        RECT 123.080 154.610 123.460 154.990 ;
        RECT 123.120 115.605 123.400 154.610 ;
        RECT 123.080 115.225 123.460 115.605 ;
        RECT 123.120 76.220 123.400 115.225 ;
        RECT 123.080 75.840 123.460 76.220 ;
        RECT 123.120 66.885 123.400 75.840 ;
    END
  END BIT_SEL[39]
  PIN BIT_SEL[40]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 122.480 374.970 122.760 382.085 ;
        RECT 122.440 374.590 122.820 374.970 ;
        RECT 122.480 335.585 122.760 374.590 ;
        RECT 122.440 335.205 122.820 335.585 ;
        RECT 122.480 296.200 122.760 335.205 ;
        RECT 122.440 295.820 122.820 296.200 ;
        RECT 122.480 256.815 122.760 295.820 ;
        RECT 122.440 256.435 122.820 256.815 ;
        RECT 122.480 217.430 122.760 256.435 ;
        RECT 122.440 217.050 122.820 217.430 ;
        RECT 122.480 178.045 122.760 217.050 ;
        RECT 122.440 177.665 122.820 178.045 ;
        RECT 122.480 138.660 122.760 177.665 ;
        RECT 122.440 138.280 122.820 138.660 ;
        RECT 122.480 99.275 122.760 138.280 ;
        RECT 122.440 98.895 122.820 99.275 ;
        RECT 122.480 66.885 122.760 98.895 ;
    END
  END BIT_SEL[40]
  PIN BIT_SEL[41]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 121.840 350.075 122.120 382.085 ;
        RECT 121.800 349.695 122.180 350.075 ;
        RECT 121.840 310.690 122.120 349.695 ;
        RECT 121.800 310.310 122.180 310.690 ;
        RECT 121.840 271.305 122.120 310.310 ;
        RECT 121.800 270.925 122.180 271.305 ;
        RECT 121.840 231.920 122.120 270.925 ;
        RECT 121.800 231.540 122.180 231.920 ;
        RECT 121.840 192.535 122.120 231.540 ;
        RECT 121.800 192.155 122.180 192.535 ;
        RECT 121.840 153.150 122.120 192.155 ;
        RECT 121.800 152.770 122.180 153.150 ;
        RECT 121.840 113.765 122.120 152.770 ;
        RECT 121.800 113.385 122.180 113.765 ;
        RECT 121.840 74.380 122.120 113.385 ;
        RECT 121.800 74.000 122.180 74.380 ;
        RECT 121.840 66.885 122.120 74.000 ;
    END
  END BIT_SEL[41]
  PIN BIT_SEL[42]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 121.200 376.810 121.480 382.085 ;
        RECT 121.160 376.430 121.540 376.810 ;
        RECT 121.200 337.425 121.480 376.430 ;
        RECT 121.160 337.045 121.540 337.425 ;
        RECT 121.200 298.040 121.480 337.045 ;
        RECT 121.160 297.660 121.540 298.040 ;
        RECT 121.200 258.655 121.480 297.660 ;
        RECT 121.160 258.275 121.540 258.655 ;
        RECT 121.200 219.270 121.480 258.275 ;
        RECT 121.160 218.890 121.540 219.270 ;
        RECT 121.200 179.885 121.480 218.890 ;
        RECT 121.160 179.505 121.540 179.885 ;
        RECT 121.200 140.500 121.480 179.505 ;
        RECT 121.160 140.120 121.540 140.500 ;
        RECT 121.200 101.115 121.480 140.120 ;
        RECT 121.160 100.735 121.540 101.115 ;
        RECT 121.200 66.885 121.480 100.735 ;
    END
  END BIT_SEL[42]
  PIN BIT_SEL[43]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 120.560 348.230 120.840 382.085 ;
        RECT 120.520 347.850 120.900 348.230 ;
        RECT 120.560 308.845 120.840 347.850 ;
        RECT 120.520 308.465 120.900 308.845 ;
        RECT 120.560 269.460 120.840 308.465 ;
        RECT 120.520 269.080 120.900 269.460 ;
        RECT 120.560 230.075 120.840 269.080 ;
        RECT 120.520 229.695 120.900 230.075 ;
        RECT 120.560 190.690 120.840 229.695 ;
        RECT 120.520 190.310 120.900 190.690 ;
        RECT 120.560 151.305 120.840 190.310 ;
        RECT 120.520 150.925 120.900 151.305 ;
        RECT 120.560 111.920 120.840 150.925 ;
        RECT 120.520 111.540 120.900 111.920 ;
        RECT 120.560 72.535 120.840 111.540 ;
        RECT 120.520 72.155 120.900 72.535 ;
        RECT 120.560 66.885 120.840 72.155 ;
    END
  END BIT_SEL[43]
  PIN BIT_SEL[44]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 119.920 379.455 120.200 382.085 ;
        RECT 119.880 379.075 120.260 379.455 ;
        RECT 119.920 340.070 120.200 379.075 ;
        RECT 119.880 339.690 120.260 340.070 ;
        RECT 119.920 300.685 120.200 339.690 ;
        RECT 119.880 300.305 120.260 300.685 ;
        RECT 119.920 261.300 120.200 300.305 ;
        RECT 119.880 260.920 120.260 261.300 ;
        RECT 119.920 221.915 120.200 260.920 ;
        RECT 119.880 221.535 120.260 221.915 ;
        RECT 119.920 182.530 120.200 221.535 ;
        RECT 119.880 182.150 120.260 182.530 ;
        RECT 119.920 143.145 120.200 182.150 ;
        RECT 119.880 142.765 120.260 143.145 ;
        RECT 119.920 103.760 120.200 142.765 ;
        RECT 119.880 103.380 120.260 103.760 ;
        RECT 119.920 66.885 120.200 103.380 ;
    END
  END BIT_SEL[44]
  PIN BIT_SEL[45]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 119.280 345.590 119.560 382.085 ;
        RECT 119.240 345.210 119.620 345.590 ;
        RECT 119.280 306.205 119.560 345.210 ;
        RECT 119.240 305.825 119.620 306.205 ;
        RECT 119.280 266.820 119.560 305.825 ;
        RECT 119.240 266.440 119.620 266.820 ;
        RECT 119.280 227.435 119.560 266.440 ;
        RECT 119.240 227.055 119.620 227.435 ;
        RECT 119.280 188.050 119.560 227.055 ;
        RECT 119.240 187.670 119.620 188.050 ;
        RECT 119.280 148.665 119.560 187.670 ;
        RECT 119.240 148.285 119.620 148.665 ;
        RECT 119.280 109.280 119.560 148.285 ;
        RECT 119.240 108.900 119.620 109.280 ;
        RECT 119.280 69.895 119.560 108.900 ;
        RECT 119.240 69.515 119.620 69.895 ;
        RECT 119.280 66.885 119.560 69.515 ;
    END
  END BIT_SEL[45]
  PIN BIT_SEL[0]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 62.700 366.805 62.980 382.085 ;
        RECT 62.660 366.425 63.040 366.805 ;
        RECT 62.700 327.420 62.980 366.425 ;
        RECT 62.660 327.040 63.040 327.420 ;
        RECT 62.700 288.035 62.980 327.040 ;
        RECT 62.660 287.655 63.040 288.035 ;
        RECT 62.700 248.650 62.980 287.655 ;
        RECT 62.660 248.270 63.040 248.650 ;
        RECT 62.700 209.265 62.980 248.270 ;
        RECT 62.660 208.885 63.040 209.265 ;
        RECT 62.700 169.880 62.980 208.885 ;
        RECT 62.660 169.500 63.040 169.880 ;
        RECT 62.700 130.495 62.980 169.500 ;
        RECT 62.660 130.115 63.040 130.495 ;
        RECT 62.700 91.110 62.980 130.115 ;
        RECT 62.660 90.730 63.040 91.110 ;
        RECT 62.700 66.885 62.980 90.730 ;
    END
  END BIT_SEL[0]
  PIN BIT_SEL[1]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 62.060 358.240 62.340 382.085 ;
        RECT 62.020 357.860 62.400 358.240 ;
        RECT 62.060 318.855 62.340 357.860 ;
        RECT 62.020 318.475 62.400 318.855 ;
        RECT 62.060 279.470 62.340 318.475 ;
        RECT 62.020 279.090 62.400 279.470 ;
        RECT 62.060 240.085 62.340 279.090 ;
        RECT 62.020 239.705 62.400 240.085 ;
        RECT 62.060 200.700 62.340 239.705 ;
        RECT 62.020 200.320 62.400 200.700 ;
        RECT 62.060 161.315 62.340 200.320 ;
        RECT 62.020 160.935 62.400 161.315 ;
        RECT 62.060 121.930 62.340 160.935 ;
        RECT 62.020 121.550 62.400 121.930 ;
        RECT 62.060 82.545 62.340 121.550 ;
        RECT 62.020 82.165 62.400 82.545 ;
        RECT 62.060 66.885 62.340 82.165 ;
    END
  END BIT_SEL[1]
  PIN BIT_SEL[2]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 61.420 368.645 61.700 382.085 ;
        RECT 61.380 368.265 61.760 368.645 ;
        RECT 61.420 329.260 61.700 368.265 ;
        RECT 61.380 328.880 61.760 329.260 ;
        RECT 61.420 289.875 61.700 328.880 ;
        RECT 61.380 289.495 61.760 289.875 ;
        RECT 61.420 250.490 61.700 289.495 ;
        RECT 61.380 250.110 61.760 250.490 ;
        RECT 61.420 211.105 61.700 250.110 ;
        RECT 61.380 210.725 61.760 211.105 ;
        RECT 61.420 171.720 61.700 210.725 ;
        RECT 61.380 171.340 61.760 171.720 ;
        RECT 61.420 132.335 61.700 171.340 ;
        RECT 61.380 131.955 61.760 132.335 ;
        RECT 61.420 92.950 61.700 131.955 ;
        RECT 61.380 92.570 61.760 92.950 ;
        RECT 61.420 66.885 61.700 92.570 ;
    END
  END BIT_SEL[2]
  PIN BIT_SEL[3]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 60.780 356.400 61.060 382.085 ;
        RECT 60.740 356.020 61.120 356.400 ;
        RECT 60.780 317.015 61.060 356.020 ;
        RECT 60.740 316.635 61.120 317.015 ;
        RECT 60.780 277.630 61.060 316.635 ;
        RECT 60.740 277.250 61.120 277.630 ;
        RECT 60.780 238.245 61.060 277.250 ;
        RECT 60.740 237.865 61.120 238.245 ;
        RECT 60.780 198.860 61.060 237.865 ;
        RECT 60.740 198.480 61.120 198.860 ;
        RECT 60.780 159.475 61.060 198.480 ;
        RECT 60.740 159.095 61.120 159.475 ;
        RECT 60.780 120.090 61.060 159.095 ;
        RECT 60.740 119.710 61.120 120.090 ;
        RECT 60.780 80.705 61.060 119.710 ;
        RECT 60.740 80.325 61.120 80.705 ;
        RECT 60.780 66.885 61.060 80.325 ;
    END
  END BIT_SEL[3]
  PIN BIT_SEL[4]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 60.140 370.485 60.420 382.085 ;
        RECT 60.100 370.105 60.480 370.485 ;
        RECT 60.140 331.100 60.420 370.105 ;
        RECT 60.100 330.720 60.480 331.100 ;
        RECT 60.140 291.715 60.420 330.720 ;
        RECT 60.100 291.335 60.480 291.715 ;
        RECT 60.140 252.330 60.420 291.335 ;
        RECT 60.100 251.950 60.480 252.330 ;
        RECT 60.140 212.945 60.420 251.950 ;
        RECT 60.100 212.565 60.480 212.945 ;
        RECT 60.140 173.560 60.420 212.565 ;
        RECT 60.100 173.180 60.480 173.560 ;
        RECT 60.140 134.175 60.420 173.180 ;
        RECT 60.100 133.795 60.480 134.175 ;
        RECT 60.140 94.790 60.420 133.795 ;
        RECT 60.100 94.410 60.480 94.790 ;
        RECT 60.140 66.885 60.420 94.410 ;
    END
  END BIT_SEL[4]
  PIN BIT_SEL[17]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 94.510 358.240 94.790 382.085 ;
        RECT 94.470 357.860 94.850 358.240 ;
        RECT 94.510 318.855 94.790 357.860 ;
        RECT 94.470 318.475 94.850 318.855 ;
        RECT 94.510 279.470 94.790 318.475 ;
        RECT 94.470 279.090 94.850 279.470 ;
        RECT 94.510 240.085 94.790 279.090 ;
        RECT 94.470 239.705 94.850 240.085 ;
        RECT 94.510 200.700 94.790 239.705 ;
        RECT 94.470 200.320 94.850 200.700 ;
        RECT 94.510 161.315 94.790 200.320 ;
        RECT 94.470 160.935 94.850 161.315 ;
        RECT 94.510 121.930 94.790 160.935 ;
        RECT 94.470 121.550 94.850 121.930 ;
        RECT 94.510 82.545 94.790 121.550 ;
        RECT 94.470 82.165 94.850 82.545 ;
        RECT 94.510 66.885 94.790 82.165 ;
    END
  END BIT_SEL[17]
  PIN BIT_SEL[18]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 93.870 368.645 94.150 382.085 ;
        RECT 93.830 368.265 94.210 368.645 ;
        RECT 93.870 329.260 94.150 368.265 ;
        RECT 93.830 328.880 94.210 329.260 ;
        RECT 93.870 289.875 94.150 328.880 ;
        RECT 93.830 289.495 94.210 289.875 ;
        RECT 93.870 250.490 94.150 289.495 ;
        RECT 93.830 250.110 94.210 250.490 ;
        RECT 93.870 211.105 94.150 250.110 ;
        RECT 93.830 210.725 94.210 211.105 ;
        RECT 93.870 171.720 94.150 210.725 ;
        RECT 93.830 171.340 94.210 171.720 ;
        RECT 93.870 132.335 94.150 171.340 ;
        RECT 93.830 131.955 94.210 132.335 ;
        RECT 93.870 92.950 94.150 131.955 ;
        RECT 93.830 92.570 94.210 92.950 ;
        RECT 93.870 66.885 94.150 92.570 ;
    END
  END BIT_SEL[18]
  PIN BIT_SEL[19]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 93.230 356.400 93.510 382.085 ;
        RECT 93.190 356.020 93.570 356.400 ;
        RECT 93.230 317.015 93.510 356.020 ;
        RECT 93.190 316.635 93.570 317.015 ;
        RECT 93.230 277.630 93.510 316.635 ;
        RECT 93.190 277.250 93.570 277.630 ;
        RECT 93.230 238.245 93.510 277.250 ;
        RECT 93.190 237.865 93.570 238.245 ;
        RECT 93.230 198.860 93.510 237.865 ;
        RECT 93.190 198.480 93.570 198.860 ;
        RECT 93.230 159.475 93.510 198.480 ;
        RECT 93.190 159.095 93.570 159.475 ;
        RECT 93.230 120.090 93.510 159.095 ;
        RECT 93.190 119.710 93.570 120.090 ;
        RECT 93.230 80.705 93.510 119.710 ;
        RECT 93.190 80.325 93.570 80.705 ;
        RECT 93.230 66.885 93.510 80.325 ;
    END
  END BIT_SEL[19]
  PIN BIT_SEL[20]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 92.590 370.485 92.870 382.085 ;
        RECT 92.550 370.105 92.930 370.485 ;
        RECT 92.590 331.100 92.870 370.105 ;
        RECT 92.550 330.720 92.930 331.100 ;
        RECT 92.590 291.715 92.870 330.720 ;
        RECT 92.550 291.335 92.930 291.715 ;
        RECT 92.590 252.330 92.870 291.335 ;
        RECT 92.550 251.950 92.930 252.330 ;
        RECT 92.590 212.945 92.870 251.950 ;
        RECT 92.550 212.565 92.930 212.945 ;
        RECT 92.590 173.560 92.870 212.565 ;
        RECT 92.550 173.180 92.930 173.560 ;
        RECT 92.590 134.175 92.870 173.180 ;
        RECT 92.550 133.795 92.930 134.175 ;
        RECT 92.590 94.790 92.870 133.795 ;
        RECT 92.550 94.410 92.930 94.790 ;
        RECT 92.590 66.885 92.870 94.410 ;
    END
  END BIT_SEL[20]
  PIN BIT_SEL[21]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 91.950 354.555 92.230 382.085 ;
        RECT 91.910 354.175 92.290 354.555 ;
        RECT 91.950 315.170 92.230 354.175 ;
        RECT 91.910 314.790 92.290 315.170 ;
        RECT 91.950 275.785 92.230 314.790 ;
        RECT 91.910 275.405 92.290 275.785 ;
        RECT 91.950 236.400 92.230 275.405 ;
        RECT 91.910 236.020 92.290 236.400 ;
        RECT 91.950 197.015 92.230 236.020 ;
        RECT 91.910 196.635 92.290 197.015 ;
        RECT 91.950 157.630 92.230 196.635 ;
        RECT 91.910 157.250 92.290 157.630 ;
        RECT 91.950 118.245 92.230 157.250 ;
        RECT 91.910 117.865 92.290 118.245 ;
        RECT 91.950 78.860 92.230 117.865 ;
        RECT 91.910 78.480 92.290 78.860 ;
        RECT 91.950 66.885 92.230 78.480 ;
    END
  END BIT_SEL[21]
  PIN BIT_SEL[22]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 91.310 373.130 91.590 382.085 ;
        RECT 91.270 372.750 91.650 373.130 ;
        RECT 91.310 333.745 91.590 372.750 ;
        RECT 91.270 333.365 91.650 333.745 ;
        RECT 91.310 294.360 91.590 333.365 ;
        RECT 91.270 293.980 91.650 294.360 ;
        RECT 91.310 254.975 91.590 293.980 ;
        RECT 91.270 254.595 91.650 254.975 ;
        RECT 91.310 215.590 91.590 254.595 ;
        RECT 91.270 215.210 91.650 215.590 ;
        RECT 91.310 176.205 91.590 215.210 ;
        RECT 91.270 175.825 91.650 176.205 ;
        RECT 91.310 136.820 91.590 175.825 ;
        RECT 91.270 136.440 91.650 136.820 ;
        RECT 91.310 97.435 91.590 136.440 ;
        RECT 91.270 97.055 91.650 97.435 ;
        RECT 91.310 66.885 91.590 97.055 ;
    END
  END BIT_SEL[22]
  PIN BIT_SEL[23]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 90.670 351.915 90.950 382.085 ;
        RECT 90.630 351.535 91.010 351.915 ;
        RECT 90.670 312.530 90.950 351.535 ;
        RECT 90.630 312.150 91.010 312.530 ;
        RECT 90.670 273.145 90.950 312.150 ;
        RECT 90.630 272.765 91.010 273.145 ;
        RECT 90.670 233.760 90.950 272.765 ;
        RECT 90.630 233.380 91.010 233.760 ;
        RECT 90.670 194.375 90.950 233.380 ;
        RECT 90.630 193.995 91.010 194.375 ;
        RECT 90.670 154.990 90.950 193.995 ;
        RECT 90.630 154.610 91.010 154.990 ;
        RECT 90.670 115.605 90.950 154.610 ;
        RECT 90.630 115.225 91.010 115.605 ;
        RECT 90.670 76.220 90.950 115.225 ;
        RECT 90.630 75.840 91.010 76.220 ;
        RECT 90.670 66.885 90.950 75.840 ;
    END
  END BIT_SEL[23]
  PIN BIT_SEL[24]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 90.030 374.970 90.310 382.085 ;
        RECT 89.990 374.590 90.370 374.970 ;
        RECT 90.030 335.585 90.310 374.590 ;
        RECT 89.990 335.205 90.370 335.585 ;
        RECT 90.030 296.200 90.310 335.205 ;
        RECT 89.990 295.820 90.370 296.200 ;
        RECT 90.030 256.815 90.310 295.820 ;
        RECT 89.990 256.435 90.370 256.815 ;
        RECT 90.030 217.430 90.310 256.435 ;
        RECT 89.990 217.050 90.370 217.430 ;
        RECT 90.030 178.045 90.310 217.050 ;
        RECT 89.990 177.665 90.370 178.045 ;
        RECT 90.030 138.660 90.310 177.665 ;
        RECT 89.990 138.280 90.370 138.660 ;
        RECT 90.030 99.275 90.310 138.280 ;
        RECT 89.990 98.895 90.370 99.275 ;
        RECT 90.030 66.885 90.310 98.895 ;
    END
  END BIT_SEL[24]
  PIN BIT_SEL[25]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 89.390 350.075 89.670 382.085 ;
        RECT 89.350 349.695 89.730 350.075 ;
        RECT 89.390 310.690 89.670 349.695 ;
        RECT 89.350 310.310 89.730 310.690 ;
        RECT 89.390 271.305 89.670 310.310 ;
        RECT 89.350 270.925 89.730 271.305 ;
        RECT 89.390 231.920 89.670 270.925 ;
        RECT 89.350 231.540 89.730 231.920 ;
        RECT 89.390 192.535 89.670 231.540 ;
        RECT 89.350 192.155 89.730 192.535 ;
        RECT 89.390 153.150 89.670 192.155 ;
        RECT 89.350 152.770 89.730 153.150 ;
        RECT 89.390 113.765 89.670 152.770 ;
        RECT 89.350 113.385 89.730 113.765 ;
        RECT 89.390 74.380 89.670 113.385 ;
        RECT 89.350 74.000 89.730 74.380 ;
        RECT 89.390 66.885 89.670 74.000 ;
    END
  END BIT_SEL[25]
  PIN BIT_SEL[26]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 88.750 376.810 89.030 382.085 ;
        RECT 88.710 376.430 89.090 376.810 ;
        RECT 88.750 337.425 89.030 376.430 ;
        RECT 88.710 337.045 89.090 337.425 ;
        RECT 88.750 298.040 89.030 337.045 ;
        RECT 88.710 297.660 89.090 298.040 ;
        RECT 88.750 258.655 89.030 297.660 ;
        RECT 88.710 258.275 89.090 258.655 ;
        RECT 88.750 219.270 89.030 258.275 ;
        RECT 88.710 218.890 89.090 219.270 ;
        RECT 88.750 179.885 89.030 218.890 ;
        RECT 88.710 179.505 89.090 179.885 ;
        RECT 88.750 140.500 89.030 179.505 ;
        RECT 88.710 140.120 89.090 140.500 ;
        RECT 88.750 101.115 89.030 140.120 ;
        RECT 88.710 100.735 89.090 101.115 ;
        RECT 88.750 66.885 89.030 100.735 ;
    END
  END BIT_SEL[26]
  PIN BIT_SEL[27]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 88.110 348.230 88.390 382.085 ;
        RECT 88.070 347.850 88.450 348.230 ;
        RECT 88.110 308.845 88.390 347.850 ;
        RECT 88.070 308.465 88.450 308.845 ;
        RECT 88.110 269.460 88.390 308.465 ;
        RECT 88.070 269.080 88.450 269.460 ;
        RECT 88.110 230.075 88.390 269.080 ;
        RECT 88.070 229.695 88.450 230.075 ;
        RECT 88.110 190.690 88.390 229.695 ;
        RECT 88.070 190.310 88.450 190.690 ;
        RECT 88.110 151.305 88.390 190.310 ;
        RECT 88.070 150.925 88.450 151.305 ;
        RECT 88.110 111.920 88.390 150.925 ;
        RECT 88.070 111.540 88.450 111.920 ;
        RECT 88.110 72.535 88.390 111.540 ;
        RECT 88.070 72.155 88.450 72.535 ;
        RECT 88.110 66.885 88.390 72.155 ;
    END
  END BIT_SEL[27]
  PIN BIT_SEL[28]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 87.470 379.455 87.750 382.085 ;
        RECT 87.430 379.075 87.810 379.455 ;
        RECT 87.470 340.070 87.750 379.075 ;
        RECT 87.430 339.690 87.810 340.070 ;
        RECT 87.470 300.685 87.750 339.690 ;
        RECT 87.430 300.305 87.810 300.685 ;
        RECT 87.470 261.300 87.750 300.305 ;
        RECT 87.430 260.920 87.810 261.300 ;
        RECT 87.470 221.915 87.750 260.920 ;
        RECT 87.430 221.535 87.810 221.915 ;
        RECT 87.470 182.530 87.750 221.535 ;
        RECT 87.430 182.150 87.810 182.530 ;
        RECT 87.470 143.145 87.750 182.150 ;
        RECT 87.430 142.765 87.810 143.145 ;
        RECT 87.470 103.760 87.750 142.765 ;
        RECT 87.430 103.380 87.810 103.760 ;
        RECT 87.470 66.885 87.750 103.380 ;
    END
  END BIT_SEL[28]
  PIN BIT_SEL[29]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 86.830 345.590 87.110 382.085 ;
        RECT 86.790 345.210 87.170 345.590 ;
        RECT 86.830 306.205 87.110 345.210 ;
        RECT 86.790 305.825 87.170 306.205 ;
        RECT 86.830 266.820 87.110 305.825 ;
        RECT 86.790 266.440 87.170 266.820 ;
        RECT 86.830 227.435 87.110 266.440 ;
        RECT 86.790 227.055 87.170 227.435 ;
        RECT 86.830 188.050 87.110 227.055 ;
        RECT 86.790 187.670 87.170 188.050 ;
        RECT 86.830 148.665 87.110 187.670 ;
        RECT 86.790 148.285 87.170 148.665 ;
        RECT 86.830 109.280 87.110 148.285 ;
        RECT 86.790 108.900 87.170 109.280 ;
        RECT 86.830 69.895 87.110 108.900 ;
        RECT 86.790 69.515 87.170 69.895 ;
        RECT 86.830 66.885 87.110 69.515 ;
    END
  END BIT_SEL[29]
  PIN BIT_SEL[30]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 86.190 381.295 86.470 382.085 ;
        RECT 86.150 380.915 86.530 381.295 ;
        RECT 86.190 341.910 86.470 380.915 ;
        RECT 86.150 341.530 86.530 341.910 ;
        RECT 86.190 302.525 86.470 341.530 ;
        RECT 86.150 302.145 86.530 302.525 ;
        RECT 86.190 263.140 86.470 302.145 ;
        RECT 86.150 262.760 86.530 263.140 ;
        RECT 86.190 223.755 86.470 262.760 ;
        RECT 86.150 223.375 86.530 223.755 ;
        RECT 86.190 184.370 86.470 223.375 ;
        RECT 86.150 183.990 86.530 184.370 ;
        RECT 86.190 144.985 86.470 183.990 ;
        RECT 86.150 144.605 86.530 144.985 ;
        RECT 86.190 105.600 86.470 144.605 ;
        RECT 86.150 105.220 86.530 105.600 ;
        RECT 86.190 66.885 86.470 105.220 ;
    END
  END BIT_SEL[30]
  PIN BIT_SEL[31]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 85.550 343.750 85.830 382.085 ;
        RECT 85.510 343.370 85.890 343.750 ;
        RECT 85.550 304.365 85.830 343.370 ;
        RECT 85.510 303.985 85.890 304.365 ;
        RECT 85.550 264.980 85.830 303.985 ;
        RECT 85.510 264.600 85.890 264.980 ;
        RECT 85.550 225.595 85.830 264.600 ;
        RECT 85.510 225.215 85.890 225.595 ;
        RECT 85.550 186.210 85.830 225.215 ;
        RECT 85.510 185.830 85.890 186.210 ;
        RECT 85.550 146.825 85.830 185.830 ;
        RECT 85.510 146.445 85.890 146.825 ;
        RECT 85.550 107.440 85.830 146.445 ;
        RECT 85.510 107.060 85.890 107.440 ;
        RECT 85.550 68.055 85.830 107.060 ;
        RECT 85.510 67.675 85.890 68.055 ;
        RECT 85.550 66.885 85.830 67.675 ;
    END
  END BIT_SEL[31]
  PIN BIT_SEL[5]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 59.500 354.555 59.780 382.085 ;
        RECT 59.460 354.175 59.840 354.555 ;
        RECT 59.500 315.170 59.780 354.175 ;
        RECT 59.460 314.790 59.840 315.170 ;
        RECT 59.500 275.785 59.780 314.790 ;
        RECT 59.460 275.405 59.840 275.785 ;
        RECT 59.500 236.400 59.780 275.405 ;
        RECT 59.460 236.020 59.840 236.400 ;
        RECT 59.500 197.015 59.780 236.020 ;
        RECT 59.460 196.635 59.840 197.015 ;
        RECT 59.500 157.630 59.780 196.635 ;
        RECT 59.460 157.250 59.840 157.630 ;
        RECT 59.500 118.245 59.780 157.250 ;
        RECT 59.460 117.865 59.840 118.245 ;
        RECT 59.500 78.860 59.780 117.865 ;
        RECT 59.460 78.480 59.840 78.860 ;
        RECT 59.500 66.885 59.780 78.480 ;
    END
  END BIT_SEL[5]
  PIN BIT_SEL[6]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 58.860 373.130 59.140 382.085 ;
        RECT 58.820 372.750 59.200 373.130 ;
        RECT 58.860 333.745 59.140 372.750 ;
        RECT 58.820 333.365 59.200 333.745 ;
        RECT 58.860 294.360 59.140 333.365 ;
        RECT 58.820 293.980 59.200 294.360 ;
        RECT 58.860 254.975 59.140 293.980 ;
        RECT 58.820 254.595 59.200 254.975 ;
        RECT 58.860 215.590 59.140 254.595 ;
        RECT 58.820 215.210 59.200 215.590 ;
        RECT 58.860 176.205 59.140 215.210 ;
        RECT 58.820 175.825 59.200 176.205 ;
        RECT 58.860 136.820 59.140 175.825 ;
        RECT 58.820 136.440 59.200 136.820 ;
        RECT 58.860 97.435 59.140 136.440 ;
        RECT 58.820 97.055 59.200 97.435 ;
        RECT 58.860 66.885 59.140 97.055 ;
    END
  END BIT_SEL[6]
  PIN BIT_SEL[7]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 58.220 351.915 58.500 382.085 ;
        RECT 58.180 351.535 58.560 351.915 ;
        RECT 58.220 312.530 58.500 351.535 ;
        RECT 58.180 312.150 58.560 312.530 ;
        RECT 58.220 273.145 58.500 312.150 ;
        RECT 58.180 272.765 58.560 273.145 ;
        RECT 58.220 233.760 58.500 272.765 ;
        RECT 58.180 233.380 58.560 233.760 ;
        RECT 58.220 194.375 58.500 233.380 ;
        RECT 58.180 193.995 58.560 194.375 ;
        RECT 58.220 154.990 58.500 193.995 ;
        RECT 58.180 154.610 58.560 154.990 ;
        RECT 58.220 115.605 58.500 154.610 ;
        RECT 58.180 115.225 58.560 115.605 ;
        RECT 58.220 76.220 58.500 115.225 ;
        RECT 58.180 75.840 58.560 76.220 ;
        RECT 58.220 66.885 58.500 75.840 ;
    END
  END BIT_SEL[7]
  PIN BIT_SEL[8]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 57.580 374.970 57.860 382.085 ;
        RECT 57.540 374.590 57.920 374.970 ;
        RECT 57.580 335.585 57.860 374.590 ;
        RECT 57.540 335.205 57.920 335.585 ;
        RECT 57.580 296.200 57.860 335.205 ;
        RECT 57.540 295.820 57.920 296.200 ;
        RECT 57.580 256.815 57.860 295.820 ;
        RECT 57.540 256.435 57.920 256.815 ;
        RECT 57.580 217.430 57.860 256.435 ;
        RECT 57.540 217.050 57.920 217.430 ;
        RECT 57.580 178.045 57.860 217.050 ;
        RECT 57.540 177.665 57.920 178.045 ;
        RECT 57.580 138.660 57.860 177.665 ;
        RECT 57.540 138.280 57.920 138.660 ;
        RECT 57.580 99.275 57.860 138.280 ;
        RECT 57.540 98.895 57.920 99.275 ;
        RECT 57.580 66.885 57.860 98.895 ;
    END
  END BIT_SEL[8]
  PIN BIT_SEL[9]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 56.940 350.075 57.220 382.085 ;
        RECT 56.900 349.695 57.280 350.075 ;
        RECT 56.940 310.690 57.220 349.695 ;
        RECT 56.900 310.310 57.280 310.690 ;
        RECT 56.940 271.305 57.220 310.310 ;
        RECT 56.900 270.925 57.280 271.305 ;
        RECT 56.940 231.920 57.220 270.925 ;
        RECT 56.900 231.540 57.280 231.920 ;
        RECT 56.940 192.535 57.220 231.540 ;
        RECT 56.900 192.155 57.280 192.535 ;
        RECT 56.940 153.150 57.220 192.155 ;
        RECT 56.900 152.770 57.280 153.150 ;
        RECT 56.940 113.765 57.220 152.770 ;
        RECT 56.900 113.385 57.280 113.765 ;
        RECT 56.940 74.380 57.220 113.385 ;
        RECT 56.900 74.000 57.280 74.380 ;
        RECT 56.940 66.885 57.220 74.000 ;
    END
  END BIT_SEL[9]
  PIN BIT_SEL[10]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 56.300 376.810 56.580 382.085 ;
        RECT 56.260 376.430 56.640 376.810 ;
        RECT 56.300 337.425 56.580 376.430 ;
        RECT 56.260 337.045 56.640 337.425 ;
        RECT 56.300 298.040 56.580 337.045 ;
        RECT 56.260 297.660 56.640 298.040 ;
        RECT 56.300 258.655 56.580 297.660 ;
        RECT 56.260 258.275 56.640 258.655 ;
        RECT 56.300 219.270 56.580 258.275 ;
        RECT 56.260 218.890 56.640 219.270 ;
        RECT 56.300 179.885 56.580 218.890 ;
        RECT 56.260 179.505 56.640 179.885 ;
        RECT 56.300 140.500 56.580 179.505 ;
        RECT 56.260 140.120 56.640 140.500 ;
        RECT 56.300 101.115 56.580 140.120 ;
        RECT 56.260 100.735 56.640 101.115 ;
        RECT 56.300 66.885 56.580 100.735 ;
    END
  END BIT_SEL[10]
  PIN BIT_SEL[11]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 55.660 348.230 55.940 382.085 ;
        RECT 55.620 347.850 56.000 348.230 ;
        RECT 55.660 308.845 55.940 347.850 ;
        RECT 55.620 308.465 56.000 308.845 ;
        RECT 55.660 269.460 55.940 308.465 ;
        RECT 55.620 269.080 56.000 269.460 ;
        RECT 55.660 230.075 55.940 269.080 ;
        RECT 55.620 229.695 56.000 230.075 ;
        RECT 55.660 190.690 55.940 229.695 ;
        RECT 55.620 190.310 56.000 190.690 ;
        RECT 55.660 151.305 55.940 190.310 ;
        RECT 55.620 150.925 56.000 151.305 ;
        RECT 55.660 111.920 55.940 150.925 ;
        RECT 55.620 111.540 56.000 111.920 ;
        RECT 55.660 72.535 55.940 111.540 ;
        RECT 55.620 72.155 56.000 72.535 ;
        RECT 55.660 66.885 55.940 72.155 ;
    END
  END BIT_SEL[11]
  PIN BIT_SEL[12]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 55.020 379.455 55.300 382.085 ;
        RECT 54.980 379.075 55.360 379.455 ;
        RECT 55.020 340.070 55.300 379.075 ;
        RECT 54.980 339.690 55.360 340.070 ;
        RECT 55.020 300.685 55.300 339.690 ;
        RECT 54.980 300.305 55.360 300.685 ;
        RECT 55.020 261.300 55.300 300.305 ;
        RECT 54.980 260.920 55.360 261.300 ;
        RECT 55.020 221.915 55.300 260.920 ;
        RECT 54.980 221.535 55.360 221.915 ;
        RECT 55.020 182.530 55.300 221.535 ;
        RECT 54.980 182.150 55.360 182.530 ;
        RECT 55.020 143.145 55.300 182.150 ;
        RECT 54.980 142.765 55.360 143.145 ;
        RECT 55.020 103.760 55.300 142.765 ;
        RECT 54.980 103.380 55.360 103.760 ;
        RECT 55.020 66.885 55.300 103.380 ;
    END
  END BIT_SEL[12]
  PIN BIT_SEL[13]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 54.380 345.590 54.660 382.085 ;
        RECT 54.340 345.210 54.720 345.590 ;
        RECT 54.380 306.205 54.660 345.210 ;
        RECT 54.340 305.825 54.720 306.205 ;
        RECT 54.380 266.820 54.660 305.825 ;
        RECT 54.340 266.440 54.720 266.820 ;
        RECT 54.380 227.435 54.660 266.440 ;
        RECT 54.340 227.055 54.720 227.435 ;
        RECT 54.380 188.050 54.660 227.055 ;
        RECT 54.340 187.670 54.720 188.050 ;
        RECT 54.380 148.665 54.660 187.670 ;
        RECT 54.340 148.285 54.720 148.665 ;
        RECT 54.380 109.280 54.660 148.285 ;
        RECT 54.340 108.900 54.720 109.280 ;
        RECT 54.380 69.895 54.660 108.900 ;
        RECT 54.340 69.515 54.720 69.895 ;
        RECT 54.380 66.885 54.660 69.515 ;
    END
  END BIT_SEL[13]
  PIN BIT_SEL[14]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 53.740 381.295 54.020 382.085 ;
        RECT 53.700 380.915 54.080 381.295 ;
        RECT 53.740 341.910 54.020 380.915 ;
        RECT 53.700 341.530 54.080 341.910 ;
        RECT 53.740 302.525 54.020 341.530 ;
        RECT 53.700 302.145 54.080 302.525 ;
        RECT 53.740 263.140 54.020 302.145 ;
        RECT 53.700 262.760 54.080 263.140 ;
        RECT 53.740 223.755 54.020 262.760 ;
        RECT 53.700 223.375 54.080 223.755 ;
        RECT 53.740 184.370 54.020 223.375 ;
        RECT 53.700 183.990 54.080 184.370 ;
        RECT 53.740 144.985 54.020 183.990 ;
        RECT 53.700 144.605 54.080 144.985 ;
        RECT 53.740 105.600 54.020 144.605 ;
        RECT 53.700 105.220 54.080 105.600 ;
        RECT 53.740 66.885 54.020 105.220 ;
    END
  END BIT_SEL[14]
  PIN BIT_SEL[15]
    ANTENNAGATEAREA 146.399994 ;
    PORT
      LAYER Metal4 ;
        RECT 53.100 343.750 53.380 382.085 ;
        RECT 53.060 343.370 53.440 343.750 ;
        RECT 53.100 304.365 53.380 343.370 ;
        RECT 53.060 303.985 53.440 304.365 ;
        RECT 53.100 264.980 53.380 303.985 ;
        RECT 53.060 264.600 53.440 264.980 ;
        RECT 53.100 225.595 53.380 264.600 ;
        RECT 53.060 225.215 53.440 225.595 ;
        RECT 53.100 186.210 53.380 225.215 ;
        RECT 53.060 185.830 53.440 186.210 ;
        RECT 53.100 146.825 53.380 185.830 ;
        RECT 53.060 146.445 53.440 146.825 ;
        RECT 53.100 107.440 53.380 146.445 ;
        RECT 53.060 107.060 53.440 107.440 ;
        RECT 53.100 68.055 53.380 107.060 ;
        RECT 53.060 67.675 53.440 68.055 ;
        RECT 53.100 66.885 53.380 67.675 ;
    END
  END BIT_SEL[15]
  OBS
      LAYER Metal1 ;
        RECT 25.090 363.855 25.690 382.710 ;
        RECT 29.010 363.855 29.610 382.710 ;
        RECT 31.650 381.475 62.170 381.855 ;
        RECT 64.100 381.475 94.620 381.855 ;
        RECT 96.550 381.475 127.070 381.855 ;
        RECT 129.000 381.475 159.520 381.855 ;
        RECT 30.800 381.220 31.420 381.405 ;
        RECT 62.400 381.220 63.020 381.405 ;
        RECT 30.800 380.990 63.020 381.220 ;
        RECT 30.800 380.805 31.420 380.990 ;
        RECT 62.400 380.805 63.020 380.990 ;
        RECT 63.250 381.220 63.870 381.405 ;
        RECT 94.850 381.220 95.470 381.405 ;
        RECT 63.250 380.990 95.470 381.220 ;
        RECT 63.250 380.805 63.870 380.990 ;
        RECT 94.850 380.805 95.470 380.990 ;
        RECT 95.700 381.220 96.320 381.405 ;
        RECT 127.300 381.220 127.920 381.405 ;
        RECT 95.700 380.990 127.920 381.220 ;
        RECT 95.700 380.805 96.320 380.990 ;
        RECT 127.300 380.805 127.920 380.990 ;
        RECT 128.150 381.220 128.770 381.405 ;
        RECT 159.750 381.220 160.370 381.405 ;
        RECT 128.150 380.990 160.370 381.220 ;
        RECT 128.150 380.805 128.770 380.990 ;
        RECT 159.750 380.805 160.370 380.990 ;
        RECT 58.400 380.725 60.020 380.735 ;
        RECT 90.850 380.725 92.470 380.735 ;
        RECT 123.300 380.725 124.920 380.735 ;
        RECT 155.750 380.725 157.370 380.735 ;
        RECT 31.650 380.355 62.170 380.725 ;
        RECT 64.100 380.355 94.620 380.725 ;
        RECT 96.550 380.355 127.070 380.725 ;
        RECT 129.000 380.355 159.520 380.725 ;
        RECT 31.650 379.635 62.170 380.015 ;
        RECT 64.100 379.635 94.620 380.015 ;
        RECT 96.550 379.635 127.070 380.015 ;
        RECT 129.000 379.635 159.520 380.015 ;
        RECT 30.800 379.380 31.420 379.565 ;
        RECT 62.400 379.380 63.020 379.565 ;
        RECT 30.800 379.150 63.020 379.380 ;
        RECT 30.800 378.965 31.420 379.150 ;
        RECT 62.400 378.965 63.020 379.150 ;
        RECT 63.250 379.380 63.870 379.565 ;
        RECT 94.850 379.380 95.470 379.565 ;
        RECT 63.250 379.150 95.470 379.380 ;
        RECT 63.250 378.965 63.870 379.150 ;
        RECT 94.850 378.965 95.470 379.150 ;
        RECT 95.700 379.380 96.320 379.565 ;
        RECT 127.300 379.380 127.920 379.565 ;
        RECT 95.700 379.150 127.920 379.380 ;
        RECT 95.700 378.965 96.320 379.150 ;
        RECT 127.300 378.965 127.920 379.150 ;
        RECT 128.150 379.380 128.770 379.565 ;
        RECT 159.750 379.380 160.370 379.565 ;
        RECT 128.150 379.150 160.370 379.380 ;
        RECT 128.150 378.965 128.770 379.150 ;
        RECT 159.750 378.965 160.370 379.150 ;
        RECT 54.560 378.885 56.180 378.895 ;
        RECT 87.010 378.885 88.630 378.895 ;
        RECT 119.460 378.885 121.080 378.895 ;
        RECT 151.910 378.885 153.530 378.895 ;
        RECT 31.650 378.515 62.170 378.885 ;
        RECT 64.100 378.515 94.620 378.885 ;
        RECT 96.550 378.515 127.070 378.885 ;
        RECT 129.000 378.515 159.520 378.885 ;
        RECT 31.660 377.720 62.160 378.160 ;
        RECT 64.110 377.720 94.610 378.160 ;
        RECT 96.560 377.720 127.060 378.160 ;
        RECT 129.010 377.720 159.510 378.160 ;
        RECT 31.650 376.990 62.170 377.370 ;
        RECT 64.100 376.990 94.620 377.370 ;
        RECT 96.550 376.990 127.070 377.370 ;
        RECT 129.000 376.990 159.520 377.370 ;
        RECT 30.800 376.735 31.420 376.920 ;
        RECT 62.400 376.735 63.020 376.920 ;
        RECT 30.800 376.505 63.020 376.735 ;
        RECT 30.800 376.320 31.420 376.505 ;
        RECT 62.400 376.320 63.020 376.505 ;
        RECT 63.250 376.735 63.870 376.920 ;
        RECT 94.850 376.735 95.470 376.920 ;
        RECT 63.250 376.505 95.470 376.735 ;
        RECT 63.250 376.320 63.870 376.505 ;
        RECT 94.850 376.320 95.470 376.505 ;
        RECT 95.700 376.735 96.320 376.920 ;
        RECT 127.300 376.735 127.920 376.920 ;
        RECT 95.700 376.505 127.920 376.735 ;
        RECT 95.700 376.320 96.320 376.505 ;
        RECT 127.300 376.320 127.920 376.505 ;
        RECT 128.150 376.735 128.770 376.920 ;
        RECT 159.750 376.735 160.370 376.920 ;
        RECT 128.150 376.505 160.370 376.735 ;
        RECT 128.150 376.320 128.770 376.505 ;
        RECT 159.750 376.320 160.370 376.505 ;
        RECT 50.720 376.240 52.340 376.250 ;
        RECT 83.170 376.240 84.790 376.250 ;
        RECT 115.620 376.240 117.240 376.250 ;
        RECT 148.070 376.240 149.690 376.250 ;
        RECT 31.650 375.870 62.170 376.240 ;
        RECT 64.100 375.870 94.620 376.240 ;
        RECT 96.550 375.870 127.070 376.240 ;
        RECT 129.000 375.870 159.520 376.240 ;
        RECT 31.650 375.150 62.170 375.530 ;
        RECT 64.100 375.150 94.620 375.530 ;
        RECT 96.550 375.150 127.070 375.530 ;
        RECT 129.000 375.150 159.520 375.530 ;
        RECT 30.800 374.895 31.420 375.080 ;
        RECT 62.400 374.895 63.020 375.080 ;
        RECT 30.800 374.665 63.020 374.895 ;
        RECT 30.800 374.480 31.420 374.665 ;
        RECT 62.400 374.480 63.020 374.665 ;
        RECT 63.250 374.895 63.870 375.080 ;
        RECT 94.850 374.895 95.470 375.080 ;
        RECT 63.250 374.665 95.470 374.895 ;
        RECT 63.250 374.480 63.870 374.665 ;
        RECT 94.850 374.480 95.470 374.665 ;
        RECT 95.700 374.895 96.320 375.080 ;
        RECT 127.300 374.895 127.920 375.080 ;
        RECT 95.700 374.665 127.920 374.895 ;
        RECT 95.700 374.480 96.320 374.665 ;
        RECT 127.300 374.480 127.920 374.665 ;
        RECT 128.150 374.895 128.770 375.080 ;
        RECT 159.750 374.895 160.370 375.080 ;
        RECT 128.150 374.665 160.370 374.895 ;
        RECT 128.150 374.480 128.770 374.665 ;
        RECT 159.750 374.480 160.370 374.665 ;
        RECT 46.880 374.400 48.500 374.410 ;
        RECT 79.330 374.400 80.950 374.410 ;
        RECT 111.780 374.400 113.400 374.410 ;
        RECT 144.230 374.400 145.850 374.410 ;
        RECT 31.650 374.030 62.170 374.400 ;
        RECT 64.100 374.030 94.620 374.400 ;
        RECT 96.550 374.030 127.070 374.400 ;
        RECT 129.000 374.030 159.520 374.400 ;
        RECT 31.650 373.310 62.170 373.690 ;
        RECT 64.100 373.310 94.620 373.690 ;
        RECT 96.550 373.310 127.070 373.690 ;
        RECT 129.000 373.310 159.520 373.690 ;
        RECT 30.800 373.055 31.420 373.240 ;
        RECT 62.400 373.055 63.020 373.240 ;
        RECT 30.800 372.825 63.020 373.055 ;
        RECT 30.800 372.640 31.420 372.825 ;
        RECT 62.400 372.640 63.020 372.825 ;
        RECT 63.250 373.055 63.870 373.240 ;
        RECT 94.850 373.055 95.470 373.240 ;
        RECT 63.250 372.825 95.470 373.055 ;
        RECT 63.250 372.640 63.870 372.825 ;
        RECT 94.850 372.640 95.470 372.825 ;
        RECT 95.700 373.055 96.320 373.240 ;
        RECT 127.300 373.055 127.920 373.240 ;
        RECT 95.700 372.825 127.920 373.055 ;
        RECT 95.700 372.640 96.320 372.825 ;
        RECT 127.300 372.640 127.920 372.825 ;
        RECT 128.150 373.055 128.770 373.240 ;
        RECT 159.750 373.055 160.370 373.240 ;
        RECT 128.150 372.825 160.370 373.055 ;
        RECT 128.150 372.640 128.770 372.825 ;
        RECT 159.750 372.640 160.370 372.825 ;
        RECT 43.040 372.560 44.660 372.570 ;
        RECT 75.490 372.560 77.110 372.570 ;
        RECT 107.940 372.560 109.560 372.570 ;
        RECT 140.390 372.560 142.010 372.570 ;
        RECT 31.650 372.190 62.170 372.560 ;
        RECT 64.100 372.190 94.620 372.560 ;
        RECT 96.550 372.190 127.070 372.560 ;
        RECT 129.000 372.190 159.520 372.560 ;
        RECT 31.660 371.395 62.160 371.835 ;
        RECT 64.110 371.395 94.610 371.835 ;
        RECT 96.560 371.395 127.060 371.835 ;
        RECT 129.010 371.395 159.510 371.835 ;
        RECT 31.650 370.665 62.170 371.045 ;
        RECT 64.100 370.665 94.620 371.045 ;
        RECT 96.550 370.665 127.070 371.045 ;
        RECT 129.000 370.665 159.520 371.045 ;
        RECT 30.800 370.410 31.420 370.595 ;
        RECT 62.400 370.410 63.020 370.595 ;
        RECT 30.800 370.180 63.020 370.410 ;
        RECT 30.800 369.995 31.420 370.180 ;
        RECT 62.400 369.995 63.020 370.180 ;
        RECT 63.250 370.410 63.870 370.595 ;
        RECT 94.850 370.410 95.470 370.595 ;
        RECT 63.250 370.180 95.470 370.410 ;
        RECT 63.250 369.995 63.870 370.180 ;
        RECT 94.850 369.995 95.470 370.180 ;
        RECT 95.700 370.410 96.320 370.595 ;
        RECT 127.300 370.410 127.920 370.595 ;
        RECT 95.700 370.180 127.920 370.410 ;
        RECT 95.700 369.995 96.320 370.180 ;
        RECT 127.300 369.995 127.920 370.180 ;
        RECT 128.150 370.410 128.770 370.595 ;
        RECT 159.750 370.410 160.370 370.595 ;
        RECT 128.150 370.180 160.370 370.410 ;
        RECT 128.150 369.995 128.770 370.180 ;
        RECT 159.750 369.995 160.370 370.180 ;
        RECT 39.200 369.915 40.820 369.925 ;
        RECT 71.650 369.915 73.270 369.925 ;
        RECT 104.100 369.915 105.720 369.925 ;
        RECT 136.550 369.915 138.170 369.925 ;
        RECT 31.650 369.545 62.170 369.915 ;
        RECT 64.100 369.545 94.620 369.915 ;
        RECT 96.550 369.545 127.070 369.915 ;
        RECT 129.000 369.545 159.520 369.915 ;
        RECT 31.650 368.825 62.170 369.205 ;
        RECT 64.100 368.825 94.620 369.205 ;
        RECT 96.550 368.825 127.070 369.205 ;
        RECT 129.000 368.825 159.520 369.205 ;
        RECT 30.800 368.570 31.420 368.755 ;
        RECT 62.400 368.570 63.020 368.755 ;
        RECT 30.800 368.340 63.020 368.570 ;
        RECT 30.800 368.155 31.420 368.340 ;
        RECT 62.400 368.155 63.020 368.340 ;
        RECT 63.250 368.570 63.870 368.755 ;
        RECT 94.850 368.570 95.470 368.755 ;
        RECT 63.250 368.340 95.470 368.570 ;
        RECT 63.250 368.155 63.870 368.340 ;
        RECT 94.850 368.155 95.470 368.340 ;
        RECT 95.700 368.570 96.320 368.755 ;
        RECT 127.300 368.570 127.920 368.755 ;
        RECT 95.700 368.340 127.920 368.570 ;
        RECT 95.700 368.155 96.320 368.340 ;
        RECT 127.300 368.155 127.920 368.340 ;
        RECT 128.150 368.570 128.770 368.755 ;
        RECT 159.750 368.570 160.370 368.755 ;
        RECT 128.150 368.340 160.370 368.570 ;
        RECT 128.150 368.155 128.770 368.340 ;
        RECT 159.750 368.155 160.370 368.340 ;
        RECT 35.360 368.075 36.980 368.085 ;
        RECT 67.810 368.075 69.430 368.085 ;
        RECT 100.260 368.075 101.880 368.085 ;
        RECT 132.710 368.075 134.330 368.085 ;
        RECT 31.650 367.705 62.170 368.075 ;
        RECT 64.100 367.705 94.620 368.075 ;
        RECT 96.550 367.705 127.070 368.075 ;
        RECT 129.000 367.705 159.520 368.075 ;
        RECT 31.650 366.985 62.170 367.365 ;
        RECT 64.100 366.985 94.620 367.365 ;
        RECT 96.550 366.985 127.070 367.365 ;
        RECT 129.000 366.985 159.520 367.365 ;
        RECT 30.800 366.730 31.420 366.915 ;
        RECT 62.400 366.730 63.020 366.915 ;
        RECT 30.800 366.500 63.020 366.730 ;
        RECT 30.800 366.315 31.420 366.500 ;
        RECT 62.400 366.315 63.020 366.500 ;
        RECT 63.250 366.730 63.870 366.915 ;
        RECT 94.850 366.730 95.470 366.915 ;
        RECT 63.250 366.500 95.470 366.730 ;
        RECT 63.250 366.315 63.870 366.500 ;
        RECT 94.850 366.315 95.470 366.500 ;
        RECT 95.700 366.730 96.320 366.915 ;
        RECT 127.300 366.730 127.920 366.915 ;
        RECT 95.700 366.500 127.920 366.730 ;
        RECT 95.700 366.315 96.320 366.500 ;
        RECT 127.300 366.315 127.920 366.500 ;
        RECT 128.150 366.730 128.770 366.915 ;
        RECT 159.750 366.730 160.370 366.915 ;
        RECT 128.150 366.500 160.370 366.730 ;
        RECT 128.150 366.315 128.770 366.500 ;
        RECT 159.750 366.315 160.370 366.500 ;
        RECT 31.650 365.865 62.170 366.235 ;
        RECT 64.100 365.865 94.620 366.235 ;
        RECT 96.550 365.865 127.070 366.235 ;
        RECT 129.000 365.865 159.520 366.235 ;
        RECT 25.090 363.515 27.380 363.855 ;
        RECT 28.125 363.515 29.610 363.855 ;
        RECT 25.090 362.880 25.690 363.515 ;
        RECT 25.090 362.650 26.670 362.880 ;
        RECT 25.090 360.610 25.690 362.650 ;
        RECT 27.100 362.420 27.460 362.505 ;
        RECT 25.970 362.190 27.460 362.420 ;
        RECT 25.970 362.040 26.330 362.190 ;
        RECT 25.920 361.405 26.870 361.810 ;
        RECT 25.090 360.380 26.380 360.610 ;
        RECT 25.090 359.420 25.690 360.380 ;
        RECT 26.610 360.060 26.870 361.405 ;
        RECT 27.100 360.755 27.460 362.190 ;
        RECT 27.690 360.855 28.040 362.055 ;
        RECT 28.400 361.445 28.780 363.090 ;
        RECT 27.480 360.060 27.830 360.120 ;
        RECT 28.400 360.060 28.740 360.665 ;
        RECT 26.610 359.800 28.740 360.060 ;
        RECT 27.480 359.740 27.830 359.800 ;
        RECT 29.010 359.520 29.610 363.515 ;
        RECT 31.455 363.080 33.205 365.865 ;
        RECT 33.845 363.080 34.655 364.080 ;
        RECT 35.295 363.080 37.045 365.375 ;
        RECT 37.685 363.080 38.495 364.080 ;
        RECT 39.135 363.080 40.885 365.375 ;
        RECT 41.525 363.080 42.335 364.080 ;
        RECT 42.975 363.080 44.725 365.375 ;
        RECT 45.365 363.080 46.175 364.080 ;
        RECT 46.815 363.080 48.565 365.375 ;
        RECT 49.205 363.080 50.015 364.080 ;
        RECT 50.655 363.080 52.405 365.375 ;
        RECT 53.045 363.080 53.855 364.080 ;
        RECT 54.495 363.080 56.245 365.375 ;
        RECT 56.885 363.080 57.695 364.080 ;
        RECT 58.335 363.080 60.085 365.375 ;
        RECT 60.725 363.080 61.535 364.080 ;
        RECT 63.905 363.080 65.655 365.865 ;
        RECT 66.295 363.080 67.105 364.080 ;
        RECT 67.745 363.080 69.495 365.375 ;
        RECT 70.135 363.080 70.945 364.080 ;
        RECT 71.585 363.080 73.335 365.375 ;
        RECT 73.975 363.080 74.785 364.080 ;
        RECT 75.425 363.080 77.175 365.375 ;
        RECT 77.815 363.080 78.625 364.080 ;
        RECT 79.265 363.080 81.015 365.375 ;
        RECT 81.655 363.080 82.465 364.080 ;
        RECT 83.105 363.080 84.855 365.375 ;
        RECT 85.495 363.080 86.305 364.080 ;
        RECT 86.945 363.080 88.695 365.375 ;
        RECT 89.335 363.080 90.145 364.080 ;
        RECT 90.785 363.080 92.535 365.375 ;
        RECT 93.175 363.080 93.985 364.080 ;
        RECT 96.355 363.080 98.105 365.865 ;
        RECT 98.745 363.080 99.555 364.080 ;
        RECT 100.195 363.080 101.945 365.375 ;
        RECT 102.585 363.080 103.395 364.080 ;
        RECT 104.035 363.080 105.785 365.375 ;
        RECT 106.425 363.080 107.235 364.080 ;
        RECT 107.875 363.080 109.625 365.375 ;
        RECT 110.265 363.080 111.075 364.080 ;
        RECT 111.715 363.080 113.465 365.375 ;
        RECT 114.105 363.080 114.915 364.080 ;
        RECT 115.555 363.080 117.305 365.375 ;
        RECT 117.945 363.080 118.755 364.080 ;
        RECT 119.395 363.080 121.145 365.375 ;
        RECT 121.785 363.080 122.595 364.080 ;
        RECT 123.235 363.080 124.985 365.375 ;
        RECT 125.625 363.080 126.435 364.080 ;
        RECT 128.805 363.080 130.555 365.865 ;
        RECT 131.195 363.080 132.005 364.080 ;
        RECT 132.645 363.080 134.395 365.375 ;
        RECT 135.035 363.080 135.845 364.080 ;
        RECT 136.485 363.080 138.235 365.375 ;
        RECT 138.875 363.080 139.685 364.080 ;
        RECT 140.325 363.080 142.075 365.375 ;
        RECT 142.715 363.080 143.525 364.080 ;
        RECT 144.165 363.080 145.915 365.375 ;
        RECT 146.555 363.080 147.365 364.080 ;
        RECT 148.005 363.080 149.755 365.375 ;
        RECT 150.395 363.080 151.205 364.080 ;
        RECT 151.845 363.080 153.595 365.375 ;
        RECT 154.235 363.080 155.045 364.080 ;
        RECT 155.685 363.080 157.435 365.375 ;
        RECT 158.075 363.080 158.885 364.080 ;
        RECT 161.300 363.270 161.670 381.780 ;
        RECT 162.320 378.145 162.690 381.780 ;
        RECT 162.315 377.765 162.695 378.145 ;
        RECT 162.320 375.145 162.690 377.765 ;
        RECT 162.315 374.765 162.695 375.145 ;
        RECT 162.320 372.145 162.690 374.765 ;
        RECT 162.315 371.765 162.695 372.145 ;
        RECT 162.320 369.145 162.690 371.765 ;
        RECT 162.315 368.765 162.695 369.145 ;
        RECT 162.320 366.145 162.690 368.765 ;
        RECT 162.315 365.765 162.695 366.145 ;
        RECT 161.300 362.890 161.680 363.270 ;
        RECT 161.300 361.820 161.670 362.890 ;
        RECT 31.925 360.630 32.735 361.630 ;
        RECT 25.090 359.190 26.780 359.420 ;
        RECT 28.150 359.290 29.610 359.520 ;
        RECT 25.090 357.180 25.690 359.190 ;
        RECT 27.110 358.730 28.110 359.055 ;
        RECT 25.920 358.170 28.780 358.500 ;
        RECT 25.090 356.950 26.780 357.180 ;
        RECT 25.090 354.940 25.690 356.950 ;
        RECT 27.495 356.815 27.760 358.170 ;
        RECT 29.010 357.280 29.610 359.290 ;
        RECT 33.375 358.800 35.125 361.630 ;
        RECT 35.765 360.630 36.575 361.630 ;
        RECT 37.215 359.335 38.965 361.630 ;
        RECT 39.605 360.630 40.415 361.630 ;
        RECT 41.055 359.335 42.805 361.630 ;
        RECT 43.445 360.630 44.255 361.630 ;
        RECT 44.895 359.335 46.645 361.630 ;
        RECT 47.285 360.630 48.095 361.630 ;
        RECT 48.735 359.335 50.485 361.630 ;
        RECT 51.125 360.630 51.935 361.630 ;
        RECT 52.575 359.335 54.325 361.630 ;
        RECT 54.965 360.630 55.775 361.630 ;
        RECT 56.415 359.335 58.165 361.630 ;
        RECT 58.805 360.630 59.615 361.630 ;
        RECT 60.255 359.335 62.005 361.630 ;
        RECT 64.375 360.630 65.185 361.630 ;
        RECT 65.825 358.800 67.575 361.630 ;
        RECT 68.215 360.630 69.025 361.630 ;
        RECT 69.665 359.335 71.415 361.630 ;
        RECT 72.055 360.630 72.865 361.630 ;
        RECT 73.505 359.335 75.255 361.630 ;
        RECT 75.895 360.630 76.705 361.630 ;
        RECT 77.345 359.335 79.095 361.630 ;
        RECT 79.735 360.630 80.545 361.630 ;
        RECT 81.185 359.335 82.935 361.630 ;
        RECT 83.575 360.630 84.385 361.630 ;
        RECT 85.025 359.335 86.775 361.630 ;
        RECT 87.415 360.630 88.225 361.630 ;
        RECT 88.865 359.335 90.615 361.630 ;
        RECT 91.255 360.630 92.065 361.630 ;
        RECT 92.705 359.335 94.455 361.630 ;
        RECT 96.825 360.630 97.635 361.630 ;
        RECT 98.275 358.800 100.025 361.630 ;
        RECT 100.665 360.630 101.475 361.630 ;
        RECT 102.115 359.335 103.865 361.630 ;
        RECT 104.505 360.630 105.315 361.630 ;
        RECT 105.955 359.335 107.705 361.630 ;
        RECT 108.345 360.630 109.155 361.630 ;
        RECT 109.795 359.335 111.545 361.630 ;
        RECT 112.185 360.630 112.995 361.630 ;
        RECT 113.635 359.335 115.385 361.630 ;
        RECT 116.025 360.630 116.835 361.630 ;
        RECT 117.475 359.335 119.225 361.630 ;
        RECT 119.865 360.630 120.675 361.630 ;
        RECT 121.315 359.335 123.065 361.630 ;
        RECT 123.705 360.630 124.515 361.630 ;
        RECT 125.155 359.335 126.905 361.630 ;
        RECT 129.275 360.630 130.085 361.630 ;
        RECT 130.725 358.800 132.475 361.630 ;
        RECT 133.115 360.630 133.925 361.630 ;
        RECT 134.565 359.335 136.315 361.630 ;
        RECT 136.955 360.630 137.765 361.630 ;
        RECT 138.405 359.335 140.155 361.630 ;
        RECT 140.795 360.630 141.605 361.630 ;
        RECT 142.245 359.335 143.995 361.630 ;
        RECT 144.635 360.630 145.445 361.630 ;
        RECT 146.085 359.335 147.835 361.630 ;
        RECT 148.475 360.630 149.285 361.630 ;
        RECT 149.925 359.335 151.675 361.630 ;
        RECT 152.315 360.630 153.125 361.630 ;
        RECT 153.765 359.335 155.515 361.630 ;
        RECT 156.155 360.630 156.965 361.630 ;
        RECT 157.605 359.335 159.355 361.630 ;
        RECT 161.300 361.440 161.680 361.820 ;
        RECT 31.650 358.430 62.170 358.800 ;
        RECT 64.100 358.430 94.620 358.800 ;
        RECT 96.550 358.430 127.070 358.800 ;
        RECT 129.000 358.430 159.520 358.800 ;
        RECT 30.800 358.165 31.420 358.350 ;
        RECT 62.400 358.165 63.020 358.350 ;
        RECT 30.800 357.935 63.020 358.165 ;
        RECT 30.800 357.750 31.420 357.935 ;
        RECT 62.400 357.750 63.020 357.935 ;
        RECT 63.250 358.165 63.870 358.350 ;
        RECT 94.850 358.165 95.470 358.350 ;
        RECT 63.250 357.935 95.470 358.165 ;
        RECT 63.250 357.750 63.870 357.935 ;
        RECT 94.850 357.750 95.470 357.935 ;
        RECT 95.700 358.165 96.320 358.350 ;
        RECT 127.300 358.165 127.920 358.350 ;
        RECT 95.700 357.935 127.920 358.165 ;
        RECT 95.700 357.750 96.320 357.935 ;
        RECT 127.300 357.750 127.920 357.935 ;
        RECT 128.150 358.165 128.770 358.350 ;
        RECT 159.750 358.165 160.370 358.350 ;
        RECT 128.150 357.935 160.370 358.165 ;
        RECT 128.150 357.750 128.770 357.935 ;
        RECT 159.750 357.750 160.370 357.935 ;
        RECT 31.650 357.300 62.170 357.680 ;
        RECT 64.100 357.300 94.620 357.680 ;
        RECT 96.550 357.300 127.070 357.680 ;
        RECT 129.000 357.300 159.520 357.680 ;
        RECT 28.150 357.050 29.610 357.280 ;
        RECT 27.110 356.490 28.110 356.815 ;
        RECT 25.920 355.930 28.780 356.260 ;
        RECT 29.010 355.040 29.610 357.050 ;
        RECT 31.650 356.590 62.170 356.960 ;
        RECT 64.100 356.590 94.620 356.960 ;
        RECT 96.550 356.590 127.070 356.960 ;
        RECT 129.000 356.590 159.520 356.960 ;
        RECT 37.280 356.580 38.900 356.590 ;
        RECT 69.730 356.580 71.350 356.590 ;
        RECT 102.180 356.580 103.800 356.590 ;
        RECT 134.630 356.580 136.250 356.590 ;
        RECT 30.800 356.325 31.420 356.510 ;
        RECT 62.400 356.325 63.020 356.510 ;
        RECT 30.800 356.095 63.020 356.325 ;
        RECT 30.800 355.910 31.420 356.095 ;
        RECT 62.400 355.910 63.020 356.095 ;
        RECT 63.250 356.325 63.870 356.510 ;
        RECT 94.850 356.325 95.470 356.510 ;
        RECT 63.250 356.095 95.470 356.325 ;
        RECT 63.250 355.910 63.870 356.095 ;
        RECT 94.850 355.910 95.470 356.095 ;
        RECT 95.700 356.325 96.320 356.510 ;
        RECT 127.300 356.325 127.920 356.510 ;
        RECT 95.700 356.095 127.920 356.325 ;
        RECT 95.700 355.910 96.320 356.095 ;
        RECT 127.300 355.910 127.920 356.095 ;
        RECT 128.150 356.325 128.770 356.510 ;
        RECT 159.750 356.325 160.370 356.510 ;
        RECT 128.150 356.095 160.370 356.325 ;
        RECT 128.150 355.910 128.770 356.095 ;
        RECT 159.750 355.910 160.370 356.095 ;
        RECT 31.650 355.460 62.170 355.840 ;
        RECT 64.100 355.460 94.620 355.840 ;
        RECT 96.550 355.460 127.070 355.840 ;
        RECT 129.000 355.460 159.520 355.840 ;
        RECT 25.090 354.710 26.780 354.940 ;
        RECT 28.150 354.810 29.610 355.040 ;
        RECT 25.090 352.655 25.690 354.710 ;
        RECT 27.110 354.250 28.110 354.575 ;
        RECT 29.010 352.655 29.610 354.810 ;
        RECT 31.650 354.745 62.170 355.115 ;
        RECT 64.100 354.745 94.620 355.115 ;
        RECT 96.550 354.745 127.070 355.115 ;
        RECT 129.000 354.745 159.520 355.115 ;
        RECT 41.120 354.735 42.740 354.745 ;
        RECT 73.570 354.735 75.190 354.745 ;
        RECT 106.020 354.735 107.640 354.745 ;
        RECT 138.470 354.735 140.090 354.745 ;
        RECT 30.800 354.480 31.420 354.665 ;
        RECT 62.400 354.480 63.020 354.665 ;
        RECT 30.800 354.250 63.020 354.480 ;
        RECT 30.800 354.065 31.420 354.250 ;
        RECT 62.400 354.065 63.020 354.250 ;
        RECT 63.250 354.480 63.870 354.665 ;
        RECT 94.850 354.480 95.470 354.665 ;
        RECT 63.250 354.250 95.470 354.480 ;
        RECT 63.250 354.065 63.870 354.250 ;
        RECT 94.850 354.065 95.470 354.250 ;
        RECT 95.700 354.480 96.320 354.665 ;
        RECT 127.300 354.480 127.920 354.665 ;
        RECT 95.700 354.250 127.920 354.480 ;
        RECT 95.700 354.065 96.320 354.250 ;
        RECT 127.300 354.065 127.920 354.250 ;
        RECT 128.150 354.480 128.770 354.665 ;
        RECT 159.750 354.480 160.370 354.665 ;
        RECT 128.150 354.250 160.370 354.480 ;
        RECT 128.150 354.065 128.770 354.250 ;
        RECT 159.750 354.065 160.370 354.250 ;
        RECT 31.650 353.615 62.170 353.995 ;
        RECT 64.100 353.615 94.620 353.995 ;
        RECT 96.550 353.615 127.070 353.995 ;
        RECT 129.000 353.615 159.520 353.995 ;
        RECT 31.660 352.825 62.160 353.265 ;
        RECT 64.110 352.825 94.610 353.265 ;
        RECT 96.560 352.825 127.060 353.265 ;
        RECT 129.010 352.825 159.510 353.265 ;
        RECT 25.090 352.315 27.380 352.655 ;
        RECT 28.125 352.315 29.610 352.655 ;
        RECT 25.090 324.470 25.690 352.315 ;
        RECT 29.010 324.470 29.610 352.315 ;
        RECT 31.650 352.105 62.170 352.475 ;
        RECT 64.100 352.105 94.620 352.475 ;
        RECT 96.550 352.105 127.070 352.475 ;
        RECT 129.000 352.105 159.520 352.475 ;
        RECT 44.960 352.095 46.580 352.105 ;
        RECT 77.410 352.095 79.030 352.105 ;
        RECT 109.860 352.095 111.480 352.105 ;
        RECT 142.310 352.095 143.930 352.105 ;
        RECT 30.800 351.840 31.420 352.025 ;
        RECT 62.400 351.840 63.020 352.025 ;
        RECT 30.800 351.610 63.020 351.840 ;
        RECT 30.800 351.425 31.420 351.610 ;
        RECT 62.400 351.425 63.020 351.610 ;
        RECT 63.250 351.840 63.870 352.025 ;
        RECT 94.850 351.840 95.470 352.025 ;
        RECT 63.250 351.610 95.470 351.840 ;
        RECT 63.250 351.425 63.870 351.610 ;
        RECT 94.850 351.425 95.470 351.610 ;
        RECT 95.700 351.840 96.320 352.025 ;
        RECT 127.300 351.840 127.920 352.025 ;
        RECT 95.700 351.610 127.920 351.840 ;
        RECT 95.700 351.425 96.320 351.610 ;
        RECT 127.300 351.425 127.920 351.610 ;
        RECT 128.150 351.840 128.770 352.025 ;
        RECT 159.750 351.840 160.370 352.025 ;
        RECT 128.150 351.610 160.370 351.840 ;
        RECT 128.150 351.425 128.770 351.610 ;
        RECT 159.750 351.425 160.370 351.610 ;
        RECT 31.650 350.975 62.170 351.355 ;
        RECT 64.100 350.975 94.620 351.355 ;
        RECT 96.550 350.975 127.070 351.355 ;
        RECT 129.000 350.975 159.520 351.355 ;
        RECT 31.650 350.265 62.170 350.635 ;
        RECT 64.100 350.265 94.620 350.635 ;
        RECT 96.550 350.265 127.070 350.635 ;
        RECT 129.000 350.265 159.520 350.635 ;
        RECT 48.800 350.255 50.420 350.265 ;
        RECT 81.250 350.255 82.870 350.265 ;
        RECT 113.700 350.255 115.320 350.265 ;
        RECT 146.150 350.255 147.770 350.265 ;
        RECT 30.800 350.000 31.420 350.185 ;
        RECT 62.400 350.000 63.020 350.185 ;
        RECT 30.800 349.770 63.020 350.000 ;
        RECT 30.800 349.585 31.420 349.770 ;
        RECT 62.400 349.585 63.020 349.770 ;
        RECT 63.250 350.000 63.870 350.185 ;
        RECT 94.850 350.000 95.470 350.185 ;
        RECT 63.250 349.770 95.470 350.000 ;
        RECT 63.250 349.585 63.870 349.770 ;
        RECT 94.850 349.585 95.470 349.770 ;
        RECT 95.700 350.000 96.320 350.185 ;
        RECT 127.300 350.000 127.920 350.185 ;
        RECT 95.700 349.770 127.920 350.000 ;
        RECT 95.700 349.585 96.320 349.770 ;
        RECT 127.300 349.585 127.920 349.770 ;
        RECT 128.150 350.000 128.770 350.185 ;
        RECT 159.750 350.000 160.370 350.185 ;
        RECT 128.150 349.770 160.370 350.000 ;
        RECT 128.150 349.585 128.770 349.770 ;
        RECT 159.750 349.585 160.370 349.770 ;
        RECT 31.650 349.135 62.170 349.515 ;
        RECT 64.100 349.135 94.620 349.515 ;
        RECT 96.550 349.135 127.070 349.515 ;
        RECT 129.000 349.135 159.520 349.515 ;
        RECT 31.650 348.420 62.170 348.790 ;
        RECT 64.100 348.420 94.620 348.790 ;
        RECT 96.550 348.420 127.070 348.790 ;
        RECT 129.000 348.420 159.520 348.790 ;
        RECT 52.640 348.410 54.260 348.420 ;
        RECT 85.090 348.410 86.710 348.420 ;
        RECT 117.540 348.410 119.160 348.420 ;
        RECT 149.990 348.410 151.610 348.420 ;
        RECT 30.800 348.155 31.420 348.340 ;
        RECT 62.400 348.155 63.020 348.340 ;
        RECT 30.800 347.925 63.020 348.155 ;
        RECT 30.800 347.740 31.420 347.925 ;
        RECT 62.400 347.740 63.020 347.925 ;
        RECT 63.250 348.155 63.870 348.340 ;
        RECT 94.850 348.155 95.470 348.340 ;
        RECT 63.250 347.925 95.470 348.155 ;
        RECT 63.250 347.740 63.870 347.925 ;
        RECT 94.850 347.740 95.470 347.925 ;
        RECT 95.700 348.155 96.320 348.340 ;
        RECT 127.300 348.155 127.920 348.340 ;
        RECT 95.700 347.925 127.920 348.155 ;
        RECT 95.700 347.740 96.320 347.925 ;
        RECT 127.300 347.740 127.920 347.925 ;
        RECT 128.150 348.155 128.770 348.340 ;
        RECT 159.750 348.155 160.370 348.340 ;
        RECT 128.150 347.925 160.370 348.155 ;
        RECT 128.150 347.740 128.770 347.925 ;
        RECT 159.750 347.740 160.370 347.925 ;
        RECT 31.650 347.290 62.170 347.670 ;
        RECT 64.100 347.290 94.620 347.670 ;
        RECT 96.550 347.290 127.070 347.670 ;
        RECT 129.000 347.290 159.520 347.670 ;
        RECT 31.660 346.500 62.160 346.940 ;
        RECT 64.110 346.500 94.610 346.940 ;
        RECT 96.560 346.500 127.060 346.940 ;
        RECT 129.010 346.500 159.510 346.940 ;
        RECT 31.650 345.780 62.170 346.150 ;
        RECT 64.100 345.780 94.620 346.150 ;
        RECT 96.550 345.780 127.070 346.150 ;
        RECT 129.000 345.780 159.520 346.150 ;
        RECT 56.480 345.770 58.100 345.780 ;
        RECT 88.930 345.770 90.550 345.780 ;
        RECT 121.380 345.770 123.000 345.780 ;
        RECT 153.830 345.770 155.450 345.780 ;
        RECT 30.800 345.515 31.420 345.700 ;
        RECT 62.400 345.515 63.020 345.700 ;
        RECT 30.800 345.285 63.020 345.515 ;
        RECT 30.800 345.100 31.420 345.285 ;
        RECT 62.400 345.100 63.020 345.285 ;
        RECT 63.250 345.515 63.870 345.700 ;
        RECT 94.850 345.515 95.470 345.700 ;
        RECT 63.250 345.285 95.470 345.515 ;
        RECT 63.250 345.100 63.870 345.285 ;
        RECT 94.850 345.100 95.470 345.285 ;
        RECT 95.700 345.515 96.320 345.700 ;
        RECT 127.300 345.515 127.920 345.700 ;
        RECT 95.700 345.285 127.920 345.515 ;
        RECT 95.700 345.100 96.320 345.285 ;
        RECT 127.300 345.100 127.920 345.285 ;
        RECT 128.150 345.515 128.770 345.700 ;
        RECT 159.750 345.515 160.370 345.700 ;
        RECT 128.150 345.285 160.370 345.515 ;
        RECT 128.150 345.100 128.770 345.285 ;
        RECT 159.750 345.100 160.370 345.285 ;
        RECT 31.650 344.650 62.170 345.030 ;
        RECT 64.100 344.650 94.620 345.030 ;
        RECT 96.550 344.650 127.070 345.030 ;
        RECT 129.000 344.650 159.520 345.030 ;
        RECT 31.650 343.940 62.170 344.310 ;
        RECT 64.100 343.940 94.620 344.310 ;
        RECT 96.550 343.940 127.070 344.310 ;
        RECT 129.000 343.940 159.520 344.310 ;
        RECT 60.320 343.930 61.940 343.940 ;
        RECT 92.770 343.930 94.390 343.940 ;
        RECT 125.220 343.930 126.840 343.940 ;
        RECT 157.670 343.930 159.290 343.940 ;
        RECT 30.800 343.675 31.420 343.860 ;
        RECT 62.400 343.675 63.020 343.860 ;
        RECT 30.800 343.445 63.020 343.675 ;
        RECT 30.800 343.260 31.420 343.445 ;
        RECT 62.400 343.260 63.020 343.445 ;
        RECT 63.250 343.675 63.870 343.860 ;
        RECT 94.850 343.675 95.470 343.860 ;
        RECT 63.250 343.445 95.470 343.675 ;
        RECT 63.250 343.260 63.870 343.445 ;
        RECT 94.850 343.260 95.470 343.445 ;
        RECT 95.700 343.675 96.320 343.860 ;
        RECT 127.300 343.675 127.920 343.860 ;
        RECT 95.700 343.445 127.920 343.675 ;
        RECT 95.700 343.260 96.320 343.445 ;
        RECT 127.300 343.260 127.920 343.445 ;
        RECT 128.150 343.675 128.770 343.860 ;
        RECT 159.750 343.675 160.370 343.860 ;
        RECT 128.150 343.445 160.370 343.675 ;
        RECT 161.300 343.510 161.670 361.440 ;
        RECT 162.320 360.145 162.690 365.765 ;
        RECT 163.340 363.270 163.710 381.780 ;
        RECT 164.360 378.145 164.730 381.780 ;
        RECT 164.355 377.765 164.735 378.145 ;
        RECT 164.360 375.145 164.730 377.765 ;
        RECT 164.355 374.765 164.735 375.145 ;
        RECT 164.360 372.145 164.730 374.765 ;
        RECT 164.355 371.765 164.735 372.145 ;
        RECT 164.360 369.145 164.730 371.765 ;
        RECT 164.355 368.765 164.735 369.145 ;
        RECT 164.360 366.145 164.730 368.765 ;
        RECT 164.355 365.765 164.735 366.145 ;
        RECT 163.340 362.890 163.720 363.270 ;
        RECT 163.340 361.820 163.710 362.890 ;
        RECT 163.340 361.440 163.720 361.820 ;
        RECT 162.315 359.765 162.695 360.145 ;
        RECT 162.320 357.145 162.690 359.765 ;
        RECT 162.315 356.765 162.695 357.145 ;
        RECT 162.320 354.145 162.690 356.765 ;
        RECT 162.315 353.765 162.695 354.145 ;
        RECT 162.320 351.145 162.690 353.765 ;
        RECT 162.315 350.765 162.695 351.145 ;
        RECT 162.320 348.145 162.690 350.765 ;
        RECT 162.315 347.765 162.695 348.145 ;
        RECT 162.320 345.145 162.690 347.765 ;
        RECT 162.315 344.765 162.695 345.145 ;
        RECT 162.320 343.510 162.690 344.765 ;
        RECT 163.340 343.510 163.710 361.440 ;
        RECT 164.360 360.145 164.730 365.765 ;
        RECT 164.355 359.765 164.735 360.145 ;
        RECT 164.360 357.145 164.730 359.765 ;
        RECT 164.355 356.765 164.735 357.145 ;
        RECT 164.360 354.145 164.730 356.765 ;
        RECT 164.355 353.765 164.735 354.145 ;
        RECT 164.360 351.145 164.730 353.765 ;
        RECT 164.355 350.765 164.735 351.145 ;
        RECT 164.360 348.145 164.730 350.765 ;
        RECT 164.355 347.765 164.735 348.145 ;
        RECT 164.360 345.145 164.730 347.765 ;
        RECT 164.355 344.765 164.735 345.145 ;
        RECT 164.360 343.510 164.730 344.765 ;
        RECT 165.380 343.510 165.760 381.780 ;
        RECT 166.110 343.520 166.550 381.770 ;
        RECT 128.150 343.260 128.770 343.445 ;
        RECT 159.750 343.260 160.370 343.445 ;
        RECT 31.650 342.810 62.170 343.190 ;
        RECT 64.100 342.810 94.620 343.190 ;
        RECT 96.550 342.810 127.070 343.190 ;
        RECT 129.000 342.810 159.520 343.190 ;
        RECT 31.650 342.090 62.170 342.470 ;
        RECT 64.100 342.090 94.620 342.470 ;
        RECT 96.550 342.090 127.070 342.470 ;
        RECT 129.000 342.090 159.520 342.470 ;
        RECT 30.800 341.835 31.420 342.020 ;
        RECT 62.400 341.835 63.020 342.020 ;
        RECT 30.800 341.605 63.020 341.835 ;
        RECT 30.800 341.420 31.420 341.605 ;
        RECT 62.400 341.420 63.020 341.605 ;
        RECT 63.250 341.835 63.870 342.020 ;
        RECT 94.850 341.835 95.470 342.020 ;
        RECT 63.250 341.605 95.470 341.835 ;
        RECT 63.250 341.420 63.870 341.605 ;
        RECT 94.850 341.420 95.470 341.605 ;
        RECT 95.700 341.835 96.320 342.020 ;
        RECT 127.300 341.835 127.920 342.020 ;
        RECT 95.700 341.605 127.920 341.835 ;
        RECT 95.700 341.420 96.320 341.605 ;
        RECT 127.300 341.420 127.920 341.605 ;
        RECT 128.150 341.835 128.770 342.020 ;
        RECT 159.750 341.835 160.370 342.020 ;
        RECT 128.150 341.605 160.370 341.835 ;
        RECT 128.150 341.420 128.770 341.605 ;
        RECT 159.750 341.420 160.370 341.605 ;
        RECT 58.400 341.340 60.020 341.350 ;
        RECT 90.850 341.340 92.470 341.350 ;
        RECT 123.300 341.340 124.920 341.350 ;
        RECT 155.750 341.340 157.370 341.350 ;
        RECT 31.650 340.970 62.170 341.340 ;
        RECT 64.100 340.970 94.620 341.340 ;
        RECT 96.550 340.970 127.070 341.340 ;
        RECT 129.000 340.970 159.520 341.340 ;
        RECT 31.650 340.250 62.170 340.630 ;
        RECT 64.100 340.250 94.620 340.630 ;
        RECT 96.550 340.250 127.070 340.630 ;
        RECT 129.000 340.250 159.520 340.630 ;
        RECT 30.800 339.995 31.420 340.180 ;
        RECT 62.400 339.995 63.020 340.180 ;
        RECT 30.800 339.765 63.020 339.995 ;
        RECT 30.800 339.580 31.420 339.765 ;
        RECT 62.400 339.580 63.020 339.765 ;
        RECT 63.250 339.995 63.870 340.180 ;
        RECT 94.850 339.995 95.470 340.180 ;
        RECT 63.250 339.765 95.470 339.995 ;
        RECT 63.250 339.580 63.870 339.765 ;
        RECT 94.850 339.580 95.470 339.765 ;
        RECT 95.700 339.995 96.320 340.180 ;
        RECT 127.300 339.995 127.920 340.180 ;
        RECT 95.700 339.765 127.920 339.995 ;
        RECT 95.700 339.580 96.320 339.765 ;
        RECT 127.300 339.580 127.920 339.765 ;
        RECT 128.150 339.995 128.770 340.180 ;
        RECT 159.750 339.995 160.370 340.180 ;
        RECT 128.150 339.765 160.370 339.995 ;
        RECT 128.150 339.580 128.770 339.765 ;
        RECT 159.750 339.580 160.370 339.765 ;
        RECT 54.560 339.500 56.180 339.510 ;
        RECT 87.010 339.500 88.630 339.510 ;
        RECT 119.460 339.500 121.080 339.510 ;
        RECT 151.910 339.500 153.530 339.510 ;
        RECT 31.650 339.130 62.170 339.500 ;
        RECT 64.100 339.130 94.620 339.500 ;
        RECT 96.550 339.130 127.070 339.500 ;
        RECT 129.000 339.130 159.520 339.500 ;
        RECT 31.660 338.335 62.160 338.775 ;
        RECT 64.110 338.335 94.610 338.775 ;
        RECT 96.560 338.335 127.060 338.775 ;
        RECT 129.010 338.335 159.510 338.775 ;
        RECT 31.650 337.605 62.170 337.985 ;
        RECT 64.100 337.605 94.620 337.985 ;
        RECT 96.550 337.605 127.070 337.985 ;
        RECT 129.000 337.605 159.520 337.985 ;
        RECT 30.800 337.350 31.420 337.535 ;
        RECT 62.400 337.350 63.020 337.535 ;
        RECT 30.800 337.120 63.020 337.350 ;
        RECT 30.800 336.935 31.420 337.120 ;
        RECT 62.400 336.935 63.020 337.120 ;
        RECT 63.250 337.350 63.870 337.535 ;
        RECT 94.850 337.350 95.470 337.535 ;
        RECT 63.250 337.120 95.470 337.350 ;
        RECT 63.250 336.935 63.870 337.120 ;
        RECT 94.850 336.935 95.470 337.120 ;
        RECT 95.700 337.350 96.320 337.535 ;
        RECT 127.300 337.350 127.920 337.535 ;
        RECT 95.700 337.120 127.920 337.350 ;
        RECT 95.700 336.935 96.320 337.120 ;
        RECT 127.300 336.935 127.920 337.120 ;
        RECT 128.150 337.350 128.770 337.535 ;
        RECT 159.750 337.350 160.370 337.535 ;
        RECT 128.150 337.120 160.370 337.350 ;
        RECT 128.150 336.935 128.770 337.120 ;
        RECT 159.750 336.935 160.370 337.120 ;
        RECT 50.720 336.855 52.340 336.865 ;
        RECT 83.170 336.855 84.790 336.865 ;
        RECT 115.620 336.855 117.240 336.865 ;
        RECT 148.070 336.855 149.690 336.865 ;
        RECT 31.650 336.485 62.170 336.855 ;
        RECT 64.100 336.485 94.620 336.855 ;
        RECT 96.550 336.485 127.070 336.855 ;
        RECT 129.000 336.485 159.520 336.855 ;
        RECT 31.650 335.765 62.170 336.145 ;
        RECT 64.100 335.765 94.620 336.145 ;
        RECT 96.550 335.765 127.070 336.145 ;
        RECT 129.000 335.765 159.520 336.145 ;
        RECT 30.800 335.510 31.420 335.695 ;
        RECT 62.400 335.510 63.020 335.695 ;
        RECT 30.800 335.280 63.020 335.510 ;
        RECT 30.800 335.095 31.420 335.280 ;
        RECT 62.400 335.095 63.020 335.280 ;
        RECT 63.250 335.510 63.870 335.695 ;
        RECT 94.850 335.510 95.470 335.695 ;
        RECT 63.250 335.280 95.470 335.510 ;
        RECT 63.250 335.095 63.870 335.280 ;
        RECT 94.850 335.095 95.470 335.280 ;
        RECT 95.700 335.510 96.320 335.695 ;
        RECT 127.300 335.510 127.920 335.695 ;
        RECT 95.700 335.280 127.920 335.510 ;
        RECT 95.700 335.095 96.320 335.280 ;
        RECT 127.300 335.095 127.920 335.280 ;
        RECT 128.150 335.510 128.770 335.695 ;
        RECT 159.750 335.510 160.370 335.695 ;
        RECT 128.150 335.280 160.370 335.510 ;
        RECT 128.150 335.095 128.770 335.280 ;
        RECT 159.750 335.095 160.370 335.280 ;
        RECT 46.880 335.015 48.500 335.025 ;
        RECT 79.330 335.015 80.950 335.025 ;
        RECT 111.780 335.015 113.400 335.025 ;
        RECT 144.230 335.015 145.850 335.025 ;
        RECT 31.650 334.645 62.170 335.015 ;
        RECT 64.100 334.645 94.620 335.015 ;
        RECT 96.550 334.645 127.070 335.015 ;
        RECT 129.000 334.645 159.520 335.015 ;
        RECT 31.650 333.925 62.170 334.305 ;
        RECT 64.100 333.925 94.620 334.305 ;
        RECT 96.550 333.925 127.070 334.305 ;
        RECT 129.000 333.925 159.520 334.305 ;
        RECT 30.800 333.670 31.420 333.855 ;
        RECT 62.400 333.670 63.020 333.855 ;
        RECT 30.800 333.440 63.020 333.670 ;
        RECT 30.800 333.255 31.420 333.440 ;
        RECT 62.400 333.255 63.020 333.440 ;
        RECT 63.250 333.670 63.870 333.855 ;
        RECT 94.850 333.670 95.470 333.855 ;
        RECT 63.250 333.440 95.470 333.670 ;
        RECT 63.250 333.255 63.870 333.440 ;
        RECT 94.850 333.255 95.470 333.440 ;
        RECT 95.700 333.670 96.320 333.855 ;
        RECT 127.300 333.670 127.920 333.855 ;
        RECT 95.700 333.440 127.920 333.670 ;
        RECT 95.700 333.255 96.320 333.440 ;
        RECT 127.300 333.255 127.920 333.440 ;
        RECT 128.150 333.670 128.770 333.855 ;
        RECT 159.750 333.670 160.370 333.855 ;
        RECT 128.150 333.440 160.370 333.670 ;
        RECT 128.150 333.255 128.770 333.440 ;
        RECT 159.750 333.255 160.370 333.440 ;
        RECT 43.040 333.175 44.660 333.185 ;
        RECT 75.490 333.175 77.110 333.185 ;
        RECT 107.940 333.175 109.560 333.185 ;
        RECT 140.390 333.175 142.010 333.185 ;
        RECT 31.650 332.805 62.170 333.175 ;
        RECT 64.100 332.805 94.620 333.175 ;
        RECT 96.550 332.805 127.070 333.175 ;
        RECT 129.000 332.805 159.520 333.175 ;
        RECT 31.660 332.010 62.160 332.450 ;
        RECT 64.110 332.010 94.610 332.450 ;
        RECT 96.560 332.010 127.060 332.450 ;
        RECT 129.010 332.010 159.510 332.450 ;
        RECT 31.650 331.280 62.170 331.660 ;
        RECT 64.100 331.280 94.620 331.660 ;
        RECT 96.550 331.280 127.070 331.660 ;
        RECT 129.000 331.280 159.520 331.660 ;
        RECT 30.800 331.025 31.420 331.210 ;
        RECT 62.400 331.025 63.020 331.210 ;
        RECT 30.800 330.795 63.020 331.025 ;
        RECT 30.800 330.610 31.420 330.795 ;
        RECT 62.400 330.610 63.020 330.795 ;
        RECT 63.250 331.025 63.870 331.210 ;
        RECT 94.850 331.025 95.470 331.210 ;
        RECT 63.250 330.795 95.470 331.025 ;
        RECT 63.250 330.610 63.870 330.795 ;
        RECT 94.850 330.610 95.470 330.795 ;
        RECT 95.700 331.025 96.320 331.210 ;
        RECT 127.300 331.025 127.920 331.210 ;
        RECT 95.700 330.795 127.920 331.025 ;
        RECT 95.700 330.610 96.320 330.795 ;
        RECT 127.300 330.610 127.920 330.795 ;
        RECT 128.150 331.025 128.770 331.210 ;
        RECT 159.750 331.025 160.370 331.210 ;
        RECT 128.150 330.795 160.370 331.025 ;
        RECT 128.150 330.610 128.770 330.795 ;
        RECT 159.750 330.610 160.370 330.795 ;
        RECT 39.200 330.530 40.820 330.540 ;
        RECT 71.650 330.530 73.270 330.540 ;
        RECT 104.100 330.530 105.720 330.540 ;
        RECT 136.550 330.530 138.170 330.540 ;
        RECT 31.650 330.160 62.170 330.530 ;
        RECT 64.100 330.160 94.620 330.530 ;
        RECT 96.550 330.160 127.070 330.530 ;
        RECT 129.000 330.160 159.520 330.530 ;
        RECT 31.650 329.440 62.170 329.820 ;
        RECT 64.100 329.440 94.620 329.820 ;
        RECT 96.550 329.440 127.070 329.820 ;
        RECT 129.000 329.440 159.520 329.820 ;
        RECT 30.800 329.185 31.420 329.370 ;
        RECT 62.400 329.185 63.020 329.370 ;
        RECT 30.800 328.955 63.020 329.185 ;
        RECT 30.800 328.770 31.420 328.955 ;
        RECT 62.400 328.770 63.020 328.955 ;
        RECT 63.250 329.185 63.870 329.370 ;
        RECT 94.850 329.185 95.470 329.370 ;
        RECT 63.250 328.955 95.470 329.185 ;
        RECT 63.250 328.770 63.870 328.955 ;
        RECT 94.850 328.770 95.470 328.955 ;
        RECT 95.700 329.185 96.320 329.370 ;
        RECT 127.300 329.185 127.920 329.370 ;
        RECT 95.700 328.955 127.920 329.185 ;
        RECT 95.700 328.770 96.320 328.955 ;
        RECT 127.300 328.770 127.920 328.955 ;
        RECT 128.150 329.185 128.770 329.370 ;
        RECT 159.750 329.185 160.370 329.370 ;
        RECT 128.150 328.955 160.370 329.185 ;
        RECT 128.150 328.770 128.770 328.955 ;
        RECT 159.750 328.770 160.370 328.955 ;
        RECT 35.360 328.690 36.980 328.700 ;
        RECT 67.810 328.690 69.430 328.700 ;
        RECT 100.260 328.690 101.880 328.700 ;
        RECT 132.710 328.690 134.330 328.700 ;
        RECT 31.650 328.320 62.170 328.690 ;
        RECT 64.100 328.320 94.620 328.690 ;
        RECT 96.550 328.320 127.070 328.690 ;
        RECT 129.000 328.320 159.520 328.690 ;
        RECT 31.650 327.600 62.170 327.980 ;
        RECT 64.100 327.600 94.620 327.980 ;
        RECT 96.550 327.600 127.070 327.980 ;
        RECT 129.000 327.600 159.520 327.980 ;
        RECT 30.800 327.345 31.420 327.530 ;
        RECT 62.400 327.345 63.020 327.530 ;
        RECT 30.800 327.115 63.020 327.345 ;
        RECT 30.800 326.930 31.420 327.115 ;
        RECT 62.400 326.930 63.020 327.115 ;
        RECT 63.250 327.345 63.870 327.530 ;
        RECT 94.850 327.345 95.470 327.530 ;
        RECT 63.250 327.115 95.470 327.345 ;
        RECT 63.250 326.930 63.870 327.115 ;
        RECT 94.850 326.930 95.470 327.115 ;
        RECT 95.700 327.345 96.320 327.530 ;
        RECT 127.300 327.345 127.920 327.530 ;
        RECT 95.700 327.115 127.920 327.345 ;
        RECT 95.700 326.930 96.320 327.115 ;
        RECT 127.300 326.930 127.920 327.115 ;
        RECT 128.150 327.345 128.770 327.530 ;
        RECT 159.750 327.345 160.370 327.530 ;
        RECT 128.150 327.115 160.370 327.345 ;
        RECT 128.150 326.930 128.770 327.115 ;
        RECT 159.750 326.930 160.370 327.115 ;
        RECT 31.650 326.480 62.170 326.850 ;
        RECT 64.100 326.480 94.620 326.850 ;
        RECT 96.550 326.480 127.070 326.850 ;
        RECT 129.000 326.480 159.520 326.850 ;
        RECT 25.090 324.130 27.380 324.470 ;
        RECT 28.125 324.130 29.610 324.470 ;
        RECT 25.090 323.495 25.690 324.130 ;
        RECT 25.090 323.265 26.670 323.495 ;
        RECT 25.090 321.225 25.690 323.265 ;
        RECT 27.100 323.035 27.460 323.120 ;
        RECT 25.970 322.805 27.460 323.035 ;
        RECT 25.970 322.655 26.330 322.805 ;
        RECT 25.920 322.020 26.870 322.425 ;
        RECT 25.090 320.995 26.380 321.225 ;
        RECT 25.090 320.035 25.690 320.995 ;
        RECT 26.610 320.675 26.870 322.020 ;
        RECT 27.100 321.370 27.460 322.805 ;
        RECT 27.690 321.470 28.040 322.670 ;
        RECT 28.400 322.060 28.780 323.705 ;
        RECT 27.480 320.675 27.830 320.735 ;
        RECT 28.400 320.675 28.740 321.280 ;
        RECT 26.610 320.415 28.740 320.675 ;
        RECT 27.480 320.355 27.830 320.415 ;
        RECT 29.010 320.135 29.610 324.130 ;
        RECT 31.455 323.695 33.205 326.480 ;
        RECT 33.845 323.695 34.655 324.695 ;
        RECT 35.295 323.695 37.045 325.990 ;
        RECT 37.685 323.695 38.495 324.695 ;
        RECT 39.135 323.695 40.885 325.990 ;
        RECT 41.525 323.695 42.335 324.695 ;
        RECT 42.975 323.695 44.725 325.990 ;
        RECT 45.365 323.695 46.175 324.695 ;
        RECT 46.815 323.695 48.565 325.990 ;
        RECT 49.205 323.695 50.015 324.695 ;
        RECT 50.655 323.695 52.405 325.990 ;
        RECT 53.045 323.695 53.855 324.695 ;
        RECT 54.495 323.695 56.245 325.990 ;
        RECT 56.885 323.695 57.695 324.695 ;
        RECT 58.335 323.695 60.085 325.990 ;
        RECT 60.725 323.695 61.535 324.695 ;
        RECT 63.905 323.695 65.655 326.480 ;
        RECT 66.295 323.695 67.105 324.695 ;
        RECT 67.745 323.695 69.495 325.990 ;
        RECT 70.135 323.695 70.945 324.695 ;
        RECT 71.585 323.695 73.335 325.990 ;
        RECT 73.975 323.695 74.785 324.695 ;
        RECT 75.425 323.695 77.175 325.990 ;
        RECT 77.815 323.695 78.625 324.695 ;
        RECT 79.265 323.695 81.015 325.990 ;
        RECT 81.655 323.695 82.465 324.695 ;
        RECT 83.105 323.695 84.855 325.990 ;
        RECT 85.495 323.695 86.305 324.695 ;
        RECT 86.945 323.695 88.695 325.990 ;
        RECT 89.335 323.695 90.145 324.695 ;
        RECT 90.785 323.695 92.535 325.990 ;
        RECT 93.175 323.695 93.985 324.695 ;
        RECT 96.355 323.695 98.105 326.480 ;
        RECT 98.745 323.695 99.555 324.695 ;
        RECT 100.195 323.695 101.945 325.990 ;
        RECT 102.585 323.695 103.395 324.695 ;
        RECT 104.035 323.695 105.785 325.990 ;
        RECT 106.425 323.695 107.235 324.695 ;
        RECT 107.875 323.695 109.625 325.990 ;
        RECT 110.265 323.695 111.075 324.695 ;
        RECT 111.715 323.695 113.465 325.990 ;
        RECT 114.105 323.695 114.915 324.695 ;
        RECT 115.555 323.695 117.305 325.990 ;
        RECT 117.945 323.695 118.755 324.695 ;
        RECT 119.395 323.695 121.145 325.990 ;
        RECT 121.785 323.695 122.595 324.695 ;
        RECT 123.235 323.695 124.985 325.990 ;
        RECT 125.625 323.695 126.435 324.695 ;
        RECT 128.805 323.695 130.555 326.480 ;
        RECT 131.195 323.695 132.005 324.695 ;
        RECT 132.645 323.695 134.395 325.990 ;
        RECT 135.035 323.695 135.845 324.695 ;
        RECT 136.485 323.695 138.235 325.990 ;
        RECT 138.875 323.695 139.685 324.695 ;
        RECT 140.325 323.695 142.075 325.990 ;
        RECT 142.715 323.695 143.525 324.695 ;
        RECT 144.165 323.695 145.915 325.990 ;
        RECT 146.555 323.695 147.365 324.695 ;
        RECT 148.005 323.695 149.755 325.990 ;
        RECT 150.395 323.695 151.205 324.695 ;
        RECT 151.845 323.695 153.595 325.990 ;
        RECT 154.235 323.695 155.045 324.695 ;
        RECT 155.685 323.695 157.435 325.990 ;
        RECT 158.075 323.695 158.885 324.695 ;
        RECT 161.300 323.885 161.670 342.395 ;
        RECT 162.320 338.760 162.690 342.395 ;
        RECT 162.315 338.380 162.695 338.760 ;
        RECT 162.320 335.760 162.690 338.380 ;
        RECT 162.315 335.380 162.695 335.760 ;
        RECT 162.320 332.760 162.690 335.380 ;
        RECT 162.315 332.380 162.695 332.760 ;
        RECT 162.320 329.760 162.690 332.380 ;
        RECT 162.315 329.380 162.695 329.760 ;
        RECT 162.320 326.760 162.690 329.380 ;
        RECT 162.315 326.380 162.695 326.760 ;
        RECT 161.300 323.505 161.680 323.885 ;
        RECT 161.300 322.435 161.670 323.505 ;
        RECT 31.925 321.245 32.735 322.245 ;
        RECT 25.090 319.805 26.780 320.035 ;
        RECT 28.150 319.905 29.610 320.135 ;
        RECT 25.090 317.795 25.690 319.805 ;
        RECT 27.110 319.345 28.110 319.670 ;
        RECT 25.920 318.785 28.780 319.115 ;
        RECT 25.090 317.565 26.780 317.795 ;
        RECT 25.090 315.555 25.690 317.565 ;
        RECT 27.495 317.430 27.760 318.785 ;
        RECT 29.010 317.895 29.610 319.905 ;
        RECT 33.375 319.415 35.125 322.245 ;
        RECT 35.765 321.245 36.575 322.245 ;
        RECT 37.215 319.950 38.965 322.245 ;
        RECT 39.605 321.245 40.415 322.245 ;
        RECT 41.055 319.950 42.805 322.245 ;
        RECT 43.445 321.245 44.255 322.245 ;
        RECT 44.895 319.950 46.645 322.245 ;
        RECT 47.285 321.245 48.095 322.245 ;
        RECT 48.735 319.950 50.485 322.245 ;
        RECT 51.125 321.245 51.935 322.245 ;
        RECT 52.575 319.950 54.325 322.245 ;
        RECT 54.965 321.245 55.775 322.245 ;
        RECT 56.415 319.950 58.165 322.245 ;
        RECT 58.805 321.245 59.615 322.245 ;
        RECT 60.255 319.950 62.005 322.245 ;
        RECT 64.375 321.245 65.185 322.245 ;
        RECT 65.825 319.415 67.575 322.245 ;
        RECT 68.215 321.245 69.025 322.245 ;
        RECT 69.665 319.950 71.415 322.245 ;
        RECT 72.055 321.245 72.865 322.245 ;
        RECT 73.505 319.950 75.255 322.245 ;
        RECT 75.895 321.245 76.705 322.245 ;
        RECT 77.345 319.950 79.095 322.245 ;
        RECT 79.735 321.245 80.545 322.245 ;
        RECT 81.185 319.950 82.935 322.245 ;
        RECT 83.575 321.245 84.385 322.245 ;
        RECT 85.025 319.950 86.775 322.245 ;
        RECT 87.415 321.245 88.225 322.245 ;
        RECT 88.865 319.950 90.615 322.245 ;
        RECT 91.255 321.245 92.065 322.245 ;
        RECT 92.705 319.950 94.455 322.245 ;
        RECT 96.825 321.245 97.635 322.245 ;
        RECT 98.275 319.415 100.025 322.245 ;
        RECT 100.665 321.245 101.475 322.245 ;
        RECT 102.115 319.950 103.865 322.245 ;
        RECT 104.505 321.245 105.315 322.245 ;
        RECT 105.955 319.950 107.705 322.245 ;
        RECT 108.345 321.245 109.155 322.245 ;
        RECT 109.795 319.950 111.545 322.245 ;
        RECT 112.185 321.245 112.995 322.245 ;
        RECT 113.635 319.950 115.385 322.245 ;
        RECT 116.025 321.245 116.835 322.245 ;
        RECT 117.475 319.950 119.225 322.245 ;
        RECT 119.865 321.245 120.675 322.245 ;
        RECT 121.315 319.950 123.065 322.245 ;
        RECT 123.705 321.245 124.515 322.245 ;
        RECT 125.155 319.950 126.905 322.245 ;
        RECT 129.275 321.245 130.085 322.245 ;
        RECT 130.725 319.415 132.475 322.245 ;
        RECT 133.115 321.245 133.925 322.245 ;
        RECT 134.565 319.950 136.315 322.245 ;
        RECT 136.955 321.245 137.765 322.245 ;
        RECT 138.405 319.950 140.155 322.245 ;
        RECT 140.795 321.245 141.605 322.245 ;
        RECT 142.245 319.950 143.995 322.245 ;
        RECT 144.635 321.245 145.445 322.245 ;
        RECT 146.085 319.950 147.835 322.245 ;
        RECT 148.475 321.245 149.285 322.245 ;
        RECT 149.925 319.950 151.675 322.245 ;
        RECT 152.315 321.245 153.125 322.245 ;
        RECT 153.765 319.950 155.515 322.245 ;
        RECT 156.155 321.245 156.965 322.245 ;
        RECT 157.605 319.950 159.355 322.245 ;
        RECT 161.300 322.055 161.680 322.435 ;
        RECT 31.650 319.045 62.170 319.415 ;
        RECT 64.100 319.045 94.620 319.415 ;
        RECT 96.550 319.045 127.070 319.415 ;
        RECT 129.000 319.045 159.520 319.415 ;
        RECT 30.800 318.780 31.420 318.965 ;
        RECT 62.400 318.780 63.020 318.965 ;
        RECT 30.800 318.550 63.020 318.780 ;
        RECT 30.800 318.365 31.420 318.550 ;
        RECT 62.400 318.365 63.020 318.550 ;
        RECT 63.250 318.780 63.870 318.965 ;
        RECT 94.850 318.780 95.470 318.965 ;
        RECT 63.250 318.550 95.470 318.780 ;
        RECT 63.250 318.365 63.870 318.550 ;
        RECT 94.850 318.365 95.470 318.550 ;
        RECT 95.700 318.780 96.320 318.965 ;
        RECT 127.300 318.780 127.920 318.965 ;
        RECT 95.700 318.550 127.920 318.780 ;
        RECT 95.700 318.365 96.320 318.550 ;
        RECT 127.300 318.365 127.920 318.550 ;
        RECT 128.150 318.780 128.770 318.965 ;
        RECT 159.750 318.780 160.370 318.965 ;
        RECT 128.150 318.550 160.370 318.780 ;
        RECT 128.150 318.365 128.770 318.550 ;
        RECT 159.750 318.365 160.370 318.550 ;
        RECT 31.650 317.915 62.170 318.295 ;
        RECT 64.100 317.915 94.620 318.295 ;
        RECT 96.550 317.915 127.070 318.295 ;
        RECT 129.000 317.915 159.520 318.295 ;
        RECT 28.150 317.665 29.610 317.895 ;
        RECT 27.110 317.105 28.110 317.430 ;
        RECT 25.920 316.545 28.780 316.875 ;
        RECT 29.010 315.655 29.610 317.665 ;
        RECT 31.650 317.205 62.170 317.575 ;
        RECT 64.100 317.205 94.620 317.575 ;
        RECT 96.550 317.205 127.070 317.575 ;
        RECT 129.000 317.205 159.520 317.575 ;
        RECT 37.280 317.195 38.900 317.205 ;
        RECT 69.730 317.195 71.350 317.205 ;
        RECT 102.180 317.195 103.800 317.205 ;
        RECT 134.630 317.195 136.250 317.205 ;
        RECT 30.800 316.940 31.420 317.125 ;
        RECT 62.400 316.940 63.020 317.125 ;
        RECT 30.800 316.710 63.020 316.940 ;
        RECT 30.800 316.525 31.420 316.710 ;
        RECT 62.400 316.525 63.020 316.710 ;
        RECT 63.250 316.940 63.870 317.125 ;
        RECT 94.850 316.940 95.470 317.125 ;
        RECT 63.250 316.710 95.470 316.940 ;
        RECT 63.250 316.525 63.870 316.710 ;
        RECT 94.850 316.525 95.470 316.710 ;
        RECT 95.700 316.940 96.320 317.125 ;
        RECT 127.300 316.940 127.920 317.125 ;
        RECT 95.700 316.710 127.920 316.940 ;
        RECT 95.700 316.525 96.320 316.710 ;
        RECT 127.300 316.525 127.920 316.710 ;
        RECT 128.150 316.940 128.770 317.125 ;
        RECT 159.750 316.940 160.370 317.125 ;
        RECT 128.150 316.710 160.370 316.940 ;
        RECT 128.150 316.525 128.770 316.710 ;
        RECT 159.750 316.525 160.370 316.710 ;
        RECT 31.650 316.075 62.170 316.455 ;
        RECT 64.100 316.075 94.620 316.455 ;
        RECT 96.550 316.075 127.070 316.455 ;
        RECT 129.000 316.075 159.520 316.455 ;
        RECT 25.090 315.325 26.780 315.555 ;
        RECT 28.150 315.425 29.610 315.655 ;
        RECT 25.090 313.270 25.690 315.325 ;
        RECT 27.110 314.865 28.110 315.190 ;
        RECT 29.010 313.270 29.610 315.425 ;
        RECT 31.650 315.360 62.170 315.730 ;
        RECT 64.100 315.360 94.620 315.730 ;
        RECT 96.550 315.360 127.070 315.730 ;
        RECT 129.000 315.360 159.520 315.730 ;
        RECT 41.120 315.350 42.740 315.360 ;
        RECT 73.570 315.350 75.190 315.360 ;
        RECT 106.020 315.350 107.640 315.360 ;
        RECT 138.470 315.350 140.090 315.360 ;
        RECT 30.800 315.095 31.420 315.280 ;
        RECT 62.400 315.095 63.020 315.280 ;
        RECT 30.800 314.865 63.020 315.095 ;
        RECT 30.800 314.680 31.420 314.865 ;
        RECT 62.400 314.680 63.020 314.865 ;
        RECT 63.250 315.095 63.870 315.280 ;
        RECT 94.850 315.095 95.470 315.280 ;
        RECT 63.250 314.865 95.470 315.095 ;
        RECT 63.250 314.680 63.870 314.865 ;
        RECT 94.850 314.680 95.470 314.865 ;
        RECT 95.700 315.095 96.320 315.280 ;
        RECT 127.300 315.095 127.920 315.280 ;
        RECT 95.700 314.865 127.920 315.095 ;
        RECT 95.700 314.680 96.320 314.865 ;
        RECT 127.300 314.680 127.920 314.865 ;
        RECT 128.150 315.095 128.770 315.280 ;
        RECT 159.750 315.095 160.370 315.280 ;
        RECT 128.150 314.865 160.370 315.095 ;
        RECT 128.150 314.680 128.770 314.865 ;
        RECT 159.750 314.680 160.370 314.865 ;
        RECT 31.650 314.230 62.170 314.610 ;
        RECT 64.100 314.230 94.620 314.610 ;
        RECT 96.550 314.230 127.070 314.610 ;
        RECT 129.000 314.230 159.520 314.610 ;
        RECT 31.660 313.440 62.160 313.880 ;
        RECT 64.110 313.440 94.610 313.880 ;
        RECT 96.560 313.440 127.060 313.880 ;
        RECT 129.010 313.440 159.510 313.880 ;
        RECT 25.090 312.930 27.380 313.270 ;
        RECT 28.125 312.930 29.610 313.270 ;
        RECT 25.090 285.085 25.690 312.930 ;
        RECT 29.010 285.085 29.610 312.930 ;
        RECT 31.650 312.720 62.170 313.090 ;
        RECT 64.100 312.720 94.620 313.090 ;
        RECT 96.550 312.720 127.070 313.090 ;
        RECT 129.000 312.720 159.520 313.090 ;
        RECT 44.960 312.710 46.580 312.720 ;
        RECT 77.410 312.710 79.030 312.720 ;
        RECT 109.860 312.710 111.480 312.720 ;
        RECT 142.310 312.710 143.930 312.720 ;
        RECT 30.800 312.455 31.420 312.640 ;
        RECT 62.400 312.455 63.020 312.640 ;
        RECT 30.800 312.225 63.020 312.455 ;
        RECT 30.800 312.040 31.420 312.225 ;
        RECT 62.400 312.040 63.020 312.225 ;
        RECT 63.250 312.455 63.870 312.640 ;
        RECT 94.850 312.455 95.470 312.640 ;
        RECT 63.250 312.225 95.470 312.455 ;
        RECT 63.250 312.040 63.870 312.225 ;
        RECT 94.850 312.040 95.470 312.225 ;
        RECT 95.700 312.455 96.320 312.640 ;
        RECT 127.300 312.455 127.920 312.640 ;
        RECT 95.700 312.225 127.920 312.455 ;
        RECT 95.700 312.040 96.320 312.225 ;
        RECT 127.300 312.040 127.920 312.225 ;
        RECT 128.150 312.455 128.770 312.640 ;
        RECT 159.750 312.455 160.370 312.640 ;
        RECT 128.150 312.225 160.370 312.455 ;
        RECT 128.150 312.040 128.770 312.225 ;
        RECT 159.750 312.040 160.370 312.225 ;
        RECT 31.650 311.590 62.170 311.970 ;
        RECT 64.100 311.590 94.620 311.970 ;
        RECT 96.550 311.590 127.070 311.970 ;
        RECT 129.000 311.590 159.520 311.970 ;
        RECT 31.650 310.880 62.170 311.250 ;
        RECT 64.100 310.880 94.620 311.250 ;
        RECT 96.550 310.880 127.070 311.250 ;
        RECT 129.000 310.880 159.520 311.250 ;
        RECT 48.800 310.870 50.420 310.880 ;
        RECT 81.250 310.870 82.870 310.880 ;
        RECT 113.700 310.870 115.320 310.880 ;
        RECT 146.150 310.870 147.770 310.880 ;
        RECT 30.800 310.615 31.420 310.800 ;
        RECT 62.400 310.615 63.020 310.800 ;
        RECT 30.800 310.385 63.020 310.615 ;
        RECT 30.800 310.200 31.420 310.385 ;
        RECT 62.400 310.200 63.020 310.385 ;
        RECT 63.250 310.615 63.870 310.800 ;
        RECT 94.850 310.615 95.470 310.800 ;
        RECT 63.250 310.385 95.470 310.615 ;
        RECT 63.250 310.200 63.870 310.385 ;
        RECT 94.850 310.200 95.470 310.385 ;
        RECT 95.700 310.615 96.320 310.800 ;
        RECT 127.300 310.615 127.920 310.800 ;
        RECT 95.700 310.385 127.920 310.615 ;
        RECT 95.700 310.200 96.320 310.385 ;
        RECT 127.300 310.200 127.920 310.385 ;
        RECT 128.150 310.615 128.770 310.800 ;
        RECT 159.750 310.615 160.370 310.800 ;
        RECT 128.150 310.385 160.370 310.615 ;
        RECT 128.150 310.200 128.770 310.385 ;
        RECT 159.750 310.200 160.370 310.385 ;
        RECT 31.650 309.750 62.170 310.130 ;
        RECT 64.100 309.750 94.620 310.130 ;
        RECT 96.550 309.750 127.070 310.130 ;
        RECT 129.000 309.750 159.520 310.130 ;
        RECT 31.650 309.035 62.170 309.405 ;
        RECT 64.100 309.035 94.620 309.405 ;
        RECT 96.550 309.035 127.070 309.405 ;
        RECT 129.000 309.035 159.520 309.405 ;
        RECT 52.640 309.025 54.260 309.035 ;
        RECT 85.090 309.025 86.710 309.035 ;
        RECT 117.540 309.025 119.160 309.035 ;
        RECT 149.990 309.025 151.610 309.035 ;
        RECT 30.800 308.770 31.420 308.955 ;
        RECT 62.400 308.770 63.020 308.955 ;
        RECT 30.800 308.540 63.020 308.770 ;
        RECT 30.800 308.355 31.420 308.540 ;
        RECT 62.400 308.355 63.020 308.540 ;
        RECT 63.250 308.770 63.870 308.955 ;
        RECT 94.850 308.770 95.470 308.955 ;
        RECT 63.250 308.540 95.470 308.770 ;
        RECT 63.250 308.355 63.870 308.540 ;
        RECT 94.850 308.355 95.470 308.540 ;
        RECT 95.700 308.770 96.320 308.955 ;
        RECT 127.300 308.770 127.920 308.955 ;
        RECT 95.700 308.540 127.920 308.770 ;
        RECT 95.700 308.355 96.320 308.540 ;
        RECT 127.300 308.355 127.920 308.540 ;
        RECT 128.150 308.770 128.770 308.955 ;
        RECT 159.750 308.770 160.370 308.955 ;
        RECT 128.150 308.540 160.370 308.770 ;
        RECT 128.150 308.355 128.770 308.540 ;
        RECT 159.750 308.355 160.370 308.540 ;
        RECT 31.650 307.905 62.170 308.285 ;
        RECT 64.100 307.905 94.620 308.285 ;
        RECT 96.550 307.905 127.070 308.285 ;
        RECT 129.000 307.905 159.520 308.285 ;
        RECT 31.660 307.115 62.160 307.555 ;
        RECT 64.110 307.115 94.610 307.555 ;
        RECT 96.560 307.115 127.060 307.555 ;
        RECT 129.010 307.115 159.510 307.555 ;
        RECT 31.650 306.395 62.170 306.765 ;
        RECT 64.100 306.395 94.620 306.765 ;
        RECT 96.550 306.395 127.070 306.765 ;
        RECT 129.000 306.395 159.520 306.765 ;
        RECT 56.480 306.385 58.100 306.395 ;
        RECT 88.930 306.385 90.550 306.395 ;
        RECT 121.380 306.385 123.000 306.395 ;
        RECT 153.830 306.385 155.450 306.395 ;
        RECT 30.800 306.130 31.420 306.315 ;
        RECT 62.400 306.130 63.020 306.315 ;
        RECT 30.800 305.900 63.020 306.130 ;
        RECT 30.800 305.715 31.420 305.900 ;
        RECT 62.400 305.715 63.020 305.900 ;
        RECT 63.250 306.130 63.870 306.315 ;
        RECT 94.850 306.130 95.470 306.315 ;
        RECT 63.250 305.900 95.470 306.130 ;
        RECT 63.250 305.715 63.870 305.900 ;
        RECT 94.850 305.715 95.470 305.900 ;
        RECT 95.700 306.130 96.320 306.315 ;
        RECT 127.300 306.130 127.920 306.315 ;
        RECT 95.700 305.900 127.920 306.130 ;
        RECT 95.700 305.715 96.320 305.900 ;
        RECT 127.300 305.715 127.920 305.900 ;
        RECT 128.150 306.130 128.770 306.315 ;
        RECT 159.750 306.130 160.370 306.315 ;
        RECT 128.150 305.900 160.370 306.130 ;
        RECT 128.150 305.715 128.770 305.900 ;
        RECT 159.750 305.715 160.370 305.900 ;
        RECT 31.650 305.265 62.170 305.645 ;
        RECT 64.100 305.265 94.620 305.645 ;
        RECT 96.550 305.265 127.070 305.645 ;
        RECT 129.000 305.265 159.520 305.645 ;
        RECT 31.650 304.555 62.170 304.925 ;
        RECT 64.100 304.555 94.620 304.925 ;
        RECT 96.550 304.555 127.070 304.925 ;
        RECT 129.000 304.555 159.520 304.925 ;
        RECT 60.320 304.545 61.940 304.555 ;
        RECT 92.770 304.545 94.390 304.555 ;
        RECT 125.220 304.545 126.840 304.555 ;
        RECT 157.670 304.545 159.290 304.555 ;
        RECT 30.800 304.290 31.420 304.475 ;
        RECT 62.400 304.290 63.020 304.475 ;
        RECT 30.800 304.060 63.020 304.290 ;
        RECT 30.800 303.875 31.420 304.060 ;
        RECT 62.400 303.875 63.020 304.060 ;
        RECT 63.250 304.290 63.870 304.475 ;
        RECT 94.850 304.290 95.470 304.475 ;
        RECT 63.250 304.060 95.470 304.290 ;
        RECT 63.250 303.875 63.870 304.060 ;
        RECT 94.850 303.875 95.470 304.060 ;
        RECT 95.700 304.290 96.320 304.475 ;
        RECT 127.300 304.290 127.920 304.475 ;
        RECT 95.700 304.060 127.920 304.290 ;
        RECT 95.700 303.875 96.320 304.060 ;
        RECT 127.300 303.875 127.920 304.060 ;
        RECT 128.150 304.290 128.770 304.475 ;
        RECT 159.750 304.290 160.370 304.475 ;
        RECT 128.150 304.060 160.370 304.290 ;
        RECT 161.300 304.125 161.670 322.055 ;
        RECT 162.320 320.760 162.690 326.380 ;
        RECT 163.340 323.885 163.710 342.395 ;
        RECT 164.360 338.760 164.730 342.395 ;
        RECT 164.355 338.380 164.735 338.760 ;
        RECT 164.360 335.760 164.730 338.380 ;
        RECT 164.355 335.380 164.735 335.760 ;
        RECT 164.360 332.760 164.730 335.380 ;
        RECT 164.355 332.380 164.735 332.760 ;
        RECT 164.360 329.760 164.730 332.380 ;
        RECT 164.355 329.380 164.735 329.760 ;
        RECT 164.360 326.760 164.730 329.380 ;
        RECT 164.355 326.380 164.735 326.760 ;
        RECT 163.340 323.505 163.720 323.885 ;
        RECT 163.340 322.435 163.710 323.505 ;
        RECT 163.340 322.055 163.720 322.435 ;
        RECT 162.315 320.380 162.695 320.760 ;
        RECT 162.320 317.760 162.690 320.380 ;
        RECT 162.315 317.380 162.695 317.760 ;
        RECT 162.320 314.760 162.690 317.380 ;
        RECT 162.315 314.380 162.695 314.760 ;
        RECT 162.320 311.760 162.690 314.380 ;
        RECT 162.315 311.380 162.695 311.760 ;
        RECT 162.320 308.760 162.690 311.380 ;
        RECT 162.315 308.380 162.695 308.760 ;
        RECT 162.320 305.760 162.690 308.380 ;
        RECT 162.315 305.380 162.695 305.760 ;
        RECT 162.320 304.125 162.690 305.380 ;
        RECT 163.340 304.125 163.710 322.055 ;
        RECT 164.360 320.760 164.730 326.380 ;
        RECT 164.355 320.380 164.735 320.760 ;
        RECT 164.360 317.760 164.730 320.380 ;
        RECT 164.355 317.380 164.735 317.760 ;
        RECT 164.360 314.760 164.730 317.380 ;
        RECT 164.355 314.380 164.735 314.760 ;
        RECT 164.360 311.760 164.730 314.380 ;
        RECT 164.355 311.380 164.735 311.760 ;
        RECT 164.360 308.760 164.730 311.380 ;
        RECT 164.355 308.380 164.735 308.760 ;
        RECT 164.360 305.760 164.730 308.380 ;
        RECT 164.355 305.380 164.735 305.760 ;
        RECT 164.360 304.125 164.730 305.380 ;
        RECT 165.380 304.125 165.760 342.395 ;
        RECT 166.110 304.135 166.550 342.385 ;
        RECT 128.150 303.875 128.770 304.060 ;
        RECT 159.750 303.875 160.370 304.060 ;
        RECT 31.650 303.425 62.170 303.805 ;
        RECT 64.100 303.425 94.620 303.805 ;
        RECT 96.550 303.425 127.070 303.805 ;
        RECT 129.000 303.425 159.520 303.805 ;
        RECT 31.650 302.705 62.170 303.085 ;
        RECT 64.100 302.705 94.620 303.085 ;
        RECT 96.550 302.705 127.070 303.085 ;
        RECT 129.000 302.705 159.520 303.085 ;
        RECT 30.800 302.450 31.420 302.635 ;
        RECT 62.400 302.450 63.020 302.635 ;
        RECT 30.800 302.220 63.020 302.450 ;
        RECT 30.800 302.035 31.420 302.220 ;
        RECT 62.400 302.035 63.020 302.220 ;
        RECT 63.250 302.450 63.870 302.635 ;
        RECT 94.850 302.450 95.470 302.635 ;
        RECT 63.250 302.220 95.470 302.450 ;
        RECT 63.250 302.035 63.870 302.220 ;
        RECT 94.850 302.035 95.470 302.220 ;
        RECT 95.700 302.450 96.320 302.635 ;
        RECT 127.300 302.450 127.920 302.635 ;
        RECT 95.700 302.220 127.920 302.450 ;
        RECT 95.700 302.035 96.320 302.220 ;
        RECT 127.300 302.035 127.920 302.220 ;
        RECT 128.150 302.450 128.770 302.635 ;
        RECT 159.750 302.450 160.370 302.635 ;
        RECT 128.150 302.220 160.370 302.450 ;
        RECT 128.150 302.035 128.770 302.220 ;
        RECT 159.750 302.035 160.370 302.220 ;
        RECT 58.400 301.955 60.020 301.965 ;
        RECT 90.850 301.955 92.470 301.965 ;
        RECT 123.300 301.955 124.920 301.965 ;
        RECT 155.750 301.955 157.370 301.965 ;
        RECT 31.650 301.585 62.170 301.955 ;
        RECT 64.100 301.585 94.620 301.955 ;
        RECT 96.550 301.585 127.070 301.955 ;
        RECT 129.000 301.585 159.520 301.955 ;
        RECT 31.650 300.865 62.170 301.245 ;
        RECT 64.100 300.865 94.620 301.245 ;
        RECT 96.550 300.865 127.070 301.245 ;
        RECT 129.000 300.865 159.520 301.245 ;
        RECT 30.800 300.610 31.420 300.795 ;
        RECT 62.400 300.610 63.020 300.795 ;
        RECT 30.800 300.380 63.020 300.610 ;
        RECT 30.800 300.195 31.420 300.380 ;
        RECT 62.400 300.195 63.020 300.380 ;
        RECT 63.250 300.610 63.870 300.795 ;
        RECT 94.850 300.610 95.470 300.795 ;
        RECT 63.250 300.380 95.470 300.610 ;
        RECT 63.250 300.195 63.870 300.380 ;
        RECT 94.850 300.195 95.470 300.380 ;
        RECT 95.700 300.610 96.320 300.795 ;
        RECT 127.300 300.610 127.920 300.795 ;
        RECT 95.700 300.380 127.920 300.610 ;
        RECT 95.700 300.195 96.320 300.380 ;
        RECT 127.300 300.195 127.920 300.380 ;
        RECT 128.150 300.610 128.770 300.795 ;
        RECT 159.750 300.610 160.370 300.795 ;
        RECT 128.150 300.380 160.370 300.610 ;
        RECT 128.150 300.195 128.770 300.380 ;
        RECT 159.750 300.195 160.370 300.380 ;
        RECT 54.560 300.115 56.180 300.125 ;
        RECT 87.010 300.115 88.630 300.125 ;
        RECT 119.460 300.115 121.080 300.125 ;
        RECT 151.910 300.115 153.530 300.125 ;
        RECT 31.650 299.745 62.170 300.115 ;
        RECT 64.100 299.745 94.620 300.115 ;
        RECT 96.550 299.745 127.070 300.115 ;
        RECT 129.000 299.745 159.520 300.115 ;
        RECT 31.660 298.950 62.160 299.390 ;
        RECT 64.110 298.950 94.610 299.390 ;
        RECT 96.560 298.950 127.060 299.390 ;
        RECT 129.010 298.950 159.510 299.390 ;
        RECT 31.650 298.220 62.170 298.600 ;
        RECT 64.100 298.220 94.620 298.600 ;
        RECT 96.550 298.220 127.070 298.600 ;
        RECT 129.000 298.220 159.520 298.600 ;
        RECT 30.800 297.965 31.420 298.150 ;
        RECT 62.400 297.965 63.020 298.150 ;
        RECT 30.800 297.735 63.020 297.965 ;
        RECT 30.800 297.550 31.420 297.735 ;
        RECT 62.400 297.550 63.020 297.735 ;
        RECT 63.250 297.965 63.870 298.150 ;
        RECT 94.850 297.965 95.470 298.150 ;
        RECT 63.250 297.735 95.470 297.965 ;
        RECT 63.250 297.550 63.870 297.735 ;
        RECT 94.850 297.550 95.470 297.735 ;
        RECT 95.700 297.965 96.320 298.150 ;
        RECT 127.300 297.965 127.920 298.150 ;
        RECT 95.700 297.735 127.920 297.965 ;
        RECT 95.700 297.550 96.320 297.735 ;
        RECT 127.300 297.550 127.920 297.735 ;
        RECT 128.150 297.965 128.770 298.150 ;
        RECT 159.750 297.965 160.370 298.150 ;
        RECT 128.150 297.735 160.370 297.965 ;
        RECT 128.150 297.550 128.770 297.735 ;
        RECT 159.750 297.550 160.370 297.735 ;
        RECT 50.720 297.470 52.340 297.480 ;
        RECT 83.170 297.470 84.790 297.480 ;
        RECT 115.620 297.470 117.240 297.480 ;
        RECT 148.070 297.470 149.690 297.480 ;
        RECT 31.650 297.100 62.170 297.470 ;
        RECT 64.100 297.100 94.620 297.470 ;
        RECT 96.550 297.100 127.070 297.470 ;
        RECT 129.000 297.100 159.520 297.470 ;
        RECT 31.650 296.380 62.170 296.760 ;
        RECT 64.100 296.380 94.620 296.760 ;
        RECT 96.550 296.380 127.070 296.760 ;
        RECT 129.000 296.380 159.520 296.760 ;
        RECT 30.800 296.125 31.420 296.310 ;
        RECT 62.400 296.125 63.020 296.310 ;
        RECT 30.800 295.895 63.020 296.125 ;
        RECT 30.800 295.710 31.420 295.895 ;
        RECT 62.400 295.710 63.020 295.895 ;
        RECT 63.250 296.125 63.870 296.310 ;
        RECT 94.850 296.125 95.470 296.310 ;
        RECT 63.250 295.895 95.470 296.125 ;
        RECT 63.250 295.710 63.870 295.895 ;
        RECT 94.850 295.710 95.470 295.895 ;
        RECT 95.700 296.125 96.320 296.310 ;
        RECT 127.300 296.125 127.920 296.310 ;
        RECT 95.700 295.895 127.920 296.125 ;
        RECT 95.700 295.710 96.320 295.895 ;
        RECT 127.300 295.710 127.920 295.895 ;
        RECT 128.150 296.125 128.770 296.310 ;
        RECT 159.750 296.125 160.370 296.310 ;
        RECT 128.150 295.895 160.370 296.125 ;
        RECT 128.150 295.710 128.770 295.895 ;
        RECT 159.750 295.710 160.370 295.895 ;
        RECT 46.880 295.630 48.500 295.640 ;
        RECT 79.330 295.630 80.950 295.640 ;
        RECT 111.780 295.630 113.400 295.640 ;
        RECT 144.230 295.630 145.850 295.640 ;
        RECT 31.650 295.260 62.170 295.630 ;
        RECT 64.100 295.260 94.620 295.630 ;
        RECT 96.550 295.260 127.070 295.630 ;
        RECT 129.000 295.260 159.520 295.630 ;
        RECT 31.650 294.540 62.170 294.920 ;
        RECT 64.100 294.540 94.620 294.920 ;
        RECT 96.550 294.540 127.070 294.920 ;
        RECT 129.000 294.540 159.520 294.920 ;
        RECT 30.800 294.285 31.420 294.470 ;
        RECT 62.400 294.285 63.020 294.470 ;
        RECT 30.800 294.055 63.020 294.285 ;
        RECT 30.800 293.870 31.420 294.055 ;
        RECT 62.400 293.870 63.020 294.055 ;
        RECT 63.250 294.285 63.870 294.470 ;
        RECT 94.850 294.285 95.470 294.470 ;
        RECT 63.250 294.055 95.470 294.285 ;
        RECT 63.250 293.870 63.870 294.055 ;
        RECT 94.850 293.870 95.470 294.055 ;
        RECT 95.700 294.285 96.320 294.470 ;
        RECT 127.300 294.285 127.920 294.470 ;
        RECT 95.700 294.055 127.920 294.285 ;
        RECT 95.700 293.870 96.320 294.055 ;
        RECT 127.300 293.870 127.920 294.055 ;
        RECT 128.150 294.285 128.770 294.470 ;
        RECT 159.750 294.285 160.370 294.470 ;
        RECT 128.150 294.055 160.370 294.285 ;
        RECT 128.150 293.870 128.770 294.055 ;
        RECT 159.750 293.870 160.370 294.055 ;
        RECT 43.040 293.790 44.660 293.800 ;
        RECT 75.490 293.790 77.110 293.800 ;
        RECT 107.940 293.790 109.560 293.800 ;
        RECT 140.390 293.790 142.010 293.800 ;
        RECT 31.650 293.420 62.170 293.790 ;
        RECT 64.100 293.420 94.620 293.790 ;
        RECT 96.550 293.420 127.070 293.790 ;
        RECT 129.000 293.420 159.520 293.790 ;
        RECT 31.660 292.625 62.160 293.065 ;
        RECT 64.110 292.625 94.610 293.065 ;
        RECT 96.560 292.625 127.060 293.065 ;
        RECT 129.010 292.625 159.510 293.065 ;
        RECT 31.650 291.895 62.170 292.275 ;
        RECT 64.100 291.895 94.620 292.275 ;
        RECT 96.550 291.895 127.070 292.275 ;
        RECT 129.000 291.895 159.520 292.275 ;
        RECT 30.800 291.640 31.420 291.825 ;
        RECT 62.400 291.640 63.020 291.825 ;
        RECT 30.800 291.410 63.020 291.640 ;
        RECT 30.800 291.225 31.420 291.410 ;
        RECT 62.400 291.225 63.020 291.410 ;
        RECT 63.250 291.640 63.870 291.825 ;
        RECT 94.850 291.640 95.470 291.825 ;
        RECT 63.250 291.410 95.470 291.640 ;
        RECT 63.250 291.225 63.870 291.410 ;
        RECT 94.850 291.225 95.470 291.410 ;
        RECT 95.700 291.640 96.320 291.825 ;
        RECT 127.300 291.640 127.920 291.825 ;
        RECT 95.700 291.410 127.920 291.640 ;
        RECT 95.700 291.225 96.320 291.410 ;
        RECT 127.300 291.225 127.920 291.410 ;
        RECT 128.150 291.640 128.770 291.825 ;
        RECT 159.750 291.640 160.370 291.825 ;
        RECT 128.150 291.410 160.370 291.640 ;
        RECT 128.150 291.225 128.770 291.410 ;
        RECT 159.750 291.225 160.370 291.410 ;
        RECT 39.200 291.145 40.820 291.155 ;
        RECT 71.650 291.145 73.270 291.155 ;
        RECT 104.100 291.145 105.720 291.155 ;
        RECT 136.550 291.145 138.170 291.155 ;
        RECT 31.650 290.775 62.170 291.145 ;
        RECT 64.100 290.775 94.620 291.145 ;
        RECT 96.550 290.775 127.070 291.145 ;
        RECT 129.000 290.775 159.520 291.145 ;
        RECT 31.650 290.055 62.170 290.435 ;
        RECT 64.100 290.055 94.620 290.435 ;
        RECT 96.550 290.055 127.070 290.435 ;
        RECT 129.000 290.055 159.520 290.435 ;
        RECT 30.800 289.800 31.420 289.985 ;
        RECT 62.400 289.800 63.020 289.985 ;
        RECT 30.800 289.570 63.020 289.800 ;
        RECT 30.800 289.385 31.420 289.570 ;
        RECT 62.400 289.385 63.020 289.570 ;
        RECT 63.250 289.800 63.870 289.985 ;
        RECT 94.850 289.800 95.470 289.985 ;
        RECT 63.250 289.570 95.470 289.800 ;
        RECT 63.250 289.385 63.870 289.570 ;
        RECT 94.850 289.385 95.470 289.570 ;
        RECT 95.700 289.800 96.320 289.985 ;
        RECT 127.300 289.800 127.920 289.985 ;
        RECT 95.700 289.570 127.920 289.800 ;
        RECT 95.700 289.385 96.320 289.570 ;
        RECT 127.300 289.385 127.920 289.570 ;
        RECT 128.150 289.800 128.770 289.985 ;
        RECT 159.750 289.800 160.370 289.985 ;
        RECT 128.150 289.570 160.370 289.800 ;
        RECT 128.150 289.385 128.770 289.570 ;
        RECT 159.750 289.385 160.370 289.570 ;
        RECT 35.360 289.305 36.980 289.315 ;
        RECT 67.810 289.305 69.430 289.315 ;
        RECT 100.260 289.305 101.880 289.315 ;
        RECT 132.710 289.305 134.330 289.315 ;
        RECT 31.650 288.935 62.170 289.305 ;
        RECT 64.100 288.935 94.620 289.305 ;
        RECT 96.550 288.935 127.070 289.305 ;
        RECT 129.000 288.935 159.520 289.305 ;
        RECT 31.650 288.215 62.170 288.595 ;
        RECT 64.100 288.215 94.620 288.595 ;
        RECT 96.550 288.215 127.070 288.595 ;
        RECT 129.000 288.215 159.520 288.595 ;
        RECT 30.800 287.960 31.420 288.145 ;
        RECT 62.400 287.960 63.020 288.145 ;
        RECT 30.800 287.730 63.020 287.960 ;
        RECT 30.800 287.545 31.420 287.730 ;
        RECT 62.400 287.545 63.020 287.730 ;
        RECT 63.250 287.960 63.870 288.145 ;
        RECT 94.850 287.960 95.470 288.145 ;
        RECT 63.250 287.730 95.470 287.960 ;
        RECT 63.250 287.545 63.870 287.730 ;
        RECT 94.850 287.545 95.470 287.730 ;
        RECT 95.700 287.960 96.320 288.145 ;
        RECT 127.300 287.960 127.920 288.145 ;
        RECT 95.700 287.730 127.920 287.960 ;
        RECT 95.700 287.545 96.320 287.730 ;
        RECT 127.300 287.545 127.920 287.730 ;
        RECT 128.150 287.960 128.770 288.145 ;
        RECT 159.750 287.960 160.370 288.145 ;
        RECT 128.150 287.730 160.370 287.960 ;
        RECT 128.150 287.545 128.770 287.730 ;
        RECT 159.750 287.545 160.370 287.730 ;
        RECT 31.650 287.095 62.170 287.465 ;
        RECT 64.100 287.095 94.620 287.465 ;
        RECT 96.550 287.095 127.070 287.465 ;
        RECT 129.000 287.095 159.520 287.465 ;
        RECT 25.090 284.745 27.380 285.085 ;
        RECT 28.125 284.745 29.610 285.085 ;
        RECT 25.090 284.110 25.690 284.745 ;
        RECT 25.090 283.880 26.670 284.110 ;
        RECT 25.090 281.840 25.690 283.880 ;
        RECT 27.100 283.650 27.460 283.735 ;
        RECT 25.970 283.420 27.460 283.650 ;
        RECT 25.970 283.270 26.330 283.420 ;
        RECT 25.920 282.635 26.870 283.040 ;
        RECT 25.090 281.610 26.380 281.840 ;
        RECT 25.090 280.650 25.690 281.610 ;
        RECT 26.610 281.290 26.870 282.635 ;
        RECT 27.100 281.985 27.460 283.420 ;
        RECT 27.690 282.085 28.040 283.285 ;
        RECT 28.400 282.675 28.780 284.320 ;
        RECT 27.480 281.290 27.830 281.350 ;
        RECT 28.400 281.290 28.740 281.895 ;
        RECT 26.610 281.030 28.740 281.290 ;
        RECT 27.480 280.970 27.830 281.030 ;
        RECT 29.010 280.750 29.610 284.745 ;
        RECT 31.455 284.310 33.205 287.095 ;
        RECT 33.845 284.310 34.655 285.310 ;
        RECT 35.295 284.310 37.045 286.605 ;
        RECT 37.685 284.310 38.495 285.310 ;
        RECT 39.135 284.310 40.885 286.605 ;
        RECT 41.525 284.310 42.335 285.310 ;
        RECT 42.975 284.310 44.725 286.605 ;
        RECT 45.365 284.310 46.175 285.310 ;
        RECT 46.815 284.310 48.565 286.605 ;
        RECT 49.205 284.310 50.015 285.310 ;
        RECT 50.655 284.310 52.405 286.605 ;
        RECT 53.045 284.310 53.855 285.310 ;
        RECT 54.495 284.310 56.245 286.605 ;
        RECT 56.885 284.310 57.695 285.310 ;
        RECT 58.335 284.310 60.085 286.605 ;
        RECT 60.725 284.310 61.535 285.310 ;
        RECT 63.905 284.310 65.655 287.095 ;
        RECT 66.295 284.310 67.105 285.310 ;
        RECT 67.745 284.310 69.495 286.605 ;
        RECT 70.135 284.310 70.945 285.310 ;
        RECT 71.585 284.310 73.335 286.605 ;
        RECT 73.975 284.310 74.785 285.310 ;
        RECT 75.425 284.310 77.175 286.605 ;
        RECT 77.815 284.310 78.625 285.310 ;
        RECT 79.265 284.310 81.015 286.605 ;
        RECT 81.655 284.310 82.465 285.310 ;
        RECT 83.105 284.310 84.855 286.605 ;
        RECT 85.495 284.310 86.305 285.310 ;
        RECT 86.945 284.310 88.695 286.605 ;
        RECT 89.335 284.310 90.145 285.310 ;
        RECT 90.785 284.310 92.535 286.605 ;
        RECT 93.175 284.310 93.985 285.310 ;
        RECT 96.355 284.310 98.105 287.095 ;
        RECT 98.745 284.310 99.555 285.310 ;
        RECT 100.195 284.310 101.945 286.605 ;
        RECT 102.585 284.310 103.395 285.310 ;
        RECT 104.035 284.310 105.785 286.605 ;
        RECT 106.425 284.310 107.235 285.310 ;
        RECT 107.875 284.310 109.625 286.605 ;
        RECT 110.265 284.310 111.075 285.310 ;
        RECT 111.715 284.310 113.465 286.605 ;
        RECT 114.105 284.310 114.915 285.310 ;
        RECT 115.555 284.310 117.305 286.605 ;
        RECT 117.945 284.310 118.755 285.310 ;
        RECT 119.395 284.310 121.145 286.605 ;
        RECT 121.785 284.310 122.595 285.310 ;
        RECT 123.235 284.310 124.985 286.605 ;
        RECT 125.625 284.310 126.435 285.310 ;
        RECT 128.805 284.310 130.555 287.095 ;
        RECT 131.195 284.310 132.005 285.310 ;
        RECT 132.645 284.310 134.395 286.605 ;
        RECT 135.035 284.310 135.845 285.310 ;
        RECT 136.485 284.310 138.235 286.605 ;
        RECT 138.875 284.310 139.685 285.310 ;
        RECT 140.325 284.310 142.075 286.605 ;
        RECT 142.715 284.310 143.525 285.310 ;
        RECT 144.165 284.310 145.915 286.605 ;
        RECT 146.555 284.310 147.365 285.310 ;
        RECT 148.005 284.310 149.755 286.605 ;
        RECT 150.395 284.310 151.205 285.310 ;
        RECT 151.845 284.310 153.595 286.605 ;
        RECT 154.235 284.310 155.045 285.310 ;
        RECT 155.685 284.310 157.435 286.605 ;
        RECT 158.075 284.310 158.885 285.310 ;
        RECT 161.300 284.500 161.670 303.010 ;
        RECT 162.320 299.375 162.690 303.010 ;
        RECT 162.315 298.995 162.695 299.375 ;
        RECT 162.320 296.375 162.690 298.995 ;
        RECT 162.315 295.995 162.695 296.375 ;
        RECT 162.320 293.375 162.690 295.995 ;
        RECT 162.315 292.995 162.695 293.375 ;
        RECT 162.320 290.375 162.690 292.995 ;
        RECT 162.315 289.995 162.695 290.375 ;
        RECT 162.320 287.375 162.690 289.995 ;
        RECT 162.315 286.995 162.695 287.375 ;
        RECT 161.300 284.120 161.680 284.500 ;
        RECT 161.300 283.050 161.670 284.120 ;
        RECT 31.925 281.860 32.735 282.860 ;
        RECT 25.090 280.420 26.780 280.650 ;
        RECT 28.150 280.520 29.610 280.750 ;
        RECT 25.090 278.410 25.690 280.420 ;
        RECT 27.110 279.960 28.110 280.285 ;
        RECT 25.920 279.400 28.780 279.730 ;
        RECT 25.090 278.180 26.780 278.410 ;
        RECT 25.090 276.170 25.690 278.180 ;
        RECT 27.495 278.045 27.760 279.400 ;
        RECT 29.010 278.510 29.610 280.520 ;
        RECT 33.375 280.030 35.125 282.860 ;
        RECT 35.765 281.860 36.575 282.860 ;
        RECT 37.215 280.565 38.965 282.860 ;
        RECT 39.605 281.860 40.415 282.860 ;
        RECT 41.055 280.565 42.805 282.860 ;
        RECT 43.445 281.860 44.255 282.860 ;
        RECT 44.895 280.565 46.645 282.860 ;
        RECT 47.285 281.860 48.095 282.860 ;
        RECT 48.735 280.565 50.485 282.860 ;
        RECT 51.125 281.860 51.935 282.860 ;
        RECT 52.575 280.565 54.325 282.860 ;
        RECT 54.965 281.860 55.775 282.860 ;
        RECT 56.415 280.565 58.165 282.860 ;
        RECT 58.805 281.860 59.615 282.860 ;
        RECT 60.255 280.565 62.005 282.860 ;
        RECT 64.375 281.860 65.185 282.860 ;
        RECT 65.825 280.030 67.575 282.860 ;
        RECT 68.215 281.860 69.025 282.860 ;
        RECT 69.665 280.565 71.415 282.860 ;
        RECT 72.055 281.860 72.865 282.860 ;
        RECT 73.505 280.565 75.255 282.860 ;
        RECT 75.895 281.860 76.705 282.860 ;
        RECT 77.345 280.565 79.095 282.860 ;
        RECT 79.735 281.860 80.545 282.860 ;
        RECT 81.185 280.565 82.935 282.860 ;
        RECT 83.575 281.860 84.385 282.860 ;
        RECT 85.025 280.565 86.775 282.860 ;
        RECT 87.415 281.860 88.225 282.860 ;
        RECT 88.865 280.565 90.615 282.860 ;
        RECT 91.255 281.860 92.065 282.860 ;
        RECT 92.705 280.565 94.455 282.860 ;
        RECT 96.825 281.860 97.635 282.860 ;
        RECT 98.275 280.030 100.025 282.860 ;
        RECT 100.665 281.860 101.475 282.860 ;
        RECT 102.115 280.565 103.865 282.860 ;
        RECT 104.505 281.860 105.315 282.860 ;
        RECT 105.955 280.565 107.705 282.860 ;
        RECT 108.345 281.860 109.155 282.860 ;
        RECT 109.795 280.565 111.545 282.860 ;
        RECT 112.185 281.860 112.995 282.860 ;
        RECT 113.635 280.565 115.385 282.860 ;
        RECT 116.025 281.860 116.835 282.860 ;
        RECT 117.475 280.565 119.225 282.860 ;
        RECT 119.865 281.860 120.675 282.860 ;
        RECT 121.315 280.565 123.065 282.860 ;
        RECT 123.705 281.860 124.515 282.860 ;
        RECT 125.155 280.565 126.905 282.860 ;
        RECT 129.275 281.860 130.085 282.860 ;
        RECT 130.725 280.030 132.475 282.860 ;
        RECT 133.115 281.860 133.925 282.860 ;
        RECT 134.565 280.565 136.315 282.860 ;
        RECT 136.955 281.860 137.765 282.860 ;
        RECT 138.405 280.565 140.155 282.860 ;
        RECT 140.795 281.860 141.605 282.860 ;
        RECT 142.245 280.565 143.995 282.860 ;
        RECT 144.635 281.860 145.445 282.860 ;
        RECT 146.085 280.565 147.835 282.860 ;
        RECT 148.475 281.860 149.285 282.860 ;
        RECT 149.925 280.565 151.675 282.860 ;
        RECT 152.315 281.860 153.125 282.860 ;
        RECT 153.765 280.565 155.515 282.860 ;
        RECT 156.155 281.860 156.965 282.860 ;
        RECT 157.605 280.565 159.355 282.860 ;
        RECT 161.300 282.670 161.680 283.050 ;
        RECT 31.650 279.660 62.170 280.030 ;
        RECT 64.100 279.660 94.620 280.030 ;
        RECT 96.550 279.660 127.070 280.030 ;
        RECT 129.000 279.660 159.520 280.030 ;
        RECT 30.800 279.395 31.420 279.580 ;
        RECT 62.400 279.395 63.020 279.580 ;
        RECT 30.800 279.165 63.020 279.395 ;
        RECT 30.800 278.980 31.420 279.165 ;
        RECT 62.400 278.980 63.020 279.165 ;
        RECT 63.250 279.395 63.870 279.580 ;
        RECT 94.850 279.395 95.470 279.580 ;
        RECT 63.250 279.165 95.470 279.395 ;
        RECT 63.250 278.980 63.870 279.165 ;
        RECT 94.850 278.980 95.470 279.165 ;
        RECT 95.700 279.395 96.320 279.580 ;
        RECT 127.300 279.395 127.920 279.580 ;
        RECT 95.700 279.165 127.920 279.395 ;
        RECT 95.700 278.980 96.320 279.165 ;
        RECT 127.300 278.980 127.920 279.165 ;
        RECT 128.150 279.395 128.770 279.580 ;
        RECT 159.750 279.395 160.370 279.580 ;
        RECT 128.150 279.165 160.370 279.395 ;
        RECT 128.150 278.980 128.770 279.165 ;
        RECT 159.750 278.980 160.370 279.165 ;
        RECT 31.650 278.530 62.170 278.910 ;
        RECT 64.100 278.530 94.620 278.910 ;
        RECT 96.550 278.530 127.070 278.910 ;
        RECT 129.000 278.530 159.520 278.910 ;
        RECT 28.150 278.280 29.610 278.510 ;
        RECT 27.110 277.720 28.110 278.045 ;
        RECT 25.920 277.160 28.780 277.490 ;
        RECT 29.010 276.270 29.610 278.280 ;
        RECT 31.650 277.820 62.170 278.190 ;
        RECT 64.100 277.820 94.620 278.190 ;
        RECT 96.550 277.820 127.070 278.190 ;
        RECT 129.000 277.820 159.520 278.190 ;
        RECT 37.280 277.810 38.900 277.820 ;
        RECT 69.730 277.810 71.350 277.820 ;
        RECT 102.180 277.810 103.800 277.820 ;
        RECT 134.630 277.810 136.250 277.820 ;
        RECT 30.800 277.555 31.420 277.740 ;
        RECT 62.400 277.555 63.020 277.740 ;
        RECT 30.800 277.325 63.020 277.555 ;
        RECT 30.800 277.140 31.420 277.325 ;
        RECT 62.400 277.140 63.020 277.325 ;
        RECT 63.250 277.555 63.870 277.740 ;
        RECT 94.850 277.555 95.470 277.740 ;
        RECT 63.250 277.325 95.470 277.555 ;
        RECT 63.250 277.140 63.870 277.325 ;
        RECT 94.850 277.140 95.470 277.325 ;
        RECT 95.700 277.555 96.320 277.740 ;
        RECT 127.300 277.555 127.920 277.740 ;
        RECT 95.700 277.325 127.920 277.555 ;
        RECT 95.700 277.140 96.320 277.325 ;
        RECT 127.300 277.140 127.920 277.325 ;
        RECT 128.150 277.555 128.770 277.740 ;
        RECT 159.750 277.555 160.370 277.740 ;
        RECT 128.150 277.325 160.370 277.555 ;
        RECT 128.150 277.140 128.770 277.325 ;
        RECT 159.750 277.140 160.370 277.325 ;
        RECT 31.650 276.690 62.170 277.070 ;
        RECT 64.100 276.690 94.620 277.070 ;
        RECT 96.550 276.690 127.070 277.070 ;
        RECT 129.000 276.690 159.520 277.070 ;
        RECT 25.090 275.940 26.780 276.170 ;
        RECT 28.150 276.040 29.610 276.270 ;
        RECT 25.090 273.885 25.690 275.940 ;
        RECT 27.110 275.480 28.110 275.805 ;
        RECT 29.010 273.885 29.610 276.040 ;
        RECT 31.650 275.975 62.170 276.345 ;
        RECT 64.100 275.975 94.620 276.345 ;
        RECT 96.550 275.975 127.070 276.345 ;
        RECT 129.000 275.975 159.520 276.345 ;
        RECT 41.120 275.965 42.740 275.975 ;
        RECT 73.570 275.965 75.190 275.975 ;
        RECT 106.020 275.965 107.640 275.975 ;
        RECT 138.470 275.965 140.090 275.975 ;
        RECT 30.800 275.710 31.420 275.895 ;
        RECT 62.400 275.710 63.020 275.895 ;
        RECT 30.800 275.480 63.020 275.710 ;
        RECT 30.800 275.295 31.420 275.480 ;
        RECT 62.400 275.295 63.020 275.480 ;
        RECT 63.250 275.710 63.870 275.895 ;
        RECT 94.850 275.710 95.470 275.895 ;
        RECT 63.250 275.480 95.470 275.710 ;
        RECT 63.250 275.295 63.870 275.480 ;
        RECT 94.850 275.295 95.470 275.480 ;
        RECT 95.700 275.710 96.320 275.895 ;
        RECT 127.300 275.710 127.920 275.895 ;
        RECT 95.700 275.480 127.920 275.710 ;
        RECT 95.700 275.295 96.320 275.480 ;
        RECT 127.300 275.295 127.920 275.480 ;
        RECT 128.150 275.710 128.770 275.895 ;
        RECT 159.750 275.710 160.370 275.895 ;
        RECT 128.150 275.480 160.370 275.710 ;
        RECT 128.150 275.295 128.770 275.480 ;
        RECT 159.750 275.295 160.370 275.480 ;
        RECT 31.650 274.845 62.170 275.225 ;
        RECT 64.100 274.845 94.620 275.225 ;
        RECT 96.550 274.845 127.070 275.225 ;
        RECT 129.000 274.845 159.520 275.225 ;
        RECT 31.660 274.055 62.160 274.495 ;
        RECT 64.110 274.055 94.610 274.495 ;
        RECT 96.560 274.055 127.060 274.495 ;
        RECT 129.010 274.055 159.510 274.495 ;
        RECT 25.090 273.545 27.380 273.885 ;
        RECT 28.125 273.545 29.610 273.885 ;
        RECT 25.090 245.700 25.690 273.545 ;
        RECT 29.010 245.700 29.610 273.545 ;
        RECT 31.650 273.335 62.170 273.705 ;
        RECT 64.100 273.335 94.620 273.705 ;
        RECT 96.550 273.335 127.070 273.705 ;
        RECT 129.000 273.335 159.520 273.705 ;
        RECT 44.960 273.325 46.580 273.335 ;
        RECT 77.410 273.325 79.030 273.335 ;
        RECT 109.860 273.325 111.480 273.335 ;
        RECT 142.310 273.325 143.930 273.335 ;
        RECT 30.800 273.070 31.420 273.255 ;
        RECT 62.400 273.070 63.020 273.255 ;
        RECT 30.800 272.840 63.020 273.070 ;
        RECT 30.800 272.655 31.420 272.840 ;
        RECT 62.400 272.655 63.020 272.840 ;
        RECT 63.250 273.070 63.870 273.255 ;
        RECT 94.850 273.070 95.470 273.255 ;
        RECT 63.250 272.840 95.470 273.070 ;
        RECT 63.250 272.655 63.870 272.840 ;
        RECT 94.850 272.655 95.470 272.840 ;
        RECT 95.700 273.070 96.320 273.255 ;
        RECT 127.300 273.070 127.920 273.255 ;
        RECT 95.700 272.840 127.920 273.070 ;
        RECT 95.700 272.655 96.320 272.840 ;
        RECT 127.300 272.655 127.920 272.840 ;
        RECT 128.150 273.070 128.770 273.255 ;
        RECT 159.750 273.070 160.370 273.255 ;
        RECT 128.150 272.840 160.370 273.070 ;
        RECT 128.150 272.655 128.770 272.840 ;
        RECT 159.750 272.655 160.370 272.840 ;
        RECT 31.650 272.205 62.170 272.585 ;
        RECT 64.100 272.205 94.620 272.585 ;
        RECT 96.550 272.205 127.070 272.585 ;
        RECT 129.000 272.205 159.520 272.585 ;
        RECT 31.650 271.495 62.170 271.865 ;
        RECT 64.100 271.495 94.620 271.865 ;
        RECT 96.550 271.495 127.070 271.865 ;
        RECT 129.000 271.495 159.520 271.865 ;
        RECT 48.800 271.485 50.420 271.495 ;
        RECT 81.250 271.485 82.870 271.495 ;
        RECT 113.700 271.485 115.320 271.495 ;
        RECT 146.150 271.485 147.770 271.495 ;
        RECT 30.800 271.230 31.420 271.415 ;
        RECT 62.400 271.230 63.020 271.415 ;
        RECT 30.800 271.000 63.020 271.230 ;
        RECT 30.800 270.815 31.420 271.000 ;
        RECT 62.400 270.815 63.020 271.000 ;
        RECT 63.250 271.230 63.870 271.415 ;
        RECT 94.850 271.230 95.470 271.415 ;
        RECT 63.250 271.000 95.470 271.230 ;
        RECT 63.250 270.815 63.870 271.000 ;
        RECT 94.850 270.815 95.470 271.000 ;
        RECT 95.700 271.230 96.320 271.415 ;
        RECT 127.300 271.230 127.920 271.415 ;
        RECT 95.700 271.000 127.920 271.230 ;
        RECT 95.700 270.815 96.320 271.000 ;
        RECT 127.300 270.815 127.920 271.000 ;
        RECT 128.150 271.230 128.770 271.415 ;
        RECT 159.750 271.230 160.370 271.415 ;
        RECT 128.150 271.000 160.370 271.230 ;
        RECT 128.150 270.815 128.770 271.000 ;
        RECT 159.750 270.815 160.370 271.000 ;
        RECT 31.650 270.365 62.170 270.745 ;
        RECT 64.100 270.365 94.620 270.745 ;
        RECT 96.550 270.365 127.070 270.745 ;
        RECT 129.000 270.365 159.520 270.745 ;
        RECT 31.650 269.650 62.170 270.020 ;
        RECT 64.100 269.650 94.620 270.020 ;
        RECT 96.550 269.650 127.070 270.020 ;
        RECT 129.000 269.650 159.520 270.020 ;
        RECT 52.640 269.640 54.260 269.650 ;
        RECT 85.090 269.640 86.710 269.650 ;
        RECT 117.540 269.640 119.160 269.650 ;
        RECT 149.990 269.640 151.610 269.650 ;
        RECT 30.800 269.385 31.420 269.570 ;
        RECT 62.400 269.385 63.020 269.570 ;
        RECT 30.800 269.155 63.020 269.385 ;
        RECT 30.800 268.970 31.420 269.155 ;
        RECT 62.400 268.970 63.020 269.155 ;
        RECT 63.250 269.385 63.870 269.570 ;
        RECT 94.850 269.385 95.470 269.570 ;
        RECT 63.250 269.155 95.470 269.385 ;
        RECT 63.250 268.970 63.870 269.155 ;
        RECT 94.850 268.970 95.470 269.155 ;
        RECT 95.700 269.385 96.320 269.570 ;
        RECT 127.300 269.385 127.920 269.570 ;
        RECT 95.700 269.155 127.920 269.385 ;
        RECT 95.700 268.970 96.320 269.155 ;
        RECT 127.300 268.970 127.920 269.155 ;
        RECT 128.150 269.385 128.770 269.570 ;
        RECT 159.750 269.385 160.370 269.570 ;
        RECT 128.150 269.155 160.370 269.385 ;
        RECT 128.150 268.970 128.770 269.155 ;
        RECT 159.750 268.970 160.370 269.155 ;
        RECT 31.650 268.520 62.170 268.900 ;
        RECT 64.100 268.520 94.620 268.900 ;
        RECT 96.550 268.520 127.070 268.900 ;
        RECT 129.000 268.520 159.520 268.900 ;
        RECT 31.660 267.730 62.160 268.170 ;
        RECT 64.110 267.730 94.610 268.170 ;
        RECT 96.560 267.730 127.060 268.170 ;
        RECT 129.010 267.730 159.510 268.170 ;
        RECT 31.650 267.010 62.170 267.380 ;
        RECT 64.100 267.010 94.620 267.380 ;
        RECT 96.550 267.010 127.070 267.380 ;
        RECT 129.000 267.010 159.520 267.380 ;
        RECT 56.480 267.000 58.100 267.010 ;
        RECT 88.930 267.000 90.550 267.010 ;
        RECT 121.380 267.000 123.000 267.010 ;
        RECT 153.830 267.000 155.450 267.010 ;
        RECT 30.800 266.745 31.420 266.930 ;
        RECT 62.400 266.745 63.020 266.930 ;
        RECT 30.800 266.515 63.020 266.745 ;
        RECT 30.800 266.330 31.420 266.515 ;
        RECT 62.400 266.330 63.020 266.515 ;
        RECT 63.250 266.745 63.870 266.930 ;
        RECT 94.850 266.745 95.470 266.930 ;
        RECT 63.250 266.515 95.470 266.745 ;
        RECT 63.250 266.330 63.870 266.515 ;
        RECT 94.850 266.330 95.470 266.515 ;
        RECT 95.700 266.745 96.320 266.930 ;
        RECT 127.300 266.745 127.920 266.930 ;
        RECT 95.700 266.515 127.920 266.745 ;
        RECT 95.700 266.330 96.320 266.515 ;
        RECT 127.300 266.330 127.920 266.515 ;
        RECT 128.150 266.745 128.770 266.930 ;
        RECT 159.750 266.745 160.370 266.930 ;
        RECT 128.150 266.515 160.370 266.745 ;
        RECT 128.150 266.330 128.770 266.515 ;
        RECT 159.750 266.330 160.370 266.515 ;
        RECT 31.650 265.880 62.170 266.260 ;
        RECT 64.100 265.880 94.620 266.260 ;
        RECT 96.550 265.880 127.070 266.260 ;
        RECT 129.000 265.880 159.520 266.260 ;
        RECT 31.650 265.170 62.170 265.540 ;
        RECT 64.100 265.170 94.620 265.540 ;
        RECT 96.550 265.170 127.070 265.540 ;
        RECT 129.000 265.170 159.520 265.540 ;
        RECT 60.320 265.160 61.940 265.170 ;
        RECT 92.770 265.160 94.390 265.170 ;
        RECT 125.220 265.160 126.840 265.170 ;
        RECT 157.670 265.160 159.290 265.170 ;
        RECT 30.800 264.905 31.420 265.090 ;
        RECT 62.400 264.905 63.020 265.090 ;
        RECT 30.800 264.675 63.020 264.905 ;
        RECT 30.800 264.490 31.420 264.675 ;
        RECT 62.400 264.490 63.020 264.675 ;
        RECT 63.250 264.905 63.870 265.090 ;
        RECT 94.850 264.905 95.470 265.090 ;
        RECT 63.250 264.675 95.470 264.905 ;
        RECT 63.250 264.490 63.870 264.675 ;
        RECT 94.850 264.490 95.470 264.675 ;
        RECT 95.700 264.905 96.320 265.090 ;
        RECT 127.300 264.905 127.920 265.090 ;
        RECT 95.700 264.675 127.920 264.905 ;
        RECT 95.700 264.490 96.320 264.675 ;
        RECT 127.300 264.490 127.920 264.675 ;
        RECT 128.150 264.905 128.770 265.090 ;
        RECT 159.750 264.905 160.370 265.090 ;
        RECT 128.150 264.675 160.370 264.905 ;
        RECT 161.300 264.740 161.670 282.670 ;
        RECT 162.320 281.375 162.690 286.995 ;
        RECT 163.340 284.500 163.710 303.010 ;
        RECT 164.360 299.375 164.730 303.010 ;
        RECT 164.355 298.995 164.735 299.375 ;
        RECT 164.360 296.375 164.730 298.995 ;
        RECT 164.355 295.995 164.735 296.375 ;
        RECT 164.360 293.375 164.730 295.995 ;
        RECT 164.355 292.995 164.735 293.375 ;
        RECT 164.360 290.375 164.730 292.995 ;
        RECT 164.355 289.995 164.735 290.375 ;
        RECT 164.360 287.375 164.730 289.995 ;
        RECT 164.355 286.995 164.735 287.375 ;
        RECT 163.340 284.120 163.720 284.500 ;
        RECT 163.340 283.050 163.710 284.120 ;
        RECT 163.340 282.670 163.720 283.050 ;
        RECT 162.315 280.995 162.695 281.375 ;
        RECT 162.320 278.375 162.690 280.995 ;
        RECT 162.315 277.995 162.695 278.375 ;
        RECT 162.320 275.375 162.690 277.995 ;
        RECT 162.315 274.995 162.695 275.375 ;
        RECT 162.320 272.375 162.690 274.995 ;
        RECT 162.315 271.995 162.695 272.375 ;
        RECT 162.320 269.375 162.690 271.995 ;
        RECT 162.315 268.995 162.695 269.375 ;
        RECT 162.320 266.375 162.690 268.995 ;
        RECT 162.315 265.995 162.695 266.375 ;
        RECT 162.320 264.740 162.690 265.995 ;
        RECT 163.340 264.740 163.710 282.670 ;
        RECT 164.360 281.375 164.730 286.995 ;
        RECT 164.355 280.995 164.735 281.375 ;
        RECT 164.360 278.375 164.730 280.995 ;
        RECT 164.355 277.995 164.735 278.375 ;
        RECT 164.360 275.375 164.730 277.995 ;
        RECT 164.355 274.995 164.735 275.375 ;
        RECT 164.360 272.375 164.730 274.995 ;
        RECT 164.355 271.995 164.735 272.375 ;
        RECT 164.360 269.375 164.730 271.995 ;
        RECT 164.355 268.995 164.735 269.375 ;
        RECT 164.360 266.375 164.730 268.995 ;
        RECT 164.355 265.995 164.735 266.375 ;
        RECT 164.360 264.740 164.730 265.995 ;
        RECT 165.380 264.740 165.760 303.010 ;
        RECT 166.110 264.750 166.550 303.000 ;
        RECT 128.150 264.490 128.770 264.675 ;
        RECT 159.750 264.490 160.370 264.675 ;
        RECT 31.650 264.040 62.170 264.420 ;
        RECT 64.100 264.040 94.620 264.420 ;
        RECT 96.550 264.040 127.070 264.420 ;
        RECT 129.000 264.040 159.520 264.420 ;
        RECT 31.650 263.320 62.170 263.700 ;
        RECT 64.100 263.320 94.620 263.700 ;
        RECT 96.550 263.320 127.070 263.700 ;
        RECT 129.000 263.320 159.520 263.700 ;
        RECT 30.800 263.065 31.420 263.250 ;
        RECT 62.400 263.065 63.020 263.250 ;
        RECT 30.800 262.835 63.020 263.065 ;
        RECT 30.800 262.650 31.420 262.835 ;
        RECT 62.400 262.650 63.020 262.835 ;
        RECT 63.250 263.065 63.870 263.250 ;
        RECT 94.850 263.065 95.470 263.250 ;
        RECT 63.250 262.835 95.470 263.065 ;
        RECT 63.250 262.650 63.870 262.835 ;
        RECT 94.850 262.650 95.470 262.835 ;
        RECT 95.700 263.065 96.320 263.250 ;
        RECT 127.300 263.065 127.920 263.250 ;
        RECT 95.700 262.835 127.920 263.065 ;
        RECT 95.700 262.650 96.320 262.835 ;
        RECT 127.300 262.650 127.920 262.835 ;
        RECT 128.150 263.065 128.770 263.250 ;
        RECT 159.750 263.065 160.370 263.250 ;
        RECT 128.150 262.835 160.370 263.065 ;
        RECT 128.150 262.650 128.770 262.835 ;
        RECT 159.750 262.650 160.370 262.835 ;
        RECT 58.400 262.570 60.020 262.580 ;
        RECT 90.850 262.570 92.470 262.580 ;
        RECT 123.300 262.570 124.920 262.580 ;
        RECT 155.750 262.570 157.370 262.580 ;
        RECT 31.650 262.200 62.170 262.570 ;
        RECT 64.100 262.200 94.620 262.570 ;
        RECT 96.550 262.200 127.070 262.570 ;
        RECT 129.000 262.200 159.520 262.570 ;
        RECT 31.650 261.480 62.170 261.860 ;
        RECT 64.100 261.480 94.620 261.860 ;
        RECT 96.550 261.480 127.070 261.860 ;
        RECT 129.000 261.480 159.520 261.860 ;
        RECT 30.800 261.225 31.420 261.410 ;
        RECT 62.400 261.225 63.020 261.410 ;
        RECT 30.800 260.995 63.020 261.225 ;
        RECT 30.800 260.810 31.420 260.995 ;
        RECT 62.400 260.810 63.020 260.995 ;
        RECT 63.250 261.225 63.870 261.410 ;
        RECT 94.850 261.225 95.470 261.410 ;
        RECT 63.250 260.995 95.470 261.225 ;
        RECT 63.250 260.810 63.870 260.995 ;
        RECT 94.850 260.810 95.470 260.995 ;
        RECT 95.700 261.225 96.320 261.410 ;
        RECT 127.300 261.225 127.920 261.410 ;
        RECT 95.700 260.995 127.920 261.225 ;
        RECT 95.700 260.810 96.320 260.995 ;
        RECT 127.300 260.810 127.920 260.995 ;
        RECT 128.150 261.225 128.770 261.410 ;
        RECT 159.750 261.225 160.370 261.410 ;
        RECT 128.150 260.995 160.370 261.225 ;
        RECT 128.150 260.810 128.770 260.995 ;
        RECT 159.750 260.810 160.370 260.995 ;
        RECT 54.560 260.730 56.180 260.740 ;
        RECT 87.010 260.730 88.630 260.740 ;
        RECT 119.460 260.730 121.080 260.740 ;
        RECT 151.910 260.730 153.530 260.740 ;
        RECT 31.650 260.360 62.170 260.730 ;
        RECT 64.100 260.360 94.620 260.730 ;
        RECT 96.550 260.360 127.070 260.730 ;
        RECT 129.000 260.360 159.520 260.730 ;
        RECT 31.660 259.565 62.160 260.005 ;
        RECT 64.110 259.565 94.610 260.005 ;
        RECT 96.560 259.565 127.060 260.005 ;
        RECT 129.010 259.565 159.510 260.005 ;
        RECT 31.650 258.835 62.170 259.215 ;
        RECT 64.100 258.835 94.620 259.215 ;
        RECT 96.550 258.835 127.070 259.215 ;
        RECT 129.000 258.835 159.520 259.215 ;
        RECT 30.800 258.580 31.420 258.765 ;
        RECT 62.400 258.580 63.020 258.765 ;
        RECT 30.800 258.350 63.020 258.580 ;
        RECT 30.800 258.165 31.420 258.350 ;
        RECT 62.400 258.165 63.020 258.350 ;
        RECT 63.250 258.580 63.870 258.765 ;
        RECT 94.850 258.580 95.470 258.765 ;
        RECT 63.250 258.350 95.470 258.580 ;
        RECT 63.250 258.165 63.870 258.350 ;
        RECT 94.850 258.165 95.470 258.350 ;
        RECT 95.700 258.580 96.320 258.765 ;
        RECT 127.300 258.580 127.920 258.765 ;
        RECT 95.700 258.350 127.920 258.580 ;
        RECT 95.700 258.165 96.320 258.350 ;
        RECT 127.300 258.165 127.920 258.350 ;
        RECT 128.150 258.580 128.770 258.765 ;
        RECT 159.750 258.580 160.370 258.765 ;
        RECT 128.150 258.350 160.370 258.580 ;
        RECT 128.150 258.165 128.770 258.350 ;
        RECT 159.750 258.165 160.370 258.350 ;
        RECT 50.720 258.085 52.340 258.095 ;
        RECT 83.170 258.085 84.790 258.095 ;
        RECT 115.620 258.085 117.240 258.095 ;
        RECT 148.070 258.085 149.690 258.095 ;
        RECT 31.650 257.715 62.170 258.085 ;
        RECT 64.100 257.715 94.620 258.085 ;
        RECT 96.550 257.715 127.070 258.085 ;
        RECT 129.000 257.715 159.520 258.085 ;
        RECT 31.650 256.995 62.170 257.375 ;
        RECT 64.100 256.995 94.620 257.375 ;
        RECT 96.550 256.995 127.070 257.375 ;
        RECT 129.000 256.995 159.520 257.375 ;
        RECT 30.800 256.740 31.420 256.925 ;
        RECT 62.400 256.740 63.020 256.925 ;
        RECT 30.800 256.510 63.020 256.740 ;
        RECT 30.800 256.325 31.420 256.510 ;
        RECT 62.400 256.325 63.020 256.510 ;
        RECT 63.250 256.740 63.870 256.925 ;
        RECT 94.850 256.740 95.470 256.925 ;
        RECT 63.250 256.510 95.470 256.740 ;
        RECT 63.250 256.325 63.870 256.510 ;
        RECT 94.850 256.325 95.470 256.510 ;
        RECT 95.700 256.740 96.320 256.925 ;
        RECT 127.300 256.740 127.920 256.925 ;
        RECT 95.700 256.510 127.920 256.740 ;
        RECT 95.700 256.325 96.320 256.510 ;
        RECT 127.300 256.325 127.920 256.510 ;
        RECT 128.150 256.740 128.770 256.925 ;
        RECT 159.750 256.740 160.370 256.925 ;
        RECT 128.150 256.510 160.370 256.740 ;
        RECT 128.150 256.325 128.770 256.510 ;
        RECT 159.750 256.325 160.370 256.510 ;
        RECT 46.880 256.245 48.500 256.255 ;
        RECT 79.330 256.245 80.950 256.255 ;
        RECT 111.780 256.245 113.400 256.255 ;
        RECT 144.230 256.245 145.850 256.255 ;
        RECT 31.650 255.875 62.170 256.245 ;
        RECT 64.100 255.875 94.620 256.245 ;
        RECT 96.550 255.875 127.070 256.245 ;
        RECT 129.000 255.875 159.520 256.245 ;
        RECT 31.650 255.155 62.170 255.535 ;
        RECT 64.100 255.155 94.620 255.535 ;
        RECT 96.550 255.155 127.070 255.535 ;
        RECT 129.000 255.155 159.520 255.535 ;
        RECT 30.800 254.900 31.420 255.085 ;
        RECT 62.400 254.900 63.020 255.085 ;
        RECT 30.800 254.670 63.020 254.900 ;
        RECT 30.800 254.485 31.420 254.670 ;
        RECT 62.400 254.485 63.020 254.670 ;
        RECT 63.250 254.900 63.870 255.085 ;
        RECT 94.850 254.900 95.470 255.085 ;
        RECT 63.250 254.670 95.470 254.900 ;
        RECT 63.250 254.485 63.870 254.670 ;
        RECT 94.850 254.485 95.470 254.670 ;
        RECT 95.700 254.900 96.320 255.085 ;
        RECT 127.300 254.900 127.920 255.085 ;
        RECT 95.700 254.670 127.920 254.900 ;
        RECT 95.700 254.485 96.320 254.670 ;
        RECT 127.300 254.485 127.920 254.670 ;
        RECT 128.150 254.900 128.770 255.085 ;
        RECT 159.750 254.900 160.370 255.085 ;
        RECT 128.150 254.670 160.370 254.900 ;
        RECT 128.150 254.485 128.770 254.670 ;
        RECT 159.750 254.485 160.370 254.670 ;
        RECT 43.040 254.405 44.660 254.415 ;
        RECT 75.490 254.405 77.110 254.415 ;
        RECT 107.940 254.405 109.560 254.415 ;
        RECT 140.390 254.405 142.010 254.415 ;
        RECT 31.650 254.035 62.170 254.405 ;
        RECT 64.100 254.035 94.620 254.405 ;
        RECT 96.550 254.035 127.070 254.405 ;
        RECT 129.000 254.035 159.520 254.405 ;
        RECT 31.660 253.240 62.160 253.680 ;
        RECT 64.110 253.240 94.610 253.680 ;
        RECT 96.560 253.240 127.060 253.680 ;
        RECT 129.010 253.240 159.510 253.680 ;
        RECT 31.650 252.510 62.170 252.890 ;
        RECT 64.100 252.510 94.620 252.890 ;
        RECT 96.550 252.510 127.070 252.890 ;
        RECT 129.000 252.510 159.520 252.890 ;
        RECT 30.800 252.255 31.420 252.440 ;
        RECT 62.400 252.255 63.020 252.440 ;
        RECT 30.800 252.025 63.020 252.255 ;
        RECT 30.800 251.840 31.420 252.025 ;
        RECT 62.400 251.840 63.020 252.025 ;
        RECT 63.250 252.255 63.870 252.440 ;
        RECT 94.850 252.255 95.470 252.440 ;
        RECT 63.250 252.025 95.470 252.255 ;
        RECT 63.250 251.840 63.870 252.025 ;
        RECT 94.850 251.840 95.470 252.025 ;
        RECT 95.700 252.255 96.320 252.440 ;
        RECT 127.300 252.255 127.920 252.440 ;
        RECT 95.700 252.025 127.920 252.255 ;
        RECT 95.700 251.840 96.320 252.025 ;
        RECT 127.300 251.840 127.920 252.025 ;
        RECT 128.150 252.255 128.770 252.440 ;
        RECT 159.750 252.255 160.370 252.440 ;
        RECT 128.150 252.025 160.370 252.255 ;
        RECT 128.150 251.840 128.770 252.025 ;
        RECT 159.750 251.840 160.370 252.025 ;
        RECT 39.200 251.760 40.820 251.770 ;
        RECT 71.650 251.760 73.270 251.770 ;
        RECT 104.100 251.760 105.720 251.770 ;
        RECT 136.550 251.760 138.170 251.770 ;
        RECT 31.650 251.390 62.170 251.760 ;
        RECT 64.100 251.390 94.620 251.760 ;
        RECT 96.550 251.390 127.070 251.760 ;
        RECT 129.000 251.390 159.520 251.760 ;
        RECT 31.650 250.670 62.170 251.050 ;
        RECT 64.100 250.670 94.620 251.050 ;
        RECT 96.550 250.670 127.070 251.050 ;
        RECT 129.000 250.670 159.520 251.050 ;
        RECT 30.800 250.415 31.420 250.600 ;
        RECT 62.400 250.415 63.020 250.600 ;
        RECT 30.800 250.185 63.020 250.415 ;
        RECT 30.800 250.000 31.420 250.185 ;
        RECT 62.400 250.000 63.020 250.185 ;
        RECT 63.250 250.415 63.870 250.600 ;
        RECT 94.850 250.415 95.470 250.600 ;
        RECT 63.250 250.185 95.470 250.415 ;
        RECT 63.250 250.000 63.870 250.185 ;
        RECT 94.850 250.000 95.470 250.185 ;
        RECT 95.700 250.415 96.320 250.600 ;
        RECT 127.300 250.415 127.920 250.600 ;
        RECT 95.700 250.185 127.920 250.415 ;
        RECT 95.700 250.000 96.320 250.185 ;
        RECT 127.300 250.000 127.920 250.185 ;
        RECT 128.150 250.415 128.770 250.600 ;
        RECT 159.750 250.415 160.370 250.600 ;
        RECT 128.150 250.185 160.370 250.415 ;
        RECT 128.150 250.000 128.770 250.185 ;
        RECT 159.750 250.000 160.370 250.185 ;
        RECT 35.360 249.920 36.980 249.930 ;
        RECT 67.810 249.920 69.430 249.930 ;
        RECT 100.260 249.920 101.880 249.930 ;
        RECT 132.710 249.920 134.330 249.930 ;
        RECT 31.650 249.550 62.170 249.920 ;
        RECT 64.100 249.550 94.620 249.920 ;
        RECT 96.550 249.550 127.070 249.920 ;
        RECT 129.000 249.550 159.520 249.920 ;
        RECT 31.650 248.830 62.170 249.210 ;
        RECT 64.100 248.830 94.620 249.210 ;
        RECT 96.550 248.830 127.070 249.210 ;
        RECT 129.000 248.830 159.520 249.210 ;
        RECT 30.800 248.575 31.420 248.760 ;
        RECT 62.400 248.575 63.020 248.760 ;
        RECT 30.800 248.345 63.020 248.575 ;
        RECT 30.800 248.160 31.420 248.345 ;
        RECT 62.400 248.160 63.020 248.345 ;
        RECT 63.250 248.575 63.870 248.760 ;
        RECT 94.850 248.575 95.470 248.760 ;
        RECT 63.250 248.345 95.470 248.575 ;
        RECT 63.250 248.160 63.870 248.345 ;
        RECT 94.850 248.160 95.470 248.345 ;
        RECT 95.700 248.575 96.320 248.760 ;
        RECT 127.300 248.575 127.920 248.760 ;
        RECT 95.700 248.345 127.920 248.575 ;
        RECT 95.700 248.160 96.320 248.345 ;
        RECT 127.300 248.160 127.920 248.345 ;
        RECT 128.150 248.575 128.770 248.760 ;
        RECT 159.750 248.575 160.370 248.760 ;
        RECT 128.150 248.345 160.370 248.575 ;
        RECT 128.150 248.160 128.770 248.345 ;
        RECT 159.750 248.160 160.370 248.345 ;
        RECT 31.650 247.710 62.170 248.080 ;
        RECT 64.100 247.710 94.620 248.080 ;
        RECT 96.550 247.710 127.070 248.080 ;
        RECT 129.000 247.710 159.520 248.080 ;
        RECT 25.090 245.360 27.380 245.700 ;
        RECT 28.125 245.360 29.610 245.700 ;
        RECT 25.090 244.725 25.690 245.360 ;
        RECT 25.090 244.495 26.670 244.725 ;
        RECT 25.090 242.455 25.690 244.495 ;
        RECT 27.100 244.265 27.460 244.350 ;
        RECT 25.970 244.035 27.460 244.265 ;
        RECT 25.970 243.885 26.330 244.035 ;
        RECT 25.920 243.250 26.870 243.655 ;
        RECT 25.090 242.225 26.380 242.455 ;
        RECT 25.090 241.265 25.690 242.225 ;
        RECT 26.610 241.905 26.870 243.250 ;
        RECT 27.100 242.600 27.460 244.035 ;
        RECT 27.690 242.700 28.040 243.900 ;
        RECT 28.400 243.290 28.780 244.935 ;
        RECT 27.480 241.905 27.830 241.965 ;
        RECT 28.400 241.905 28.740 242.510 ;
        RECT 26.610 241.645 28.740 241.905 ;
        RECT 27.480 241.585 27.830 241.645 ;
        RECT 29.010 241.365 29.610 245.360 ;
        RECT 31.455 244.925 33.205 247.710 ;
        RECT 33.845 244.925 34.655 245.925 ;
        RECT 35.295 244.925 37.045 247.220 ;
        RECT 37.685 244.925 38.495 245.925 ;
        RECT 39.135 244.925 40.885 247.220 ;
        RECT 41.525 244.925 42.335 245.925 ;
        RECT 42.975 244.925 44.725 247.220 ;
        RECT 45.365 244.925 46.175 245.925 ;
        RECT 46.815 244.925 48.565 247.220 ;
        RECT 49.205 244.925 50.015 245.925 ;
        RECT 50.655 244.925 52.405 247.220 ;
        RECT 53.045 244.925 53.855 245.925 ;
        RECT 54.495 244.925 56.245 247.220 ;
        RECT 56.885 244.925 57.695 245.925 ;
        RECT 58.335 244.925 60.085 247.220 ;
        RECT 60.725 244.925 61.535 245.925 ;
        RECT 63.905 244.925 65.655 247.710 ;
        RECT 66.295 244.925 67.105 245.925 ;
        RECT 67.745 244.925 69.495 247.220 ;
        RECT 70.135 244.925 70.945 245.925 ;
        RECT 71.585 244.925 73.335 247.220 ;
        RECT 73.975 244.925 74.785 245.925 ;
        RECT 75.425 244.925 77.175 247.220 ;
        RECT 77.815 244.925 78.625 245.925 ;
        RECT 79.265 244.925 81.015 247.220 ;
        RECT 81.655 244.925 82.465 245.925 ;
        RECT 83.105 244.925 84.855 247.220 ;
        RECT 85.495 244.925 86.305 245.925 ;
        RECT 86.945 244.925 88.695 247.220 ;
        RECT 89.335 244.925 90.145 245.925 ;
        RECT 90.785 244.925 92.535 247.220 ;
        RECT 93.175 244.925 93.985 245.925 ;
        RECT 96.355 244.925 98.105 247.710 ;
        RECT 98.745 244.925 99.555 245.925 ;
        RECT 100.195 244.925 101.945 247.220 ;
        RECT 102.585 244.925 103.395 245.925 ;
        RECT 104.035 244.925 105.785 247.220 ;
        RECT 106.425 244.925 107.235 245.925 ;
        RECT 107.875 244.925 109.625 247.220 ;
        RECT 110.265 244.925 111.075 245.925 ;
        RECT 111.715 244.925 113.465 247.220 ;
        RECT 114.105 244.925 114.915 245.925 ;
        RECT 115.555 244.925 117.305 247.220 ;
        RECT 117.945 244.925 118.755 245.925 ;
        RECT 119.395 244.925 121.145 247.220 ;
        RECT 121.785 244.925 122.595 245.925 ;
        RECT 123.235 244.925 124.985 247.220 ;
        RECT 125.625 244.925 126.435 245.925 ;
        RECT 128.805 244.925 130.555 247.710 ;
        RECT 131.195 244.925 132.005 245.925 ;
        RECT 132.645 244.925 134.395 247.220 ;
        RECT 135.035 244.925 135.845 245.925 ;
        RECT 136.485 244.925 138.235 247.220 ;
        RECT 138.875 244.925 139.685 245.925 ;
        RECT 140.325 244.925 142.075 247.220 ;
        RECT 142.715 244.925 143.525 245.925 ;
        RECT 144.165 244.925 145.915 247.220 ;
        RECT 146.555 244.925 147.365 245.925 ;
        RECT 148.005 244.925 149.755 247.220 ;
        RECT 150.395 244.925 151.205 245.925 ;
        RECT 151.845 244.925 153.595 247.220 ;
        RECT 154.235 244.925 155.045 245.925 ;
        RECT 155.685 244.925 157.435 247.220 ;
        RECT 158.075 244.925 158.885 245.925 ;
        RECT 161.300 245.115 161.670 263.625 ;
        RECT 162.320 259.990 162.690 263.625 ;
        RECT 162.315 259.610 162.695 259.990 ;
        RECT 162.320 256.990 162.690 259.610 ;
        RECT 162.315 256.610 162.695 256.990 ;
        RECT 162.320 253.990 162.690 256.610 ;
        RECT 162.315 253.610 162.695 253.990 ;
        RECT 162.320 250.990 162.690 253.610 ;
        RECT 162.315 250.610 162.695 250.990 ;
        RECT 162.320 247.990 162.690 250.610 ;
        RECT 162.315 247.610 162.695 247.990 ;
        RECT 161.300 244.735 161.680 245.115 ;
        RECT 161.300 243.665 161.670 244.735 ;
        RECT 31.925 242.475 32.735 243.475 ;
        RECT 25.090 241.035 26.780 241.265 ;
        RECT 28.150 241.135 29.610 241.365 ;
        RECT 25.090 239.025 25.690 241.035 ;
        RECT 27.110 240.575 28.110 240.900 ;
        RECT 25.920 240.015 28.780 240.345 ;
        RECT 25.090 238.795 26.780 239.025 ;
        RECT 25.090 236.785 25.690 238.795 ;
        RECT 27.495 238.660 27.760 240.015 ;
        RECT 29.010 239.125 29.610 241.135 ;
        RECT 33.375 240.645 35.125 243.475 ;
        RECT 35.765 242.475 36.575 243.475 ;
        RECT 37.215 241.180 38.965 243.475 ;
        RECT 39.605 242.475 40.415 243.475 ;
        RECT 41.055 241.180 42.805 243.475 ;
        RECT 43.445 242.475 44.255 243.475 ;
        RECT 44.895 241.180 46.645 243.475 ;
        RECT 47.285 242.475 48.095 243.475 ;
        RECT 48.735 241.180 50.485 243.475 ;
        RECT 51.125 242.475 51.935 243.475 ;
        RECT 52.575 241.180 54.325 243.475 ;
        RECT 54.965 242.475 55.775 243.475 ;
        RECT 56.415 241.180 58.165 243.475 ;
        RECT 58.805 242.475 59.615 243.475 ;
        RECT 60.255 241.180 62.005 243.475 ;
        RECT 64.375 242.475 65.185 243.475 ;
        RECT 65.825 240.645 67.575 243.475 ;
        RECT 68.215 242.475 69.025 243.475 ;
        RECT 69.665 241.180 71.415 243.475 ;
        RECT 72.055 242.475 72.865 243.475 ;
        RECT 73.505 241.180 75.255 243.475 ;
        RECT 75.895 242.475 76.705 243.475 ;
        RECT 77.345 241.180 79.095 243.475 ;
        RECT 79.735 242.475 80.545 243.475 ;
        RECT 81.185 241.180 82.935 243.475 ;
        RECT 83.575 242.475 84.385 243.475 ;
        RECT 85.025 241.180 86.775 243.475 ;
        RECT 87.415 242.475 88.225 243.475 ;
        RECT 88.865 241.180 90.615 243.475 ;
        RECT 91.255 242.475 92.065 243.475 ;
        RECT 92.705 241.180 94.455 243.475 ;
        RECT 96.825 242.475 97.635 243.475 ;
        RECT 98.275 240.645 100.025 243.475 ;
        RECT 100.665 242.475 101.475 243.475 ;
        RECT 102.115 241.180 103.865 243.475 ;
        RECT 104.505 242.475 105.315 243.475 ;
        RECT 105.955 241.180 107.705 243.475 ;
        RECT 108.345 242.475 109.155 243.475 ;
        RECT 109.795 241.180 111.545 243.475 ;
        RECT 112.185 242.475 112.995 243.475 ;
        RECT 113.635 241.180 115.385 243.475 ;
        RECT 116.025 242.475 116.835 243.475 ;
        RECT 117.475 241.180 119.225 243.475 ;
        RECT 119.865 242.475 120.675 243.475 ;
        RECT 121.315 241.180 123.065 243.475 ;
        RECT 123.705 242.475 124.515 243.475 ;
        RECT 125.155 241.180 126.905 243.475 ;
        RECT 129.275 242.475 130.085 243.475 ;
        RECT 130.725 240.645 132.475 243.475 ;
        RECT 133.115 242.475 133.925 243.475 ;
        RECT 134.565 241.180 136.315 243.475 ;
        RECT 136.955 242.475 137.765 243.475 ;
        RECT 138.405 241.180 140.155 243.475 ;
        RECT 140.795 242.475 141.605 243.475 ;
        RECT 142.245 241.180 143.995 243.475 ;
        RECT 144.635 242.475 145.445 243.475 ;
        RECT 146.085 241.180 147.835 243.475 ;
        RECT 148.475 242.475 149.285 243.475 ;
        RECT 149.925 241.180 151.675 243.475 ;
        RECT 152.315 242.475 153.125 243.475 ;
        RECT 153.765 241.180 155.515 243.475 ;
        RECT 156.155 242.475 156.965 243.475 ;
        RECT 157.605 241.180 159.355 243.475 ;
        RECT 161.300 243.285 161.680 243.665 ;
        RECT 31.650 240.275 62.170 240.645 ;
        RECT 64.100 240.275 94.620 240.645 ;
        RECT 96.550 240.275 127.070 240.645 ;
        RECT 129.000 240.275 159.520 240.645 ;
        RECT 30.800 240.010 31.420 240.195 ;
        RECT 62.400 240.010 63.020 240.195 ;
        RECT 30.800 239.780 63.020 240.010 ;
        RECT 30.800 239.595 31.420 239.780 ;
        RECT 62.400 239.595 63.020 239.780 ;
        RECT 63.250 240.010 63.870 240.195 ;
        RECT 94.850 240.010 95.470 240.195 ;
        RECT 63.250 239.780 95.470 240.010 ;
        RECT 63.250 239.595 63.870 239.780 ;
        RECT 94.850 239.595 95.470 239.780 ;
        RECT 95.700 240.010 96.320 240.195 ;
        RECT 127.300 240.010 127.920 240.195 ;
        RECT 95.700 239.780 127.920 240.010 ;
        RECT 95.700 239.595 96.320 239.780 ;
        RECT 127.300 239.595 127.920 239.780 ;
        RECT 128.150 240.010 128.770 240.195 ;
        RECT 159.750 240.010 160.370 240.195 ;
        RECT 128.150 239.780 160.370 240.010 ;
        RECT 128.150 239.595 128.770 239.780 ;
        RECT 159.750 239.595 160.370 239.780 ;
        RECT 31.650 239.145 62.170 239.525 ;
        RECT 64.100 239.145 94.620 239.525 ;
        RECT 96.550 239.145 127.070 239.525 ;
        RECT 129.000 239.145 159.520 239.525 ;
        RECT 28.150 238.895 29.610 239.125 ;
        RECT 27.110 238.335 28.110 238.660 ;
        RECT 25.920 237.775 28.780 238.105 ;
        RECT 29.010 236.885 29.610 238.895 ;
        RECT 31.650 238.435 62.170 238.805 ;
        RECT 64.100 238.435 94.620 238.805 ;
        RECT 96.550 238.435 127.070 238.805 ;
        RECT 129.000 238.435 159.520 238.805 ;
        RECT 37.280 238.425 38.900 238.435 ;
        RECT 69.730 238.425 71.350 238.435 ;
        RECT 102.180 238.425 103.800 238.435 ;
        RECT 134.630 238.425 136.250 238.435 ;
        RECT 30.800 238.170 31.420 238.355 ;
        RECT 62.400 238.170 63.020 238.355 ;
        RECT 30.800 237.940 63.020 238.170 ;
        RECT 30.800 237.755 31.420 237.940 ;
        RECT 62.400 237.755 63.020 237.940 ;
        RECT 63.250 238.170 63.870 238.355 ;
        RECT 94.850 238.170 95.470 238.355 ;
        RECT 63.250 237.940 95.470 238.170 ;
        RECT 63.250 237.755 63.870 237.940 ;
        RECT 94.850 237.755 95.470 237.940 ;
        RECT 95.700 238.170 96.320 238.355 ;
        RECT 127.300 238.170 127.920 238.355 ;
        RECT 95.700 237.940 127.920 238.170 ;
        RECT 95.700 237.755 96.320 237.940 ;
        RECT 127.300 237.755 127.920 237.940 ;
        RECT 128.150 238.170 128.770 238.355 ;
        RECT 159.750 238.170 160.370 238.355 ;
        RECT 128.150 237.940 160.370 238.170 ;
        RECT 128.150 237.755 128.770 237.940 ;
        RECT 159.750 237.755 160.370 237.940 ;
        RECT 31.650 237.305 62.170 237.685 ;
        RECT 64.100 237.305 94.620 237.685 ;
        RECT 96.550 237.305 127.070 237.685 ;
        RECT 129.000 237.305 159.520 237.685 ;
        RECT 25.090 236.555 26.780 236.785 ;
        RECT 28.150 236.655 29.610 236.885 ;
        RECT 25.090 234.500 25.690 236.555 ;
        RECT 27.110 236.095 28.110 236.420 ;
        RECT 29.010 234.500 29.610 236.655 ;
        RECT 31.650 236.590 62.170 236.960 ;
        RECT 64.100 236.590 94.620 236.960 ;
        RECT 96.550 236.590 127.070 236.960 ;
        RECT 129.000 236.590 159.520 236.960 ;
        RECT 41.120 236.580 42.740 236.590 ;
        RECT 73.570 236.580 75.190 236.590 ;
        RECT 106.020 236.580 107.640 236.590 ;
        RECT 138.470 236.580 140.090 236.590 ;
        RECT 30.800 236.325 31.420 236.510 ;
        RECT 62.400 236.325 63.020 236.510 ;
        RECT 30.800 236.095 63.020 236.325 ;
        RECT 30.800 235.910 31.420 236.095 ;
        RECT 62.400 235.910 63.020 236.095 ;
        RECT 63.250 236.325 63.870 236.510 ;
        RECT 94.850 236.325 95.470 236.510 ;
        RECT 63.250 236.095 95.470 236.325 ;
        RECT 63.250 235.910 63.870 236.095 ;
        RECT 94.850 235.910 95.470 236.095 ;
        RECT 95.700 236.325 96.320 236.510 ;
        RECT 127.300 236.325 127.920 236.510 ;
        RECT 95.700 236.095 127.920 236.325 ;
        RECT 95.700 235.910 96.320 236.095 ;
        RECT 127.300 235.910 127.920 236.095 ;
        RECT 128.150 236.325 128.770 236.510 ;
        RECT 159.750 236.325 160.370 236.510 ;
        RECT 128.150 236.095 160.370 236.325 ;
        RECT 128.150 235.910 128.770 236.095 ;
        RECT 159.750 235.910 160.370 236.095 ;
        RECT 31.650 235.460 62.170 235.840 ;
        RECT 64.100 235.460 94.620 235.840 ;
        RECT 96.550 235.460 127.070 235.840 ;
        RECT 129.000 235.460 159.520 235.840 ;
        RECT 31.660 234.670 62.160 235.110 ;
        RECT 64.110 234.670 94.610 235.110 ;
        RECT 96.560 234.670 127.060 235.110 ;
        RECT 129.010 234.670 159.510 235.110 ;
        RECT 25.090 234.160 27.380 234.500 ;
        RECT 28.125 234.160 29.610 234.500 ;
        RECT 25.090 206.315 25.690 234.160 ;
        RECT 29.010 206.315 29.610 234.160 ;
        RECT 31.650 233.950 62.170 234.320 ;
        RECT 64.100 233.950 94.620 234.320 ;
        RECT 96.550 233.950 127.070 234.320 ;
        RECT 129.000 233.950 159.520 234.320 ;
        RECT 44.960 233.940 46.580 233.950 ;
        RECT 77.410 233.940 79.030 233.950 ;
        RECT 109.860 233.940 111.480 233.950 ;
        RECT 142.310 233.940 143.930 233.950 ;
        RECT 30.800 233.685 31.420 233.870 ;
        RECT 62.400 233.685 63.020 233.870 ;
        RECT 30.800 233.455 63.020 233.685 ;
        RECT 30.800 233.270 31.420 233.455 ;
        RECT 62.400 233.270 63.020 233.455 ;
        RECT 63.250 233.685 63.870 233.870 ;
        RECT 94.850 233.685 95.470 233.870 ;
        RECT 63.250 233.455 95.470 233.685 ;
        RECT 63.250 233.270 63.870 233.455 ;
        RECT 94.850 233.270 95.470 233.455 ;
        RECT 95.700 233.685 96.320 233.870 ;
        RECT 127.300 233.685 127.920 233.870 ;
        RECT 95.700 233.455 127.920 233.685 ;
        RECT 95.700 233.270 96.320 233.455 ;
        RECT 127.300 233.270 127.920 233.455 ;
        RECT 128.150 233.685 128.770 233.870 ;
        RECT 159.750 233.685 160.370 233.870 ;
        RECT 128.150 233.455 160.370 233.685 ;
        RECT 128.150 233.270 128.770 233.455 ;
        RECT 159.750 233.270 160.370 233.455 ;
        RECT 31.650 232.820 62.170 233.200 ;
        RECT 64.100 232.820 94.620 233.200 ;
        RECT 96.550 232.820 127.070 233.200 ;
        RECT 129.000 232.820 159.520 233.200 ;
        RECT 31.650 232.110 62.170 232.480 ;
        RECT 64.100 232.110 94.620 232.480 ;
        RECT 96.550 232.110 127.070 232.480 ;
        RECT 129.000 232.110 159.520 232.480 ;
        RECT 48.800 232.100 50.420 232.110 ;
        RECT 81.250 232.100 82.870 232.110 ;
        RECT 113.700 232.100 115.320 232.110 ;
        RECT 146.150 232.100 147.770 232.110 ;
        RECT 30.800 231.845 31.420 232.030 ;
        RECT 62.400 231.845 63.020 232.030 ;
        RECT 30.800 231.615 63.020 231.845 ;
        RECT 30.800 231.430 31.420 231.615 ;
        RECT 62.400 231.430 63.020 231.615 ;
        RECT 63.250 231.845 63.870 232.030 ;
        RECT 94.850 231.845 95.470 232.030 ;
        RECT 63.250 231.615 95.470 231.845 ;
        RECT 63.250 231.430 63.870 231.615 ;
        RECT 94.850 231.430 95.470 231.615 ;
        RECT 95.700 231.845 96.320 232.030 ;
        RECT 127.300 231.845 127.920 232.030 ;
        RECT 95.700 231.615 127.920 231.845 ;
        RECT 95.700 231.430 96.320 231.615 ;
        RECT 127.300 231.430 127.920 231.615 ;
        RECT 128.150 231.845 128.770 232.030 ;
        RECT 159.750 231.845 160.370 232.030 ;
        RECT 128.150 231.615 160.370 231.845 ;
        RECT 128.150 231.430 128.770 231.615 ;
        RECT 159.750 231.430 160.370 231.615 ;
        RECT 31.650 230.980 62.170 231.360 ;
        RECT 64.100 230.980 94.620 231.360 ;
        RECT 96.550 230.980 127.070 231.360 ;
        RECT 129.000 230.980 159.520 231.360 ;
        RECT 31.650 230.265 62.170 230.635 ;
        RECT 64.100 230.265 94.620 230.635 ;
        RECT 96.550 230.265 127.070 230.635 ;
        RECT 129.000 230.265 159.520 230.635 ;
        RECT 52.640 230.255 54.260 230.265 ;
        RECT 85.090 230.255 86.710 230.265 ;
        RECT 117.540 230.255 119.160 230.265 ;
        RECT 149.990 230.255 151.610 230.265 ;
        RECT 30.800 230.000 31.420 230.185 ;
        RECT 62.400 230.000 63.020 230.185 ;
        RECT 30.800 229.770 63.020 230.000 ;
        RECT 30.800 229.585 31.420 229.770 ;
        RECT 62.400 229.585 63.020 229.770 ;
        RECT 63.250 230.000 63.870 230.185 ;
        RECT 94.850 230.000 95.470 230.185 ;
        RECT 63.250 229.770 95.470 230.000 ;
        RECT 63.250 229.585 63.870 229.770 ;
        RECT 94.850 229.585 95.470 229.770 ;
        RECT 95.700 230.000 96.320 230.185 ;
        RECT 127.300 230.000 127.920 230.185 ;
        RECT 95.700 229.770 127.920 230.000 ;
        RECT 95.700 229.585 96.320 229.770 ;
        RECT 127.300 229.585 127.920 229.770 ;
        RECT 128.150 230.000 128.770 230.185 ;
        RECT 159.750 230.000 160.370 230.185 ;
        RECT 128.150 229.770 160.370 230.000 ;
        RECT 128.150 229.585 128.770 229.770 ;
        RECT 159.750 229.585 160.370 229.770 ;
        RECT 31.650 229.135 62.170 229.515 ;
        RECT 64.100 229.135 94.620 229.515 ;
        RECT 96.550 229.135 127.070 229.515 ;
        RECT 129.000 229.135 159.520 229.515 ;
        RECT 31.660 228.345 62.160 228.785 ;
        RECT 64.110 228.345 94.610 228.785 ;
        RECT 96.560 228.345 127.060 228.785 ;
        RECT 129.010 228.345 159.510 228.785 ;
        RECT 31.650 227.625 62.170 227.995 ;
        RECT 64.100 227.625 94.620 227.995 ;
        RECT 96.550 227.625 127.070 227.995 ;
        RECT 129.000 227.625 159.520 227.995 ;
        RECT 56.480 227.615 58.100 227.625 ;
        RECT 88.930 227.615 90.550 227.625 ;
        RECT 121.380 227.615 123.000 227.625 ;
        RECT 153.830 227.615 155.450 227.625 ;
        RECT 30.800 227.360 31.420 227.545 ;
        RECT 62.400 227.360 63.020 227.545 ;
        RECT 30.800 227.130 63.020 227.360 ;
        RECT 30.800 226.945 31.420 227.130 ;
        RECT 62.400 226.945 63.020 227.130 ;
        RECT 63.250 227.360 63.870 227.545 ;
        RECT 94.850 227.360 95.470 227.545 ;
        RECT 63.250 227.130 95.470 227.360 ;
        RECT 63.250 226.945 63.870 227.130 ;
        RECT 94.850 226.945 95.470 227.130 ;
        RECT 95.700 227.360 96.320 227.545 ;
        RECT 127.300 227.360 127.920 227.545 ;
        RECT 95.700 227.130 127.920 227.360 ;
        RECT 95.700 226.945 96.320 227.130 ;
        RECT 127.300 226.945 127.920 227.130 ;
        RECT 128.150 227.360 128.770 227.545 ;
        RECT 159.750 227.360 160.370 227.545 ;
        RECT 128.150 227.130 160.370 227.360 ;
        RECT 128.150 226.945 128.770 227.130 ;
        RECT 159.750 226.945 160.370 227.130 ;
        RECT 31.650 226.495 62.170 226.875 ;
        RECT 64.100 226.495 94.620 226.875 ;
        RECT 96.550 226.495 127.070 226.875 ;
        RECT 129.000 226.495 159.520 226.875 ;
        RECT 31.650 225.785 62.170 226.155 ;
        RECT 64.100 225.785 94.620 226.155 ;
        RECT 96.550 225.785 127.070 226.155 ;
        RECT 129.000 225.785 159.520 226.155 ;
        RECT 60.320 225.775 61.940 225.785 ;
        RECT 92.770 225.775 94.390 225.785 ;
        RECT 125.220 225.775 126.840 225.785 ;
        RECT 157.670 225.775 159.290 225.785 ;
        RECT 30.800 225.520 31.420 225.705 ;
        RECT 62.400 225.520 63.020 225.705 ;
        RECT 30.800 225.290 63.020 225.520 ;
        RECT 30.800 225.105 31.420 225.290 ;
        RECT 62.400 225.105 63.020 225.290 ;
        RECT 63.250 225.520 63.870 225.705 ;
        RECT 94.850 225.520 95.470 225.705 ;
        RECT 63.250 225.290 95.470 225.520 ;
        RECT 63.250 225.105 63.870 225.290 ;
        RECT 94.850 225.105 95.470 225.290 ;
        RECT 95.700 225.520 96.320 225.705 ;
        RECT 127.300 225.520 127.920 225.705 ;
        RECT 95.700 225.290 127.920 225.520 ;
        RECT 95.700 225.105 96.320 225.290 ;
        RECT 127.300 225.105 127.920 225.290 ;
        RECT 128.150 225.520 128.770 225.705 ;
        RECT 159.750 225.520 160.370 225.705 ;
        RECT 128.150 225.290 160.370 225.520 ;
        RECT 161.300 225.355 161.670 243.285 ;
        RECT 162.320 241.990 162.690 247.610 ;
        RECT 163.340 245.115 163.710 263.625 ;
        RECT 164.360 259.990 164.730 263.625 ;
        RECT 164.355 259.610 164.735 259.990 ;
        RECT 164.360 256.990 164.730 259.610 ;
        RECT 164.355 256.610 164.735 256.990 ;
        RECT 164.360 253.990 164.730 256.610 ;
        RECT 164.355 253.610 164.735 253.990 ;
        RECT 164.360 250.990 164.730 253.610 ;
        RECT 164.355 250.610 164.735 250.990 ;
        RECT 164.360 247.990 164.730 250.610 ;
        RECT 164.355 247.610 164.735 247.990 ;
        RECT 163.340 244.735 163.720 245.115 ;
        RECT 163.340 243.665 163.710 244.735 ;
        RECT 163.340 243.285 163.720 243.665 ;
        RECT 162.315 241.610 162.695 241.990 ;
        RECT 162.320 238.990 162.690 241.610 ;
        RECT 162.315 238.610 162.695 238.990 ;
        RECT 162.320 235.990 162.690 238.610 ;
        RECT 162.315 235.610 162.695 235.990 ;
        RECT 162.320 232.990 162.690 235.610 ;
        RECT 162.315 232.610 162.695 232.990 ;
        RECT 162.320 229.990 162.690 232.610 ;
        RECT 162.315 229.610 162.695 229.990 ;
        RECT 162.320 226.990 162.690 229.610 ;
        RECT 162.315 226.610 162.695 226.990 ;
        RECT 162.320 225.355 162.690 226.610 ;
        RECT 163.340 225.355 163.710 243.285 ;
        RECT 164.360 241.990 164.730 247.610 ;
        RECT 164.355 241.610 164.735 241.990 ;
        RECT 164.360 238.990 164.730 241.610 ;
        RECT 164.355 238.610 164.735 238.990 ;
        RECT 164.360 235.990 164.730 238.610 ;
        RECT 164.355 235.610 164.735 235.990 ;
        RECT 164.360 232.990 164.730 235.610 ;
        RECT 164.355 232.610 164.735 232.990 ;
        RECT 164.360 229.990 164.730 232.610 ;
        RECT 164.355 229.610 164.735 229.990 ;
        RECT 164.360 226.990 164.730 229.610 ;
        RECT 164.355 226.610 164.735 226.990 ;
        RECT 164.360 225.355 164.730 226.610 ;
        RECT 165.380 225.355 165.760 263.625 ;
        RECT 166.110 225.365 166.550 263.615 ;
        RECT 128.150 225.105 128.770 225.290 ;
        RECT 159.750 225.105 160.370 225.290 ;
        RECT 31.650 224.655 62.170 225.035 ;
        RECT 64.100 224.655 94.620 225.035 ;
        RECT 96.550 224.655 127.070 225.035 ;
        RECT 129.000 224.655 159.520 225.035 ;
        RECT 31.650 223.935 62.170 224.315 ;
        RECT 64.100 223.935 94.620 224.315 ;
        RECT 96.550 223.935 127.070 224.315 ;
        RECT 129.000 223.935 159.520 224.315 ;
        RECT 30.800 223.680 31.420 223.865 ;
        RECT 62.400 223.680 63.020 223.865 ;
        RECT 30.800 223.450 63.020 223.680 ;
        RECT 30.800 223.265 31.420 223.450 ;
        RECT 62.400 223.265 63.020 223.450 ;
        RECT 63.250 223.680 63.870 223.865 ;
        RECT 94.850 223.680 95.470 223.865 ;
        RECT 63.250 223.450 95.470 223.680 ;
        RECT 63.250 223.265 63.870 223.450 ;
        RECT 94.850 223.265 95.470 223.450 ;
        RECT 95.700 223.680 96.320 223.865 ;
        RECT 127.300 223.680 127.920 223.865 ;
        RECT 95.700 223.450 127.920 223.680 ;
        RECT 95.700 223.265 96.320 223.450 ;
        RECT 127.300 223.265 127.920 223.450 ;
        RECT 128.150 223.680 128.770 223.865 ;
        RECT 159.750 223.680 160.370 223.865 ;
        RECT 128.150 223.450 160.370 223.680 ;
        RECT 128.150 223.265 128.770 223.450 ;
        RECT 159.750 223.265 160.370 223.450 ;
        RECT 58.400 223.185 60.020 223.195 ;
        RECT 90.850 223.185 92.470 223.195 ;
        RECT 123.300 223.185 124.920 223.195 ;
        RECT 155.750 223.185 157.370 223.195 ;
        RECT 31.650 222.815 62.170 223.185 ;
        RECT 64.100 222.815 94.620 223.185 ;
        RECT 96.550 222.815 127.070 223.185 ;
        RECT 129.000 222.815 159.520 223.185 ;
        RECT 31.650 222.095 62.170 222.475 ;
        RECT 64.100 222.095 94.620 222.475 ;
        RECT 96.550 222.095 127.070 222.475 ;
        RECT 129.000 222.095 159.520 222.475 ;
        RECT 30.800 221.840 31.420 222.025 ;
        RECT 62.400 221.840 63.020 222.025 ;
        RECT 30.800 221.610 63.020 221.840 ;
        RECT 30.800 221.425 31.420 221.610 ;
        RECT 62.400 221.425 63.020 221.610 ;
        RECT 63.250 221.840 63.870 222.025 ;
        RECT 94.850 221.840 95.470 222.025 ;
        RECT 63.250 221.610 95.470 221.840 ;
        RECT 63.250 221.425 63.870 221.610 ;
        RECT 94.850 221.425 95.470 221.610 ;
        RECT 95.700 221.840 96.320 222.025 ;
        RECT 127.300 221.840 127.920 222.025 ;
        RECT 95.700 221.610 127.920 221.840 ;
        RECT 95.700 221.425 96.320 221.610 ;
        RECT 127.300 221.425 127.920 221.610 ;
        RECT 128.150 221.840 128.770 222.025 ;
        RECT 159.750 221.840 160.370 222.025 ;
        RECT 128.150 221.610 160.370 221.840 ;
        RECT 128.150 221.425 128.770 221.610 ;
        RECT 159.750 221.425 160.370 221.610 ;
        RECT 54.560 221.345 56.180 221.355 ;
        RECT 87.010 221.345 88.630 221.355 ;
        RECT 119.460 221.345 121.080 221.355 ;
        RECT 151.910 221.345 153.530 221.355 ;
        RECT 31.650 220.975 62.170 221.345 ;
        RECT 64.100 220.975 94.620 221.345 ;
        RECT 96.550 220.975 127.070 221.345 ;
        RECT 129.000 220.975 159.520 221.345 ;
        RECT 31.660 220.180 62.160 220.620 ;
        RECT 64.110 220.180 94.610 220.620 ;
        RECT 96.560 220.180 127.060 220.620 ;
        RECT 129.010 220.180 159.510 220.620 ;
        RECT 31.650 219.450 62.170 219.830 ;
        RECT 64.100 219.450 94.620 219.830 ;
        RECT 96.550 219.450 127.070 219.830 ;
        RECT 129.000 219.450 159.520 219.830 ;
        RECT 30.800 219.195 31.420 219.380 ;
        RECT 62.400 219.195 63.020 219.380 ;
        RECT 30.800 218.965 63.020 219.195 ;
        RECT 30.800 218.780 31.420 218.965 ;
        RECT 62.400 218.780 63.020 218.965 ;
        RECT 63.250 219.195 63.870 219.380 ;
        RECT 94.850 219.195 95.470 219.380 ;
        RECT 63.250 218.965 95.470 219.195 ;
        RECT 63.250 218.780 63.870 218.965 ;
        RECT 94.850 218.780 95.470 218.965 ;
        RECT 95.700 219.195 96.320 219.380 ;
        RECT 127.300 219.195 127.920 219.380 ;
        RECT 95.700 218.965 127.920 219.195 ;
        RECT 95.700 218.780 96.320 218.965 ;
        RECT 127.300 218.780 127.920 218.965 ;
        RECT 128.150 219.195 128.770 219.380 ;
        RECT 159.750 219.195 160.370 219.380 ;
        RECT 128.150 218.965 160.370 219.195 ;
        RECT 128.150 218.780 128.770 218.965 ;
        RECT 159.750 218.780 160.370 218.965 ;
        RECT 50.720 218.700 52.340 218.710 ;
        RECT 83.170 218.700 84.790 218.710 ;
        RECT 115.620 218.700 117.240 218.710 ;
        RECT 148.070 218.700 149.690 218.710 ;
        RECT 31.650 218.330 62.170 218.700 ;
        RECT 64.100 218.330 94.620 218.700 ;
        RECT 96.550 218.330 127.070 218.700 ;
        RECT 129.000 218.330 159.520 218.700 ;
        RECT 31.650 217.610 62.170 217.990 ;
        RECT 64.100 217.610 94.620 217.990 ;
        RECT 96.550 217.610 127.070 217.990 ;
        RECT 129.000 217.610 159.520 217.990 ;
        RECT 30.800 217.355 31.420 217.540 ;
        RECT 62.400 217.355 63.020 217.540 ;
        RECT 30.800 217.125 63.020 217.355 ;
        RECT 30.800 216.940 31.420 217.125 ;
        RECT 62.400 216.940 63.020 217.125 ;
        RECT 63.250 217.355 63.870 217.540 ;
        RECT 94.850 217.355 95.470 217.540 ;
        RECT 63.250 217.125 95.470 217.355 ;
        RECT 63.250 216.940 63.870 217.125 ;
        RECT 94.850 216.940 95.470 217.125 ;
        RECT 95.700 217.355 96.320 217.540 ;
        RECT 127.300 217.355 127.920 217.540 ;
        RECT 95.700 217.125 127.920 217.355 ;
        RECT 95.700 216.940 96.320 217.125 ;
        RECT 127.300 216.940 127.920 217.125 ;
        RECT 128.150 217.355 128.770 217.540 ;
        RECT 159.750 217.355 160.370 217.540 ;
        RECT 128.150 217.125 160.370 217.355 ;
        RECT 128.150 216.940 128.770 217.125 ;
        RECT 159.750 216.940 160.370 217.125 ;
        RECT 46.880 216.860 48.500 216.870 ;
        RECT 79.330 216.860 80.950 216.870 ;
        RECT 111.780 216.860 113.400 216.870 ;
        RECT 144.230 216.860 145.850 216.870 ;
        RECT 31.650 216.490 62.170 216.860 ;
        RECT 64.100 216.490 94.620 216.860 ;
        RECT 96.550 216.490 127.070 216.860 ;
        RECT 129.000 216.490 159.520 216.860 ;
        RECT 31.650 215.770 62.170 216.150 ;
        RECT 64.100 215.770 94.620 216.150 ;
        RECT 96.550 215.770 127.070 216.150 ;
        RECT 129.000 215.770 159.520 216.150 ;
        RECT 30.800 215.515 31.420 215.700 ;
        RECT 62.400 215.515 63.020 215.700 ;
        RECT 30.800 215.285 63.020 215.515 ;
        RECT 30.800 215.100 31.420 215.285 ;
        RECT 62.400 215.100 63.020 215.285 ;
        RECT 63.250 215.515 63.870 215.700 ;
        RECT 94.850 215.515 95.470 215.700 ;
        RECT 63.250 215.285 95.470 215.515 ;
        RECT 63.250 215.100 63.870 215.285 ;
        RECT 94.850 215.100 95.470 215.285 ;
        RECT 95.700 215.515 96.320 215.700 ;
        RECT 127.300 215.515 127.920 215.700 ;
        RECT 95.700 215.285 127.920 215.515 ;
        RECT 95.700 215.100 96.320 215.285 ;
        RECT 127.300 215.100 127.920 215.285 ;
        RECT 128.150 215.515 128.770 215.700 ;
        RECT 159.750 215.515 160.370 215.700 ;
        RECT 128.150 215.285 160.370 215.515 ;
        RECT 128.150 215.100 128.770 215.285 ;
        RECT 159.750 215.100 160.370 215.285 ;
        RECT 43.040 215.020 44.660 215.030 ;
        RECT 75.490 215.020 77.110 215.030 ;
        RECT 107.940 215.020 109.560 215.030 ;
        RECT 140.390 215.020 142.010 215.030 ;
        RECT 31.650 214.650 62.170 215.020 ;
        RECT 64.100 214.650 94.620 215.020 ;
        RECT 96.550 214.650 127.070 215.020 ;
        RECT 129.000 214.650 159.520 215.020 ;
        RECT 31.660 213.855 62.160 214.295 ;
        RECT 64.110 213.855 94.610 214.295 ;
        RECT 96.560 213.855 127.060 214.295 ;
        RECT 129.010 213.855 159.510 214.295 ;
        RECT 31.650 213.125 62.170 213.505 ;
        RECT 64.100 213.125 94.620 213.505 ;
        RECT 96.550 213.125 127.070 213.505 ;
        RECT 129.000 213.125 159.520 213.505 ;
        RECT 30.800 212.870 31.420 213.055 ;
        RECT 62.400 212.870 63.020 213.055 ;
        RECT 30.800 212.640 63.020 212.870 ;
        RECT 30.800 212.455 31.420 212.640 ;
        RECT 62.400 212.455 63.020 212.640 ;
        RECT 63.250 212.870 63.870 213.055 ;
        RECT 94.850 212.870 95.470 213.055 ;
        RECT 63.250 212.640 95.470 212.870 ;
        RECT 63.250 212.455 63.870 212.640 ;
        RECT 94.850 212.455 95.470 212.640 ;
        RECT 95.700 212.870 96.320 213.055 ;
        RECT 127.300 212.870 127.920 213.055 ;
        RECT 95.700 212.640 127.920 212.870 ;
        RECT 95.700 212.455 96.320 212.640 ;
        RECT 127.300 212.455 127.920 212.640 ;
        RECT 128.150 212.870 128.770 213.055 ;
        RECT 159.750 212.870 160.370 213.055 ;
        RECT 128.150 212.640 160.370 212.870 ;
        RECT 128.150 212.455 128.770 212.640 ;
        RECT 159.750 212.455 160.370 212.640 ;
        RECT 39.200 212.375 40.820 212.385 ;
        RECT 71.650 212.375 73.270 212.385 ;
        RECT 104.100 212.375 105.720 212.385 ;
        RECT 136.550 212.375 138.170 212.385 ;
        RECT 31.650 212.005 62.170 212.375 ;
        RECT 64.100 212.005 94.620 212.375 ;
        RECT 96.550 212.005 127.070 212.375 ;
        RECT 129.000 212.005 159.520 212.375 ;
        RECT 31.650 211.285 62.170 211.665 ;
        RECT 64.100 211.285 94.620 211.665 ;
        RECT 96.550 211.285 127.070 211.665 ;
        RECT 129.000 211.285 159.520 211.665 ;
        RECT 30.800 211.030 31.420 211.215 ;
        RECT 62.400 211.030 63.020 211.215 ;
        RECT 30.800 210.800 63.020 211.030 ;
        RECT 30.800 210.615 31.420 210.800 ;
        RECT 62.400 210.615 63.020 210.800 ;
        RECT 63.250 211.030 63.870 211.215 ;
        RECT 94.850 211.030 95.470 211.215 ;
        RECT 63.250 210.800 95.470 211.030 ;
        RECT 63.250 210.615 63.870 210.800 ;
        RECT 94.850 210.615 95.470 210.800 ;
        RECT 95.700 211.030 96.320 211.215 ;
        RECT 127.300 211.030 127.920 211.215 ;
        RECT 95.700 210.800 127.920 211.030 ;
        RECT 95.700 210.615 96.320 210.800 ;
        RECT 127.300 210.615 127.920 210.800 ;
        RECT 128.150 211.030 128.770 211.215 ;
        RECT 159.750 211.030 160.370 211.215 ;
        RECT 128.150 210.800 160.370 211.030 ;
        RECT 128.150 210.615 128.770 210.800 ;
        RECT 159.750 210.615 160.370 210.800 ;
        RECT 35.360 210.535 36.980 210.545 ;
        RECT 67.810 210.535 69.430 210.545 ;
        RECT 100.260 210.535 101.880 210.545 ;
        RECT 132.710 210.535 134.330 210.545 ;
        RECT 31.650 210.165 62.170 210.535 ;
        RECT 64.100 210.165 94.620 210.535 ;
        RECT 96.550 210.165 127.070 210.535 ;
        RECT 129.000 210.165 159.520 210.535 ;
        RECT 31.650 209.445 62.170 209.825 ;
        RECT 64.100 209.445 94.620 209.825 ;
        RECT 96.550 209.445 127.070 209.825 ;
        RECT 129.000 209.445 159.520 209.825 ;
        RECT 30.800 209.190 31.420 209.375 ;
        RECT 62.400 209.190 63.020 209.375 ;
        RECT 30.800 208.960 63.020 209.190 ;
        RECT 30.800 208.775 31.420 208.960 ;
        RECT 62.400 208.775 63.020 208.960 ;
        RECT 63.250 209.190 63.870 209.375 ;
        RECT 94.850 209.190 95.470 209.375 ;
        RECT 63.250 208.960 95.470 209.190 ;
        RECT 63.250 208.775 63.870 208.960 ;
        RECT 94.850 208.775 95.470 208.960 ;
        RECT 95.700 209.190 96.320 209.375 ;
        RECT 127.300 209.190 127.920 209.375 ;
        RECT 95.700 208.960 127.920 209.190 ;
        RECT 95.700 208.775 96.320 208.960 ;
        RECT 127.300 208.775 127.920 208.960 ;
        RECT 128.150 209.190 128.770 209.375 ;
        RECT 159.750 209.190 160.370 209.375 ;
        RECT 128.150 208.960 160.370 209.190 ;
        RECT 128.150 208.775 128.770 208.960 ;
        RECT 159.750 208.775 160.370 208.960 ;
        RECT 31.650 208.325 62.170 208.695 ;
        RECT 64.100 208.325 94.620 208.695 ;
        RECT 96.550 208.325 127.070 208.695 ;
        RECT 129.000 208.325 159.520 208.695 ;
        RECT 25.090 205.975 27.380 206.315 ;
        RECT 28.125 205.975 29.610 206.315 ;
        RECT 25.090 205.340 25.690 205.975 ;
        RECT 25.090 205.110 26.670 205.340 ;
        RECT 25.090 203.070 25.690 205.110 ;
        RECT 27.100 204.880 27.460 204.965 ;
        RECT 25.970 204.650 27.460 204.880 ;
        RECT 25.970 204.500 26.330 204.650 ;
        RECT 25.920 203.865 26.870 204.270 ;
        RECT 25.090 202.840 26.380 203.070 ;
        RECT 25.090 201.880 25.690 202.840 ;
        RECT 26.610 202.520 26.870 203.865 ;
        RECT 27.100 203.215 27.460 204.650 ;
        RECT 27.690 203.315 28.040 204.515 ;
        RECT 28.400 203.905 28.780 205.550 ;
        RECT 27.480 202.520 27.830 202.580 ;
        RECT 28.400 202.520 28.740 203.125 ;
        RECT 26.610 202.260 28.740 202.520 ;
        RECT 27.480 202.200 27.830 202.260 ;
        RECT 29.010 201.980 29.610 205.975 ;
        RECT 31.455 205.540 33.205 208.325 ;
        RECT 33.845 205.540 34.655 206.540 ;
        RECT 35.295 205.540 37.045 207.835 ;
        RECT 37.685 205.540 38.495 206.540 ;
        RECT 39.135 205.540 40.885 207.835 ;
        RECT 41.525 205.540 42.335 206.540 ;
        RECT 42.975 205.540 44.725 207.835 ;
        RECT 45.365 205.540 46.175 206.540 ;
        RECT 46.815 205.540 48.565 207.835 ;
        RECT 49.205 205.540 50.015 206.540 ;
        RECT 50.655 205.540 52.405 207.835 ;
        RECT 53.045 205.540 53.855 206.540 ;
        RECT 54.495 205.540 56.245 207.835 ;
        RECT 56.885 205.540 57.695 206.540 ;
        RECT 58.335 205.540 60.085 207.835 ;
        RECT 60.725 205.540 61.535 206.540 ;
        RECT 63.905 205.540 65.655 208.325 ;
        RECT 66.295 205.540 67.105 206.540 ;
        RECT 67.745 205.540 69.495 207.835 ;
        RECT 70.135 205.540 70.945 206.540 ;
        RECT 71.585 205.540 73.335 207.835 ;
        RECT 73.975 205.540 74.785 206.540 ;
        RECT 75.425 205.540 77.175 207.835 ;
        RECT 77.815 205.540 78.625 206.540 ;
        RECT 79.265 205.540 81.015 207.835 ;
        RECT 81.655 205.540 82.465 206.540 ;
        RECT 83.105 205.540 84.855 207.835 ;
        RECT 85.495 205.540 86.305 206.540 ;
        RECT 86.945 205.540 88.695 207.835 ;
        RECT 89.335 205.540 90.145 206.540 ;
        RECT 90.785 205.540 92.535 207.835 ;
        RECT 93.175 205.540 93.985 206.540 ;
        RECT 96.355 205.540 98.105 208.325 ;
        RECT 98.745 205.540 99.555 206.540 ;
        RECT 100.195 205.540 101.945 207.835 ;
        RECT 102.585 205.540 103.395 206.540 ;
        RECT 104.035 205.540 105.785 207.835 ;
        RECT 106.425 205.540 107.235 206.540 ;
        RECT 107.875 205.540 109.625 207.835 ;
        RECT 110.265 205.540 111.075 206.540 ;
        RECT 111.715 205.540 113.465 207.835 ;
        RECT 114.105 205.540 114.915 206.540 ;
        RECT 115.555 205.540 117.305 207.835 ;
        RECT 117.945 205.540 118.755 206.540 ;
        RECT 119.395 205.540 121.145 207.835 ;
        RECT 121.785 205.540 122.595 206.540 ;
        RECT 123.235 205.540 124.985 207.835 ;
        RECT 125.625 205.540 126.435 206.540 ;
        RECT 128.805 205.540 130.555 208.325 ;
        RECT 131.195 205.540 132.005 206.540 ;
        RECT 132.645 205.540 134.395 207.835 ;
        RECT 135.035 205.540 135.845 206.540 ;
        RECT 136.485 205.540 138.235 207.835 ;
        RECT 138.875 205.540 139.685 206.540 ;
        RECT 140.325 205.540 142.075 207.835 ;
        RECT 142.715 205.540 143.525 206.540 ;
        RECT 144.165 205.540 145.915 207.835 ;
        RECT 146.555 205.540 147.365 206.540 ;
        RECT 148.005 205.540 149.755 207.835 ;
        RECT 150.395 205.540 151.205 206.540 ;
        RECT 151.845 205.540 153.595 207.835 ;
        RECT 154.235 205.540 155.045 206.540 ;
        RECT 155.685 205.540 157.435 207.835 ;
        RECT 158.075 205.540 158.885 206.540 ;
        RECT 161.300 205.730 161.670 224.240 ;
        RECT 162.320 220.605 162.690 224.240 ;
        RECT 162.315 220.225 162.695 220.605 ;
        RECT 162.320 217.605 162.690 220.225 ;
        RECT 162.315 217.225 162.695 217.605 ;
        RECT 162.320 214.605 162.690 217.225 ;
        RECT 162.315 214.225 162.695 214.605 ;
        RECT 162.320 211.605 162.690 214.225 ;
        RECT 162.315 211.225 162.695 211.605 ;
        RECT 162.320 208.605 162.690 211.225 ;
        RECT 162.315 208.225 162.695 208.605 ;
        RECT 161.300 205.350 161.680 205.730 ;
        RECT 161.300 204.280 161.670 205.350 ;
        RECT 31.925 203.090 32.735 204.090 ;
        RECT 25.090 201.650 26.780 201.880 ;
        RECT 28.150 201.750 29.610 201.980 ;
        RECT 25.090 199.640 25.690 201.650 ;
        RECT 27.110 201.190 28.110 201.515 ;
        RECT 25.920 200.630 28.780 200.960 ;
        RECT 25.090 199.410 26.780 199.640 ;
        RECT 25.090 197.400 25.690 199.410 ;
        RECT 27.495 199.275 27.760 200.630 ;
        RECT 29.010 199.740 29.610 201.750 ;
        RECT 33.375 201.260 35.125 204.090 ;
        RECT 35.765 203.090 36.575 204.090 ;
        RECT 37.215 201.795 38.965 204.090 ;
        RECT 39.605 203.090 40.415 204.090 ;
        RECT 41.055 201.795 42.805 204.090 ;
        RECT 43.445 203.090 44.255 204.090 ;
        RECT 44.895 201.795 46.645 204.090 ;
        RECT 47.285 203.090 48.095 204.090 ;
        RECT 48.735 201.795 50.485 204.090 ;
        RECT 51.125 203.090 51.935 204.090 ;
        RECT 52.575 201.795 54.325 204.090 ;
        RECT 54.965 203.090 55.775 204.090 ;
        RECT 56.415 201.795 58.165 204.090 ;
        RECT 58.805 203.090 59.615 204.090 ;
        RECT 60.255 201.795 62.005 204.090 ;
        RECT 64.375 203.090 65.185 204.090 ;
        RECT 65.825 201.260 67.575 204.090 ;
        RECT 68.215 203.090 69.025 204.090 ;
        RECT 69.665 201.795 71.415 204.090 ;
        RECT 72.055 203.090 72.865 204.090 ;
        RECT 73.505 201.795 75.255 204.090 ;
        RECT 75.895 203.090 76.705 204.090 ;
        RECT 77.345 201.795 79.095 204.090 ;
        RECT 79.735 203.090 80.545 204.090 ;
        RECT 81.185 201.795 82.935 204.090 ;
        RECT 83.575 203.090 84.385 204.090 ;
        RECT 85.025 201.795 86.775 204.090 ;
        RECT 87.415 203.090 88.225 204.090 ;
        RECT 88.865 201.795 90.615 204.090 ;
        RECT 91.255 203.090 92.065 204.090 ;
        RECT 92.705 201.795 94.455 204.090 ;
        RECT 96.825 203.090 97.635 204.090 ;
        RECT 98.275 201.260 100.025 204.090 ;
        RECT 100.665 203.090 101.475 204.090 ;
        RECT 102.115 201.795 103.865 204.090 ;
        RECT 104.505 203.090 105.315 204.090 ;
        RECT 105.955 201.795 107.705 204.090 ;
        RECT 108.345 203.090 109.155 204.090 ;
        RECT 109.795 201.795 111.545 204.090 ;
        RECT 112.185 203.090 112.995 204.090 ;
        RECT 113.635 201.795 115.385 204.090 ;
        RECT 116.025 203.090 116.835 204.090 ;
        RECT 117.475 201.795 119.225 204.090 ;
        RECT 119.865 203.090 120.675 204.090 ;
        RECT 121.315 201.795 123.065 204.090 ;
        RECT 123.705 203.090 124.515 204.090 ;
        RECT 125.155 201.795 126.905 204.090 ;
        RECT 129.275 203.090 130.085 204.090 ;
        RECT 130.725 201.260 132.475 204.090 ;
        RECT 133.115 203.090 133.925 204.090 ;
        RECT 134.565 201.795 136.315 204.090 ;
        RECT 136.955 203.090 137.765 204.090 ;
        RECT 138.405 201.795 140.155 204.090 ;
        RECT 140.795 203.090 141.605 204.090 ;
        RECT 142.245 201.795 143.995 204.090 ;
        RECT 144.635 203.090 145.445 204.090 ;
        RECT 146.085 201.795 147.835 204.090 ;
        RECT 148.475 203.090 149.285 204.090 ;
        RECT 149.925 201.795 151.675 204.090 ;
        RECT 152.315 203.090 153.125 204.090 ;
        RECT 153.765 201.795 155.515 204.090 ;
        RECT 156.155 203.090 156.965 204.090 ;
        RECT 157.605 201.795 159.355 204.090 ;
        RECT 161.300 203.900 161.680 204.280 ;
        RECT 31.650 200.890 62.170 201.260 ;
        RECT 64.100 200.890 94.620 201.260 ;
        RECT 96.550 200.890 127.070 201.260 ;
        RECT 129.000 200.890 159.520 201.260 ;
        RECT 30.800 200.625 31.420 200.810 ;
        RECT 62.400 200.625 63.020 200.810 ;
        RECT 30.800 200.395 63.020 200.625 ;
        RECT 30.800 200.210 31.420 200.395 ;
        RECT 62.400 200.210 63.020 200.395 ;
        RECT 63.250 200.625 63.870 200.810 ;
        RECT 94.850 200.625 95.470 200.810 ;
        RECT 63.250 200.395 95.470 200.625 ;
        RECT 63.250 200.210 63.870 200.395 ;
        RECT 94.850 200.210 95.470 200.395 ;
        RECT 95.700 200.625 96.320 200.810 ;
        RECT 127.300 200.625 127.920 200.810 ;
        RECT 95.700 200.395 127.920 200.625 ;
        RECT 95.700 200.210 96.320 200.395 ;
        RECT 127.300 200.210 127.920 200.395 ;
        RECT 128.150 200.625 128.770 200.810 ;
        RECT 159.750 200.625 160.370 200.810 ;
        RECT 128.150 200.395 160.370 200.625 ;
        RECT 128.150 200.210 128.770 200.395 ;
        RECT 159.750 200.210 160.370 200.395 ;
        RECT 31.650 199.760 62.170 200.140 ;
        RECT 64.100 199.760 94.620 200.140 ;
        RECT 96.550 199.760 127.070 200.140 ;
        RECT 129.000 199.760 159.520 200.140 ;
        RECT 28.150 199.510 29.610 199.740 ;
        RECT 27.110 198.950 28.110 199.275 ;
        RECT 25.920 198.390 28.780 198.720 ;
        RECT 29.010 197.500 29.610 199.510 ;
        RECT 31.650 199.050 62.170 199.420 ;
        RECT 64.100 199.050 94.620 199.420 ;
        RECT 96.550 199.050 127.070 199.420 ;
        RECT 129.000 199.050 159.520 199.420 ;
        RECT 37.280 199.040 38.900 199.050 ;
        RECT 69.730 199.040 71.350 199.050 ;
        RECT 102.180 199.040 103.800 199.050 ;
        RECT 134.630 199.040 136.250 199.050 ;
        RECT 30.800 198.785 31.420 198.970 ;
        RECT 62.400 198.785 63.020 198.970 ;
        RECT 30.800 198.555 63.020 198.785 ;
        RECT 30.800 198.370 31.420 198.555 ;
        RECT 62.400 198.370 63.020 198.555 ;
        RECT 63.250 198.785 63.870 198.970 ;
        RECT 94.850 198.785 95.470 198.970 ;
        RECT 63.250 198.555 95.470 198.785 ;
        RECT 63.250 198.370 63.870 198.555 ;
        RECT 94.850 198.370 95.470 198.555 ;
        RECT 95.700 198.785 96.320 198.970 ;
        RECT 127.300 198.785 127.920 198.970 ;
        RECT 95.700 198.555 127.920 198.785 ;
        RECT 95.700 198.370 96.320 198.555 ;
        RECT 127.300 198.370 127.920 198.555 ;
        RECT 128.150 198.785 128.770 198.970 ;
        RECT 159.750 198.785 160.370 198.970 ;
        RECT 128.150 198.555 160.370 198.785 ;
        RECT 128.150 198.370 128.770 198.555 ;
        RECT 159.750 198.370 160.370 198.555 ;
        RECT 31.650 197.920 62.170 198.300 ;
        RECT 64.100 197.920 94.620 198.300 ;
        RECT 96.550 197.920 127.070 198.300 ;
        RECT 129.000 197.920 159.520 198.300 ;
        RECT 25.090 197.170 26.780 197.400 ;
        RECT 28.150 197.270 29.610 197.500 ;
        RECT 25.090 195.115 25.690 197.170 ;
        RECT 27.110 196.710 28.110 197.035 ;
        RECT 29.010 195.115 29.610 197.270 ;
        RECT 31.650 197.205 62.170 197.575 ;
        RECT 64.100 197.205 94.620 197.575 ;
        RECT 96.550 197.205 127.070 197.575 ;
        RECT 129.000 197.205 159.520 197.575 ;
        RECT 41.120 197.195 42.740 197.205 ;
        RECT 73.570 197.195 75.190 197.205 ;
        RECT 106.020 197.195 107.640 197.205 ;
        RECT 138.470 197.195 140.090 197.205 ;
        RECT 30.800 196.940 31.420 197.125 ;
        RECT 62.400 196.940 63.020 197.125 ;
        RECT 30.800 196.710 63.020 196.940 ;
        RECT 30.800 196.525 31.420 196.710 ;
        RECT 62.400 196.525 63.020 196.710 ;
        RECT 63.250 196.940 63.870 197.125 ;
        RECT 94.850 196.940 95.470 197.125 ;
        RECT 63.250 196.710 95.470 196.940 ;
        RECT 63.250 196.525 63.870 196.710 ;
        RECT 94.850 196.525 95.470 196.710 ;
        RECT 95.700 196.940 96.320 197.125 ;
        RECT 127.300 196.940 127.920 197.125 ;
        RECT 95.700 196.710 127.920 196.940 ;
        RECT 95.700 196.525 96.320 196.710 ;
        RECT 127.300 196.525 127.920 196.710 ;
        RECT 128.150 196.940 128.770 197.125 ;
        RECT 159.750 196.940 160.370 197.125 ;
        RECT 128.150 196.710 160.370 196.940 ;
        RECT 128.150 196.525 128.770 196.710 ;
        RECT 159.750 196.525 160.370 196.710 ;
        RECT 31.650 196.075 62.170 196.455 ;
        RECT 64.100 196.075 94.620 196.455 ;
        RECT 96.550 196.075 127.070 196.455 ;
        RECT 129.000 196.075 159.520 196.455 ;
        RECT 31.660 195.285 62.160 195.725 ;
        RECT 64.110 195.285 94.610 195.725 ;
        RECT 96.560 195.285 127.060 195.725 ;
        RECT 129.010 195.285 159.510 195.725 ;
        RECT 25.090 194.775 27.380 195.115 ;
        RECT 28.125 194.775 29.610 195.115 ;
        RECT 25.090 166.930 25.690 194.775 ;
        RECT 29.010 166.930 29.610 194.775 ;
        RECT 31.650 194.565 62.170 194.935 ;
        RECT 64.100 194.565 94.620 194.935 ;
        RECT 96.550 194.565 127.070 194.935 ;
        RECT 129.000 194.565 159.520 194.935 ;
        RECT 44.960 194.555 46.580 194.565 ;
        RECT 77.410 194.555 79.030 194.565 ;
        RECT 109.860 194.555 111.480 194.565 ;
        RECT 142.310 194.555 143.930 194.565 ;
        RECT 30.800 194.300 31.420 194.485 ;
        RECT 62.400 194.300 63.020 194.485 ;
        RECT 30.800 194.070 63.020 194.300 ;
        RECT 30.800 193.885 31.420 194.070 ;
        RECT 62.400 193.885 63.020 194.070 ;
        RECT 63.250 194.300 63.870 194.485 ;
        RECT 94.850 194.300 95.470 194.485 ;
        RECT 63.250 194.070 95.470 194.300 ;
        RECT 63.250 193.885 63.870 194.070 ;
        RECT 94.850 193.885 95.470 194.070 ;
        RECT 95.700 194.300 96.320 194.485 ;
        RECT 127.300 194.300 127.920 194.485 ;
        RECT 95.700 194.070 127.920 194.300 ;
        RECT 95.700 193.885 96.320 194.070 ;
        RECT 127.300 193.885 127.920 194.070 ;
        RECT 128.150 194.300 128.770 194.485 ;
        RECT 159.750 194.300 160.370 194.485 ;
        RECT 128.150 194.070 160.370 194.300 ;
        RECT 128.150 193.885 128.770 194.070 ;
        RECT 159.750 193.885 160.370 194.070 ;
        RECT 31.650 193.435 62.170 193.815 ;
        RECT 64.100 193.435 94.620 193.815 ;
        RECT 96.550 193.435 127.070 193.815 ;
        RECT 129.000 193.435 159.520 193.815 ;
        RECT 31.650 192.725 62.170 193.095 ;
        RECT 64.100 192.725 94.620 193.095 ;
        RECT 96.550 192.725 127.070 193.095 ;
        RECT 129.000 192.725 159.520 193.095 ;
        RECT 48.800 192.715 50.420 192.725 ;
        RECT 81.250 192.715 82.870 192.725 ;
        RECT 113.700 192.715 115.320 192.725 ;
        RECT 146.150 192.715 147.770 192.725 ;
        RECT 30.800 192.460 31.420 192.645 ;
        RECT 62.400 192.460 63.020 192.645 ;
        RECT 30.800 192.230 63.020 192.460 ;
        RECT 30.800 192.045 31.420 192.230 ;
        RECT 62.400 192.045 63.020 192.230 ;
        RECT 63.250 192.460 63.870 192.645 ;
        RECT 94.850 192.460 95.470 192.645 ;
        RECT 63.250 192.230 95.470 192.460 ;
        RECT 63.250 192.045 63.870 192.230 ;
        RECT 94.850 192.045 95.470 192.230 ;
        RECT 95.700 192.460 96.320 192.645 ;
        RECT 127.300 192.460 127.920 192.645 ;
        RECT 95.700 192.230 127.920 192.460 ;
        RECT 95.700 192.045 96.320 192.230 ;
        RECT 127.300 192.045 127.920 192.230 ;
        RECT 128.150 192.460 128.770 192.645 ;
        RECT 159.750 192.460 160.370 192.645 ;
        RECT 128.150 192.230 160.370 192.460 ;
        RECT 128.150 192.045 128.770 192.230 ;
        RECT 159.750 192.045 160.370 192.230 ;
        RECT 31.650 191.595 62.170 191.975 ;
        RECT 64.100 191.595 94.620 191.975 ;
        RECT 96.550 191.595 127.070 191.975 ;
        RECT 129.000 191.595 159.520 191.975 ;
        RECT 31.650 190.880 62.170 191.250 ;
        RECT 64.100 190.880 94.620 191.250 ;
        RECT 96.550 190.880 127.070 191.250 ;
        RECT 129.000 190.880 159.520 191.250 ;
        RECT 52.640 190.870 54.260 190.880 ;
        RECT 85.090 190.870 86.710 190.880 ;
        RECT 117.540 190.870 119.160 190.880 ;
        RECT 149.990 190.870 151.610 190.880 ;
        RECT 30.800 190.615 31.420 190.800 ;
        RECT 62.400 190.615 63.020 190.800 ;
        RECT 30.800 190.385 63.020 190.615 ;
        RECT 30.800 190.200 31.420 190.385 ;
        RECT 62.400 190.200 63.020 190.385 ;
        RECT 63.250 190.615 63.870 190.800 ;
        RECT 94.850 190.615 95.470 190.800 ;
        RECT 63.250 190.385 95.470 190.615 ;
        RECT 63.250 190.200 63.870 190.385 ;
        RECT 94.850 190.200 95.470 190.385 ;
        RECT 95.700 190.615 96.320 190.800 ;
        RECT 127.300 190.615 127.920 190.800 ;
        RECT 95.700 190.385 127.920 190.615 ;
        RECT 95.700 190.200 96.320 190.385 ;
        RECT 127.300 190.200 127.920 190.385 ;
        RECT 128.150 190.615 128.770 190.800 ;
        RECT 159.750 190.615 160.370 190.800 ;
        RECT 128.150 190.385 160.370 190.615 ;
        RECT 128.150 190.200 128.770 190.385 ;
        RECT 159.750 190.200 160.370 190.385 ;
        RECT 31.650 189.750 62.170 190.130 ;
        RECT 64.100 189.750 94.620 190.130 ;
        RECT 96.550 189.750 127.070 190.130 ;
        RECT 129.000 189.750 159.520 190.130 ;
        RECT 31.660 188.960 62.160 189.400 ;
        RECT 64.110 188.960 94.610 189.400 ;
        RECT 96.560 188.960 127.060 189.400 ;
        RECT 129.010 188.960 159.510 189.400 ;
        RECT 31.650 188.240 62.170 188.610 ;
        RECT 64.100 188.240 94.620 188.610 ;
        RECT 96.550 188.240 127.070 188.610 ;
        RECT 129.000 188.240 159.520 188.610 ;
        RECT 56.480 188.230 58.100 188.240 ;
        RECT 88.930 188.230 90.550 188.240 ;
        RECT 121.380 188.230 123.000 188.240 ;
        RECT 153.830 188.230 155.450 188.240 ;
        RECT 30.800 187.975 31.420 188.160 ;
        RECT 62.400 187.975 63.020 188.160 ;
        RECT 30.800 187.745 63.020 187.975 ;
        RECT 30.800 187.560 31.420 187.745 ;
        RECT 62.400 187.560 63.020 187.745 ;
        RECT 63.250 187.975 63.870 188.160 ;
        RECT 94.850 187.975 95.470 188.160 ;
        RECT 63.250 187.745 95.470 187.975 ;
        RECT 63.250 187.560 63.870 187.745 ;
        RECT 94.850 187.560 95.470 187.745 ;
        RECT 95.700 187.975 96.320 188.160 ;
        RECT 127.300 187.975 127.920 188.160 ;
        RECT 95.700 187.745 127.920 187.975 ;
        RECT 95.700 187.560 96.320 187.745 ;
        RECT 127.300 187.560 127.920 187.745 ;
        RECT 128.150 187.975 128.770 188.160 ;
        RECT 159.750 187.975 160.370 188.160 ;
        RECT 128.150 187.745 160.370 187.975 ;
        RECT 128.150 187.560 128.770 187.745 ;
        RECT 159.750 187.560 160.370 187.745 ;
        RECT 31.650 187.110 62.170 187.490 ;
        RECT 64.100 187.110 94.620 187.490 ;
        RECT 96.550 187.110 127.070 187.490 ;
        RECT 129.000 187.110 159.520 187.490 ;
        RECT 31.650 186.400 62.170 186.770 ;
        RECT 64.100 186.400 94.620 186.770 ;
        RECT 96.550 186.400 127.070 186.770 ;
        RECT 129.000 186.400 159.520 186.770 ;
        RECT 60.320 186.390 61.940 186.400 ;
        RECT 92.770 186.390 94.390 186.400 ;
        RECT 125.220 186.390 126.840 186.400 ;
        RECT 157.670 186.390 159.290 186.400 ;
        RECT 30.800 186.135 31.420 186.320 ;
        RECT 62.400 186.135 63.020 186.320 ;
        RECT 30.800 185.905 63.020 186.135 ;
        RECT 30.800 185.720 31.420 185.905 ;
        RECT 62.400 185.720 63.020 185.905 ;
        RECT 63.250 186.135 63.870 186.320 ;
        RECT 94.850 186.135 95.470 186.320 ;
        RECT 63.250 185.905 95.470 186.135 ;
        RECT 63.250 185.720 63.870 185.905 ;
        RECT 94.850 185.720 95.470 185.905 ;
        RECT 95.700 186.135 96.320 186.320 ;
        RECT 127.300 186.135 127.920 186.320 ;
        RECT 95.700 185.905 127.920 186.135 ;
        RECT 95.700 185.720 96.320 185.905 ;
        RECT 127.300 185.720 127.920 185.905 ;
        RECT 128.150 186.135 128.770 186.320 ;
        RECT 159.750 186.135 160.370 186.320 ;
        RECT 128.150 185.905 160.370 186.135 ;
        RECT 161.300 185.970 161.670 203.900 ;
        RECT 162.320 202.605 162.690 208.225 ;
        RECT 163.340 205.730 163.710 224.240 ;
        RECT 164.360 220.605 164.730 224.240 ;
        RECT 164.355 220.225 164.735 220.605 ;
        RECT 164.360 217.605 164.730 220.225 ;
        RECT 164.355 217.225 164.735 217.605 ;
        RECT 164.360 214.605 164.730 217.225 ;
        RECT 164.355 214.225 164.735 214.605 ;
        RECT 164.360 211.605 164.730 214.225 ;
        RECT 164.355 211.225 164.735 211.605 ;
        RECT 164.360 208.605 164.730 211.225 ;
        RECT 164.355 208.225 164.735 208.605 ;
        RECT 163.340 205.350 163.720 205.730 ;
        RECT 163.340 204.280 163.710 205.350 ;
        RECT 163.340 203.900 163.720 204.280 ;
        RECT 162.315 202.225 162.695 202.605 ;
        RECT 162.320 199.605 162.690 202.225 ;
        RECT 162.315 199.225 162.695 199.605 ;
        RECT 162.320 196.605 162.690 199.225 ;
        RECT 162.315 196.225 162.695 196.605 ;
        RECT 162.320 193.605 162.690 196.225 ;
        RECT 162.315 193.225 162.695 193.605 ;
        RECT 162.320 190.605 162.690 193.225 ;
        RECT 162.315 190.225 162.695 190.605 ;
        RECT 162.320 187.605 162.690 190.225 ;
        RECT 162.315 187.225 162.695 187.605 ;
        RECT 162.320 185.970 162.690 187.225 ;
        RECT 163.340 185.970 163.710 203.900 ;
        RECT 164.360 202.605 164.730 208.225 ;
        RECT 164.355 202.225 164.735 202.605 ;
        RECT 164.360 199.605 164.730 202.225 ;
        RECT 164.355 199.225 164.735 199.605 ;
        RECT 164.360 196.605 164.730 199.225 ;
        RECT 164.355 196.225 164.735 196.605 ;
        RECT 164.360 193.605 164.730 196.225 ;
        RECT 164.355 193.225 164.735 193.605 ;
        RECT 164.360 190.605 164.730 193.225 ;
        RECT 164.355 190.225 164.735 190.605 ;
        RECT 164.360 187.605 164.730 190.225 ;
        RECT 164.355 187.225 164.735 187.605 ;
        RECT 164.360 185.970 164.730 187.225 ;
        RECT 165.380 185.970 165.760 224.240 ;
        RECT 166.110 185.980 166.550 224.230 ;
        RECT 128.150 185.720 128.770 185.905 ;
        RECT 159.750 185.720 160.370 185.905 ;
        RECT 31.650 185.270 62.170 185.650 ;
        RECT 64.100 185.270 94.620 185.650 ;
        RECT 96.550 185.270 127.070 185.650 ;
        RECT 129.000 185.270 159.520 185.650 ;
        RECT 31.650 184.550 62.170 184.930 ;
        RECT 64.100 184.550 94.620 184.930 ;
        RECT 96.550 184.550 127.070 184.930 ;
        RECT 129.000 184.550 159.520 184.930 ;
        RECT 30.800 184.295 31.420 184.480 ;
        RECT 62.400 184.295 63.020 184.480 ;
        RECT 30.800 184.065 63.020 184.295 ;
        RECT 30.800 183.880 31.420 184.065 ;
        RECT 62.400 183.880 63.020 184.065 ;
        RECT 63.250 184.295 63.870 184.480 ;
        RECT 94.850 184.295 95.470 184.480 ;
        RECT 63.250 184.065 95.470 184.295 ;
        RECT 63.250 183.880 63.870 184.065 ;
        RECT 94.850 183.880 95.470 184.065 ;
        RECT 95.700 184.295 96.320 184.480 ;
        RECT 127.300 184.295 127.920 184.480 ;
        RECT 95.700 184.065 127.920 184.295 ;
        RECT 95.700 183.880 96.320 184.065 ;
        RECT 127.300 183.880 127.920 184.065 ;
        RECT 128.150 184.295 128.770 184.480 ;
        RECT 159.750 184.295 160.370 184.480 ;
        RECT 128.150 184.065 160.370 184.295 ;
        RECT 128.150 183.880 128.770 184.065 ;
        RECT 159.750 183.880 160.370 184.065 ;
        RECT 58.400 183.800 60.020 183.810 ;
        RECT 90.850 183.800 92.470 183.810 ;
        RECT 123.300 183.800 124.920 183.810 ;
        RECT 155.750 183.800 157.370 183.810 ;
        RECT 31.650 183.430 62.170 183.800 ;
        RECT 64.100 183.430 94.620 183.800 ;
        RECT 96.550 183.430 127.070 183.800 ;
        RECT 129.000 183.430 159.520 183.800 ;
        RECT 31.650 182.710 62.170 183.090 ;
        RECT 64.100 182.710 94.620 183.090 ;
        RECT 96.550 182.710 127.070 183.090 ;
        RECT 129.000 182.710 159.520 183.090 ;
        RECT 30.800 182.455 31.420 182.640 ;
        RECT 62.400 182.455 63.020 182.640 ;
        RECT 30.800 182.225 63.020 182.455 ;
        RECT 30.800 182.040 31.420 182.225 ;
        RECT 62.400 182.040 63.020 182.225 ;
        RECT 63.250 182.455 63.870 182.640 ;
        RECT 94.850 182.455 95.470 182.640 ;
        RECT 63.250 182.225 95.470 182.455 ;
        RECT 63.250 182.040 63.870 182.225 ;
        RECT 94.850 182.040 95.470 182.225 ;
        RECT 95.700 182.455 96.320 182.640 ;
        RECT 127.300 182.455 127.920 182.640 ;
        RECT 95.700 182.225 127.920 182.455 ;
        RECT 95.700 182.040 96.320 182.225 ;
        RECT 127.300 182.040 127.920 182.225 ;
        RECT 128.150 182.455 128.770 182.640 ;
        RECT 159.750 182.455 160.370 182.640 ;
        RECT 128.150 182.225 160.370 182.455 ;
        RECT 128.150 182.040 128.770 182.225 ;
        RECT 159.750 182.040 160.370 182.225 ;
        RECT 54.560 181.960 56.180 181.970 ;
        RECT 87.010 181.960 88.630 181.970 ;
        RECT 119.460 181.960 121.080 181.970 ;
        RECT 151.910 181.960 153.530 181.970 ;
        RECT 31.650 181.590 62.170 181.960 ;
        RECT 64.100 181.590 94.620 181.960 ;
        RECT 96.550 181.590 127.070 181.960 ;
        RECT 129.000 181.590 159.520 181.960 ;
        RECT 31.660 180.795 62.160 181.235 ;
        RECT 64.110 180.795 94.610 181.235 ;
        RECT 96.560 180.795 127.060 181.235 ;
        RECT 129.010 180.795 159.510 181.235 ;
        RECT 31.650 180.065 62.170 180.445 ;
        RECT 64.100 180.065 94.620 180.445 ;
        RECT 96.550 180.065 127.070 180.445 ;
        RECT 129.000 180.065 159.520 180.445 ;
        RECT 30.800 179.810 31.420 179.995 ;
        RECT 62.400 179.810 63.020 179.995 ;
        RECT 30.800 179.580 63.020 179.810 ;
        RECT 30.800 179.395 31.420 179.580 ;
        RECT 62.400 179.395 63.020 179.580 ;
        RECT 63.250 179.810 63.870 179.995 ;
        RECT 94.850 179.810 95.470 179.995 ;
        RECT 63.250 179.580 95.470 179.810 ;
        RECT 63.250 179.395 63.870 179.580 ;
        RECT 94.850 179.395 95.470 179.580 ;
        RECT 95.700 179.810 96.320 179.995 ;
        RECT 127.300 179.810 127.920 179.995 ;
        RECT 95.700 179.580 127.920 179.810 ;
        RECT 95.700 179.395 96.320 179.580 ;
        RECT 127.300 179.395 127.920 179.580 ;
        RECT 128.150 179.810 128.770 179.995 ;
        RECT 159.750 179.810 160.370 179.995 ;
        RECT 128.150 179.580 160.370 179.810 ;
        RECT 128.150 179.395 128.770 179.580 ;
        RECT 159.750 179.395 160.370 179.580 ;
        RECT 50.720 179.315 52.340 179.325 ;
        RECT 83.170 179.315 84.790 179.325 ;
        RECT 115.620 179.315 117.240 179.325 ;
        RECT 148.070 179.315 149.690 179.325 ;
        RECT 31.650 178.945 62.170 179.315 ;
        RECT 64.100 178.945 94.620 179.315 ;
        RECT 96.550 178.945 127.070 179.315 ;
        RECT 129.000 178.945 159.520 179.315 ;
        RECT 31.650 178.225 62.170 178.605 ;
        RECT 64.100 178.225 94.620 178.605 ;
        RECT 96.550 178.225 127.070 178.605 ;
        RECT 129.000 178.225 159.520 178.605 ;
        RECT 30.800 177.970 31.420 178.155 ;
        RECT 62.400 177.970 63.020 178.155 ;
        RECT 30.800 177.740 63.020 177.970 ;
        RECT 30.800 177.555 31.420 177.740 ;
        RECT 62.400 177.555 63.020 177.740 ;
        RECT 63.250 177.970 63.870 178.155 ;
        RECT 94.850 177.970 95.470 178.155 ;
        RECT 63.250 177.740 95.470 177.970 ;
        RECT 63.250 177.555 63.870 177.740 ;
        RECT 94.850 177.555 95.470 177.740 ;
        RECT 95.700 177.970 96.320 178.155 ;
        RECT 127.300 177.970 127.920 178.155 ;
        RECT 95.700 177.740 127.920 177.970 ;
        RECT 95.700 177.555 96.320 177.740 ;
        RECT 127.300 177.555 127.920 177.740 ;
        RECT 128.150 177.970 128.770 178.155 ;
        RECT 159.750 177.970 160.370 178.155 ;
        RECT 128.150 177.740 160.370 177.970 ;
        RECT 128.150 177.555 128.770 177.740 ;
        RECT 159.750 177.555 160.370 177.740 ;
        RECT 46.880 177.475 48.500 177.485 ;
        RECT 79.330 177.475 80.950 177.485 ;
        RECT 111.780 177.475 113.400 177.485 ;
        RECT 144.230 177.475 145.850 177.485 ;
        RECT 31.650 177.105 62.170 177.475 ;
        RECT 64.100 177.105 94.620 177.475 ;
        RECT 96.550 177.105 127.070 177.475 ;
        RECT 129.000 177.105 159.520 177.475 ;
        RECT 31.650 176.385 62.170 176.765 ;
        RECT 64.100 176.385 94.620 176.765 ;
        RECT 96.550 176.385 127.070 176.765 ;
        RECT 129.000 176.385 159.520 176.765 ;
        RECT 30.800 176.130 31.420 176.315 ;
        RECT 62.400 176.130 63.020 176.315 ;
        RECT 30.800 175.900 63.020 176.130 ;
        RECT 30.800 175.715 31.420 175.900 ;
        RECT 62.400 175.715 63.020 175.900 ;
        RECT 63.250 176.130 63.870 176.315 ;
        RECT 94.850 176.130 95.470 176.315 ;
        RECT 63.250 175.900 95.470 176.130 ;
        RECT 63.250 175.715 63.870 175.900 ;
        RECT 94.850 175.715 95.470 175.900 ;
        RECT 95.700 176.130 96.320 176.315 ;
        RECT 127.300 176.130 127.920 176.315 ;
        RECT 95.700 175.900 127.920 176.130 ;
        RECT 95.700 175.715 96.320 175.900 ;
        RECT 127.300 175.715 127.920 175.900 ;
        RECT 128.150 176.130 128.770 176.315 ;
        RECT 159.750 176.130 160.370 176.315 ;
        RECT 128.150 175.900 160.370 176.130 ;
        RECT 128.150 175.715 128.770 175.900 ;
        RECT 159.750 175.715 160.370 175.900 ;
        RECT 43.040 175.635 44.660 175.645 ;
        RECT 75.490 175.635 77.110 175.645 ;
        RECT 107.940 175.635 109.560 175.645 ;
        RECT 140.390 175.635 142.010 175.645 ;
        RECT 31.650 175.265 62.170 175.635 ;
        RECT 64.100 175.265 94.620 175.635 ;
        RECT 96.550 175.265 127.070 175.635 ;
        RECT 129.000 175.265 159.520 175.635 ;
        RECT 31.660 174.470 62.160 174.910 ;
        RECT 64.110 174.470 94.610 174.910 ;
        RECT 96.560 174.470 127.060 174.910 ;
        RECT 129.010 174.470 159.510 174.910 ;
        RECT 31.650 173.740 62.170 174.120 ;
        RECT 64.100 173.740 94.620 174.120 ;
        RECT 96.550 173.740 127.070 174.120 ;
        RECT 129.000 173.740 159.520 174.120 ;
        RECT 30.800 173.485 31.420 173.670 ;
        RECT 62.400 173.485 63.020 173.670 ;
        RECT 30.800 173.255 63.020 173.485 ;
        RECT 30.800 173.070 31.420 173.255 ;
        RECT 62.400 173.070 63.020 173.255 ;
        RECT 63.250 173.485 63.870 173.670 ;
        RECT 94.850 173.485 95.470 173.670 ;
        RECT 63.250 173.255 95.470 173.485 ;
        RECT 63.250 173.070 63.870 173.255 ;
        RECT 94.850 173.070 95.470 173.255 ;
        RECT 95.700 173.485 96.320 173.670 ;
        RECT 127.300 173.485 127.920 173.670 ;
        RECT 95.700 173.255 127.920 173.485 ;
        RECT 95.700 173.070 96.320 173.255 ;
        RECT 127.300 173.070 127.920 173.255 ;
        RECT 128.150 173.485 128.770 173.670 ;
        RECT 159.750 173.485 160.370 173.670 ;
        RECT 128.150 173.255 160.370 173.485 ;
        RECT 128.150 173.070 128.770 173.255 ;
        RECT 159.750 173.070 160.370 173.255 ;
        RECT 39.200 172.990 40.820 173.000 ;
        RECT 71.650 172.990 73.270 173.000 ;
        RECT 104.100 172.990 105.720 173.000 ;
        RECT 136.550 172.990 138.170 173.000 ;
        RECT 31.650 172.620 62.170 172.990 ;
        RECT 64.100 172.620 94.620 172.990 ;
        RECT 96.550 172.620 127.070 172.990 ;
        RECT 129.000 172.620 159.520 172.990 ;
        RECT 31.650 171.900 62.170 172.280 ;
        RECT 64.100 171.900 94.620 172.280 ;
        RECT 96.550 171.900 127.070 172.280 ;
        RECT 129.000 171.900 159.520 172.280 ;
        RECT 30.800 171.645 31.420 171.830 ;
        RECT 62.400 171.645 63.020 171.830 ;
        RECT 30.800 171.415 63.020 171.645 ;
        RECT 30.800 171.230 31.420 171.415 ;
        RECT 62.400 171.230 63.020 171.415 ;
        RECT 63.250 171.645 63.870 171.830 ;
        RECT 94.850 171.645 95.470 171.830 ;
        RECT 63.250 171.415 95.470 171.645 ;
        RECT 63.250 171.230 63.870 171.415 ;
        RECT 94.850 171.230 95.470 171.415 ;
        RECT 95.700 171.645 96.320 171.830 ;
        RECT 127.300 171.645 127.920 171.830 ;
        RECT 95.700 171.415 127.920 171.645 ;
        RECT 95.700 171.230 96.320 171.415 ;
        RECT 127.300 171.230 127.920 171.415 ;
        RECT 128.150 171.645 128.770 171.830 ;
        RECT 159.750 171.645 160.370 171.830 ;
        RECT 128.150 171.415 160.370 171.645 ;
        RECT 128.150 171.230 128.770 171.415 ;
        RECT 159.750 171.230 160.370 171.415 ;
        RECT 35.360 171.150 36.980 171.160 ;
        RECT 67.810 171.150 69.430 171.160 ;
        RECT 100.260 171.150 101.880 171.160 ;
        RECT 132.710 171.150 134.330 171.160 ;
        RECT 31.650 170.780 62.170 171.150 ;
        RECT 64.100 170.780 94.620 171.150 ;
        RECT 96.550 170.780 127.070 171.150 ;
        RECT 129.000 170.780 159.520 171.150 ;
        RECT 31.650 170.060 62.170 170.440 ;
        RECT 64.100 170.060 94.620 170.440 ;
        RECT 96.550 170.060 127.070 170.440 ;
        RECT 129.000 170.060 159.520 170.440 ;
        RECT 30.800 169.805 31.420 169.990 ;
        RECT 62.400 169.805 63.020 169.990 ;
        RECT 30.800 169.575 63.020 169.805 ;
        RECT 30.800 169.390 31.420 169.575 ;
        RECT 62.400 169.390 63.020 169.575 ;
        RECT 63.250 169.805 63.870 169.990 ;
        RECT 94.850 169.805 95.470 169.990 ;
        RECT 63.250 169.575 95.470 169.805 ;
        RECT 63.250 169.390 63.870 169.575 ;
        RECT 94.850 169.390 95.470 169.575 ;
        RECT 95.700 169.805 96.320 169.990 ;
        RECT 127.300 169.805 127.920 169.990 ;
        RECT 95.700 169.575 127.920 169.805 ;
        RECT 95.700 169.390 96.320 169.575 ;
        RECT 127.300 169.390 127.920 169.575 ;
        RECT 128.150 169.805 128.770 169.990 ;
        RECT 159.750 169.805 160.370 169.990 ;
        RECT 128.150 169.575 160.370 169.805 ;
        RECT 128.150 169.390 128.770 169.575 ;
        RECT 159.750 169.390 160.370 169.575 ;
        RECT 31.650 168.940 62.170 169.310 ;
        RECT 64.100 168.940 94.620 169.310 ;
        RECT 96.550 168.940 127.070 169.310 ;
        RECT 129.000 168.940 159.520 169.310 ;
        RECT 25.090 166.590 27.380 166.930 ;
        RECT 28.125 166.590 29.610 166.930 ;
        RECT 25.090 165.955 25.690 166.590 ;
        RECT 25.090 165.725 26.670 165.955 ;
        RECT 25.090 163.685 25.690 165.725 ;
        RECT 27.100 165.495 27.460 165.580 ;
        RECT 25.970 165.265 27.460 165.495 ;
        RECT 25.970 165.115 26.330 165.265 ;
        RECT 25.920 164.480 26.870 164.885 ;
        RECT 25.090 163.455 26.380 163.685 ;
        RECT 25.090 162.495 25.690 163.455 ;
        RECT 26.610 163.135 26.870 164.480 ;
        RECT 27.100 163.830 27.460 165.265 ;
        RECT 27.690 163.930 28.040 165.130 ;
        RECT 28.400 164.520 28.780 166.165 ;
        RECT 27.480 163.135 27.830 163.195 ;
        RECT 28.400 163.135 28.740 163.740 ;
        RECT 26.610 162.875 28.740 163.135 ;
        RECT 27.480 162.815 27.830 162.875 ;
        RECT 29.010 162.595 29.610 166.590 ;
        RECT 31.455 166.155 33.205 168.940 ;
        RECT 33.845 166.155 34.655 167.155 ;
        RECT 35.295 166.155 37.045 168.450 ;
        RECT 37.685 166.155 38.495 167.155 ;
        RECT 39.135 166.155 40.885 168.450 ;
        RECT 41.525 166.155 42.335 167.155 ;
        RECT 42.975 166.155 44.725 168.450 ;
        RECT 45.365 166.155 46.175 167.155 ;
        RECT 46.815 166.155 48.565 168.450 ;
        RECT 49.205 166.155 50.015 167.155 ;
        RECT 50.655 166.155 52.405 168.450 ;
        RECT 53.045 166.155 53.855 167.155 ;
        RECT 54.495 166.155 56.245 168.450 ;
        RECT 56.885 166.155 57.695 167.155 ;
        RECT 58.335 166.155 60.085 168.450 ;
        RECT 60.725 166.155 61.535 167.155 ;
        RECT 63.905 166.155 65.655 168.940 ;
        RECT 66.295 166.155 67.105 167.155 ;
        RECT 67.745 166.155 69.495 168.450 ;
        RECT 70.135 166.155 70.945 167.155 ;
        RECT 71.585 166.155 73.335 168.450 ;
        RECT 73.975 166.155 74.785 167.155 ;
        RECT 75.425 166.155 77.175 168.450 ;
        RECT 77.815 166.155 78.625 167.155 ;
        RECT 79.265 166.155 81.015 168.450 ;
        RECT 81.655 166.155 82.465 167.155 ;
        RECT 83.105 166.155 84.855 168.450 ;
        RECT 85.495 166.155 86.305 167.155 ;
        RECT 86.945 166.155 88.695 168.450 ;
        RECT 89.335 166.155 90.145 167.155 ;
        RECT 90.785 166.155 92.535 168.450 ;
        RECT 93.175 166.155 93.985 167.155 ;
        RECT 96.355 166.155 98.105 168.940 ;
        RECT 98.745 166.155 99.555 167.155 ;
        RECT 100.195 166.155 101.945 168.450 ;
        RECT 102.585 166.155 103.395 167.155 ;
        RECT 104.035 166.155 105.785 168.450 ;
        RECT 106.425 166.155 107.235 167.155 ;
        RECT 107.875 166.155 109.625 168.450 ;
        RECT 110.265 166.155 111.075 167.155 ;
        RECT 111.715 166.155 113.465 168.450 ;
        RECT 114.105 166.155 114.915 167.155 ;
        RECT 115.555 166.155 117.305 168.450 ;
        RECT 117.945 166.155 118.755 167.155 ;
        RECT 119.395 166.155 121.145 168.450 ;
        RECT 121.785 166.155 122.595 167.155 ;
        RECT 123.235 166.155 124.985 168.450 ;
        RECT 125.625 166.155 126.435 167.155 ;
        RECT 128.805 166.155 130.555 168.940 ;
        RECT 131.195 166.155 132.005 167.155 ;
        RECT 132.645 166.155 134.395 168.450 ;
        RECT 135.035 166.155 135.845 167.155 ;
        RECT 136.485 166.155 138.235 168.450 ;
        RECT 138.875 166.155 139.685 167.155 ;
        RECT 140.325 166.155 142.075 168.450 ;
        RECT 142.715 166.155 143.525 167.155 ;
        RECT 144.165 166.155 145.915 168.450 ;
        RECT 146.555 166.155 147.365 167.155 ;
        RECT 148.005 166.155 149.755 168.450 ;
        RECT 150.395 166.155 151.205 167.155 ;
        RECT 151.845 166.155 153.595 168.450 ;
        RECT 154.235 166.155 155.045 167.155 ;
        RECT 155.685 166.155 157.435 168.450 ;
        RECT 158.075 166.155 158.885 167.155 ;
        RECT 161.300 166.345 161.670 184.855 ;
        RECT 162.320 181.220 162.690 184.855 ;
        RECT 162.315 180.840 162.695 181.220 ;
        RECT 162.320 178.220 162.690 180.840 ;
        RECT 162.315 177.840 162.695 178.220 ;
        RECT 162.320 175.220 162.690 177.840 ;
        RECT 162.315 174.840 162.695 175.220 ;
        RECT 162.320 172.220 162.690 174.840 ;
        RECT 162.315 171.840 162.695 172.220 ;
        RECT 162.320 169.220 162.690 171.840 ;
        RECT 162.315 168.840 162.695 169.220 ;
        RECT 161.300 165.965 161.680 166.345 ;
        RECT 161.300 164.895 161.670 165.965 ;
        RECT 31.925 163.705 32.735 164.705 ;
        RECT 25.090 162.265 26.780 162.495 ;
        RECT 28.150 162.365 29.610 162.595 ;
        RECT 25.090 160.255 25.690 162.265 ;
        RECT 27.110 161.805 28.110 162.130 ;
        RECT 25.920 161.245 28.780 161.575 ;
        RECT 25.090 160.025 26.780 160.255 ;
        RECT 25.090 158.015 25.690 160.025 ;
        RECT 27.495 159.890 27.760 161.245 ;
        RECT 29.010 160.355 29.610 162.365 ;
        RECT 33.375 161.875 35.125 164.705 ;
        RECT 35.765 163.705 36.575 164.705 ;
        RECT 37.215 162.410 38.965 164.705 ;
        RECT 39.605 163.705 40.415 164.705 ;
        RECT 41.055 162.410 42.805 164.705 ;
        RECT 43.445 163.705 44.255 164.705 ;
        RECT 44.895 162.410 46.645 164.705 ;
        RECT 47.285 163.705 48.095 164.705 ;
        RECT 48.735 162.410 50.485 164.705 ;
        RECT 51.125 163.705 51.935 164.705 ;
        RECT 52.575 162.410 54.325 164.705 ;
        RECT 54.965 163.705 55.775 164.705 ;
        RECT 56.415 162.410 58.165 164.705 ;
        RECT 58.805 163.705 59.615 164.705 ;
        RECT 60.255 162.410 62.005 164.705 ;
        RECT 64.375 163.705 65.185 164.705 ;
        RECT 65.825 161.875 67.575 164.705 ;
        RECT 68.215 163.705 69.025 164.705 ;
        RECT 69.665 162.410 71.415 164.705 ;
        RECT 72.055 163.705 72.865 164.705 ;
        RECT 73.505 162.410 75.255 164.705 ;
        RECT 75.895 163.705 76.705 164.705 ;
        RECT 77.345 162.410 79.095 164.705 ;
        RECT 79.735 163.705 80.545 164.705 ;
        RECT 81.185 162.410 82.935 164.705 ;
        RECT 83.575 163.705 84.385 164.705 ;
        RECT 85.025 162.410 86.775 164.705 ;
        RECT 87.415 163.705 88.225 164.705 ;
        RECT 88.865 162.410 90.615 164.705 ;
        RECT 91.255 163.705 92.065 164.705 ;
        RECT 92.705 162.410 94.455 164.705 ;
        RECT 96.825 163.705 97.635 164.705 ;
        RECT 98.275 161.875 100.025 164.705 ;
        RECT 100.665 163.705 101.475 164.705 ;
        RECT 102.115 162.410 103.865 164.705 ;
        RECT 104.505 163.705 105.315 164.705 ;
        RECT 105.955 162.410 107.705 164.705 ;
        RECT 108.345 163.705 109.155 164.705 ;
        RECT 109.795 162.410 111.545 164.705 ;
        RECT 112.185 163.705 112.995 164.705 ;
        RECT 113.635 162.410 115.385 164.705 ;
        RECT 116.025 163.705 116.835 164.705 ;
        RECT 117.475 162.410 119.225 164.705 ;
        RECT 119.865 163.705 120.675 164.705 ;
        RECT 121.315 162.410 123.065 164.705 ;
        RECT 123.705 163.705 124.515 164.705 ;
        RECT 125.155 162.410 126.905 164.705 ;
        RECT 129.275 163.705 130.085 164.705 ;
        RECT 130.725 161.875 132.475 164.705 ;
        RECT 133.115 163.705 133.925 164.705 ;
        RECT 134.565 162.410 136.315 164.705 ;
        RECT 136.955 163.705 137.765 164.705 ;
        RECT 138.405 162.410 140.155 164.705 ;
        RECT 140.795 163.705 141.605 164.705 ;
        RECT 142.245 162.410 143.995 164.705 ;
        RECT 144.635 163.705 145.445 164.705 ;
        RECT 146.085 162.410 147.835 164.705 ;
        RECT 148.475 163.705 149.285 164.705 ;
        RECT 149.925 162.410 151.675 164.705 ;
        RECT 152.315 163.705 153.125 164.705 ;
        RECT 153.765 162.410 155.515 164.705 ;
        RECT 156.155 163.705 156.965 164.705 ;
        RECT 157.605 162.410 159.355 164.705 ;
        RECT 161.300 164.515 161.680 164.895 ;
        RECT 31.650 161.505 62.170 161.875 ;
        RECT 64.100 161.505 94.620 161.875 ;
        RECT 96.550 161.505 127.070 161.875 ;
        RECT 129.000 161.505 159.520 161.875 ;
        RECT 30.800 161.240 31.420 161.425 ;
        RECT 62.400 161.240 63.020 161.425 ;
        RECT 30.800 161.010 63.020 161.240 ;
        RECT 30.800 160.825 31.420 161.010 ;
        RECT 62.400 160.825 63.020 161.010 ;
        RECT 63.250 161.240 63.870 161.425 ;
        RECT 94.850 161.240 95.470 161.425 ;
        RECT 63.250 161.010 95.470 161.240 ;
        RECT 63.250 160.825 63.870 161.010 ;
        RECT 94.850 160.825 95.470 161.010 ;
        RECT 95.700 161.240 96.320 161.425 ;
        RECT 127.300 161.240 127.920 161.425 ;
        RECT 95.700 161.010 127.920 161.240 ;
        RECT 95.700 160.825 96.320 161.010 ;
        RECT 127.300 160.825 127.920 161.010 ;
        RECT 128.150 161.240 128.770 161.425 ;
        RECT 159.750 161.240 160.370 161.425 ;
        RECT 128.150 161.010 160.370 161.240 ;
        RECT 128.150 160.825 128.770 161.010 ;
        RECT 159.750 160.825 160.370 161.010 ;
        RECT 31.650 160.375 62.170 160.755 ;
        RECT 64.100 160.375 94.620 160.755 ;
        RECT 96.550 160.375 127.070 160.755 ;
        RECT 129.000 160.375 159.520 160.755 ;
        RECT 28.150 160.125 29.610 160.355 ;
        RECT 27.110 159.565 28.110 159.890 ;
        RECT 25.920 159.005 28.780 159.335 ;
        RECT 29.010 158.115 29.610 160.125 ;
        RECT 31.650 159.665 62.170 160.035 ;
        RECT 64.100 159.665 94.620 160.035 ;
        RECT 96.550 159.665 127.070 160.035 ;
        RECT 129.000 159.665 159.520 160.035 ;
        RECT 37.280 159.655 38.900 159.665 ;
        RECT 69.730 159.655 71.350 159.665 ;
        RECT 102.180 159.655 103.800 159.665 ;
        RECT 134.630 159.655 136.250 159.665 ;
        RECT 30.800 159.400 31.420 159.585 ;
        RECT 62.400 159.400 63.020 159.585 ;
        RECT 30.800 159.170 63.020 159.400 ;
        RECT 30.800 158.985 31.420 159.170 ;
        RECT 62.400 158.985 63.020 159.170 ;
        RECT 63.250 159.400 63.870 159.585 ;
        RECT 94.850 159.400 95.470 159.585 ;
        RECT 63.250 159.170 95.470 159.400 ;
        RECT 63.250 158.985 63.870 159.170 ;
        RECT 94.850 158.985 95.470 159.170 ;
        RECT 95.700 159.400 96.320 159.585 ;
        RECT 127.300 159.400 127.920 159.585 ;
        RECT 95.700 159.170 127.920 159.400 ;
        RECT 95.700 158.985 96.320 159.170 ;
        RECT 127.300 158.985 127.920 159.170 ;
        RECT 128.150 159.400 128.770 159.585 ;
        RECT 159.750 159.400 160.370 159.585 ;
        RECT 128.150 159.170 160.370 159.400 ;
        RECT 128.150 158.985 128.770 159.170 ;
        RECT 159.750 158.985 160.370 159.170 ;
        RECT 31.650 158.535 62.170 158.915 ;
        RECT 64.100 158.535 94.620 158.915 ;
        RECT 96.550 158.535 127.070 158.915 ;
        RECT 129.000 158.535 159.520 158.915 ;
        RECT 25.090 157.785 26.780 158.015 ;
        RECT 28.150 157.885 29.610 158.115 ;
        RECT 25.090 155.730 25.690 157.785 ;
        RECT 27.110 157.325 28.110 157.650 ;
        RECT 29.010 155.730 29.610 157.885 ;
        RECT 31.650 157.820 62.170 158.190 ;
        RECT 64.100 157.820 94.620 158.190 ;
        RECT 96.550 157.820 127.070 158.190 ;
        RECT 129.000 157.820 159.520 158.190 ;
        RECT 41.120 157.810 42.740 157.820 ;
        RECT 73.570 157.810 75.190 157.820 ;
        RECT 106.020 157.810 107.640 157.820 ;
        RECT 138.470 157.810 140.090 157.820 ;
        RECT 30.800 157.555 31.420 157.740 ;
        RECT 62.400 157.555 63.020 157.740 ;
        RECT 30.800 157.325 63.020 157.555 ;
        RECT 30.800 157.140 31.420 157.325 ;
        RECT 62.400 157.140 63.020 157.325 ;
        RECT 63.250 157.555 63.870 157.740 ;
        RECT 94.850 157.555 95.470 157.740 ;
        RECT 63.250 157.325 95.470 157.555 ;
        RECT 63.250 157.140 63.870 157.325 ;
        RECT 94.850 157.140 95.470 157.325 ;
        RECT 95.700 157.555 96.320 157.740 ;
        RECT 127.300 157.555 127.920 157.740 ;
        RECT 95.700 157.325 127.920 157.555 ;
        RECT 95.700 157.140 96.320 157.325 ;
        RECT 127.300 157.140 127.920 157.325 ;
        RECT 128.150 157.555 128.770 157.740 ;
        RECT 159.750 157.555 160.370 157.740 ;
        RECT 128.150 157.325 160.370 157.555 ;
        RECT 128.150 157.140 128.770 157.325 ;
        RECT 159.750 157.140 160.370 157.325 ;
        RECT 31.650 156.690 62.170 157.070 ;
        RECT 64.100 156.690 94.620 157.070 ;
        RECT 96.550 156.690 127.070 157.070 ;
        RECT 129.000 156.690 159.520 157.070 ;
        RECT 31.660 155.900 62.160 156.340 ;
        RECT 64.110 155.900 94.610 156.340 ;
        RECT 96.560 155.900 127.060 156.340 ;
        RECT 129.010 155.900 159.510 156.340 ;
        RECT 25.090 155.390 27.380 155.730 ;
        RECT 28.125 155.390 29.610 155.730 ;
        RECT 25.090 127.545 25.690 155.390 ;
        RECT 29.010 127.545 29.610 155.390 ;
        RECT 31.650 155.180 62.170 155.550 ;
        RECT 64.100 155.180 94.620 155.550 ;
        RECT 96.550 155.180 127.070 155.550 ;
        RECT 129.000 155.180 159.520 155.550 ;
        RECT 44.960 155.170 46.580 155.180 ;
        RECT 77.410 155.170 79.030 155.180 ;
        RECT 109.860 155.170 111.480 155.180 ;
        RECT 142.310 155.170 143.930 155.180 ;
        RECT 30.800 154.915 31.420 155.100 ;
        RECT 62.400 154.915 63.020 155.100 ;
        RECT 30.800 154.685 63.020 154.915 ;
        RECT 30.800 154.500 31.420 154.685 ;
        RECT 62.400 154.500 63.020 154.685 ;
        RECT 63.250 154.915 63.870 155.100 ;
        RECT 94.850 154.915 95.470 155.100 ;
        RECT 63.250 154.685 95.470 154.915 ;
        RECT 63.250 154.500 63.870 154.685 ;
        RECT 94.850 154.500 95.470 154.685 ;
        RECT 95.700 154.915 96.320 155.100 ;
        RECT 127.300 154.915 127.920 155.100 ;
        RECT 95.700 154.685 127.920 154.915 ;
        RECT 95.700 154.500 96.320 154.685 ;
        RECT 127.300 154.500 127.920 154.685 ;
        RECT 128.150 154.915 128.770 155.100 ;
        RECT 159.750 154.915 160.370 155.100 ;
        RECT 128.150 154.685 160.370 154.915 ;
        RECT 128.150 154.500 128.770 154.685 ;
        RECT 159.750 154.500 160.370 154.685 ;
        RECT 31.650 154.050 62.170 154.430 ;
        RECT 64.100 154.050 94.620 154.430 ;
        RECT 96.550 154.050 127.070 154.430 ;
        RECT 129.000 154.050 159.520 154.430 ;
        RECT 31.650 153.340 62.170 153.710 ;
        RECT 64.100 153.340 94.620 153.710 ;
        RECT 96.550 153.340 127.070 153.710 ;
        RECT 129.000 153.340 159.520 153.710 ;
        RECT 48.800 153.330 50.420 153.340 ;
        RECT 81.250 153.330 82.870 153.340 ;
        RECT 113.700 153.330 115.320 153.340 ;
        RECT 146.150 153.330 147.770 153.340 ;
        RECT 30.800 153.075 31.420 153.260 ;
        RECT 62.400 153.075 63.020 153.260 ;
        RECT 30.800 152.845 63.020 153.075 ;
        RECT 30.800 152.660 31.420 152.845 ;
        RECT 62.400 152.660 63.020 152.845 ;
        RECT 63.250 153.075 63.870 153.260 ;
        RECT 94.850 153.075 95.470 153.260 ;
        RECT 63.250 152.845 95.470 153.075 ;
        RECT 63.250 152.660 63.870 152.845 ;
        RECT 94.850 152.660 95.470 152.845 ;
        RECT 95.700 153.075 96.320 153.260 ;
        RECT 127.300 153.075 127.920 153.260 ;
        RECT 95.700 152.845 127.920 153.075 ;
        RECT 95.700 152.660 96.320 152.845 ;
        RECT 127.300 152.660 127.920 152.845 ;
        RECT 128.150 153.075 128.770 153.260 ;
        RECT 159.750 153.075 160.370 153.260 ;
        RECT 128.150 152.845 160.370 153.075 ;
        RECT 128.150 152.660 128.770 152.845 ;
        RECT 159.750 152.660 160.370 152.845 ;
        RECT 31.650 152.210 62.170 152.590 ;
        RECT 64.100 152.210 94.620 152.590 ;
        RECT 96.550 152.210 127.070 152.590 ;
        RECT 129.000 152.210 159.520 152.590 ;
        RECT 31.650 151.495 62.170 151.865 ;
        RECT 64.100 151.495 94.620 151.865 ;
        RECT 96.550 151.495 127.070 151.865 ;
        RECT 129.000 151.495 159.520 151.865 ;
        RECT 52.640 151.485 54.260 151.495 ;
        RECT 85.090 151.485 86.710 151.495 ;
        RECT 117.540 151.485 119.160 151.495 ;
        RECT 149.990 151.485 151.610 151.495 ;
        RECT 30.800 151.230 31.420 151.415 ;
        RECT 62.400 151.230 63.020 151.415 ;
        RECT 30.800 151.000 63.020 151.230 ;
        RECT 30.800 150.815 31.420 151.000 ;
        RECT 62.400 150.815 63.020 151.000 ;
        RECT 63.250 151.230 63.870 151.415 ;
        RECT 94.850 151.230 95.470 151.415 ;
        RECT 63.250 151.000 95.470 151.230 ;
        RECT 63.250 150.815 63.870 151.000 ;
        RECT 94.850 150.815 95.470 151.000 ;
        RECT 95.700 151.230 96.320 151.415 ;
        RECT 127.300 151.230 127.920 151.415 ;
        RECT 95.700 151.000 127.920 151.230 ;
        RECT 95.700 150.815 96.320 151.000 ;
        RECT 127.300 150.815 127.920 151.000 ;
        RECT 128.150 151.230 128.770 151.415 ;
        RECT 159.750 151.230 160.370 151.415 ;
        RECT 128.150 151.000 160.370 151.230 ;
        RECT 128.150 150.815 128.770 151.000 ;
        RECT 159.750 150.815 160.370 151.000 ;
        RECT 31.650 150.365 62.170 150.745 ;
        RECT 64.100 150.365 94.620 150.745 ;
        RECT 96.550 150.365 127.070 150.745 ;
        RECT 129.000 150.365 159.520 150.745 ;
        RECT 31.660 149.575 62.160 150.015 ;
        RECT 64.110 149.575 94.610 150.015 ;
        RECT 96.560 149.575 127.060 150.015 ;
        RECT 129.010 149.575 159.510 150.015 ;
        RECT 31.650 148.855 62.170 149.225 ;
        RECT 64.100 148.855 94.620 149.225 ;
        RECT 96.550 148.855 127.070 149.225 ;
        RECT 129.000 148.855 159.520 149.225 ;
        RECT 56.480 148.845 58.100 148.855 ;
        RECT 88.930 148.845 90.550 148.855 ;
        RECT 121.380 148.845 123.000 148.855 ;
        RECT 153.830 148.845 155.450 148.855 ;
        RECT 30.800 148.590 31.420 148.775 ;
        RECT 62.400 148.590 63.020 148.775 ;
        RECT 30.800 148.360 63.020 148.590 ;
        RECT 30.800 148.175 31.420 148.360 ;
        RECT 62.400 148.175 63.020 148.360 ;
        RECT 63.250 148.590 63.870 148.775 ;
        RECT 94.850 148.590 95.470 148.775 ;
        RECT 63.250 148.360 95.470 148.590 ;
        RECT 63.250 148.175 63.870 148.360 ;
        RECT 94.850 148.175 95.470 148.360 ;
        RECT 95.700 148.590 96.320 148.775 ;
        RECT 127.300 148.590 127.920 148.775 ;
        RECT 95.700 148.360 127.920 148.590 ;
        RECT 95.700 148.175 96.320 148.360 ;
        RECT 127.300 148.175 127.920 148.360 ;
        RECT 128.150 148.590 128.770 148.775 ;
        RECT 159.750 148.590 160.370 148.775 ;
        RECT 128.150 148.360 160.370 148.590 ;
        RECT 128.150 148.175 128.770 148.360 ;
        RECT 159.750 148.175 160.370 148.360 ;
        RECT 31.650 147.725 62.170 148.105 ;
        RECT 64.100 147.725 94.620 148.105 ;
        RECT 96.550 147.725 127.070 148.105 ;
        RECT 129.000 147.725 159.520 148.105 ;
        RECT 31.650 147.015 62.170 147.385 ;
        RECT 64.100 147.015 94.620 147.385 ;
        RECT 96.550 147.015 127.070 147.385 ;
        RECT 129.000 147.015 159.520 147.385 ;
        RECT 60.320 147.005 61.940 147.015 ;
        RECT 92.770 147.005 94.390 147.015 ;
        RECT 125.220 147.005 126.840 147.015 ;
        RECT 157.670 147.005 159.290 147.015 ;
        RECT 30.800 146.750 31.420 146.935 ;
        RECT 62.400 146.750 63.020 146.935 ;
        RECT 30.800 146.520 63.020 146.750 ;
        RECT 30.800 146.335 31.420 146.520 ;
        RECT 62.400 146.335 63.020 146.520 ;
        RECT 63.250 146.750 63.870 146.935 ;
        RECT 94.850 146.750 95.470 146.935 ;
        RECT 63.250 146.520 95.470 146.750 ;
        RECT 63.250 146.335 63.870 146.520 ;
        RECT 94.850 146.335 95.470 146.520 ;
        RECT 95.700 146.750 96.320 146.935 ;
        RECT 127.300 146.750 127.920 146.935 ;
        RECT 95.700 146.520 127.920 146.750 ;
        RECT 95.700 146.335 96.320 146.520 ;
        RECT 127.300 146.335 127.920 146.520 ;
        RECT 128.150 146.750 128.770 146.935 ;
        RECT 159.750 146.750 160.370 146.935 ;
        RECT 128.150 146.520 160.370 146.750 ;
        RECT 161.300 146.585 161.670 164.515 ;
        RECT 162.320 163.220 162.690 168.840 ;
        RECT 163.340 166.345 163.710 184.855 ;
        RECT 164.360 181.220 164.730 184.855 ;
        RECT 164.355 180.840 164.735 181.220 ;
        RECT 164.360 178.220 164.730 180.840 ;
        RECT 164.355 177.840 164.735 178.220 ;
        RECT 164.360 175.220 164.730 177.840 ;
        RECT 164.355 174.840 164.735 175.220 ;
        RECT 164.360 172.220 164.730 174.840 ;
        RECT 164.355 171.840 164.735 172.220 ;
        RECT 164.360 169.220 164.730 171.840 ;
        RECT 164.355 168.840 164.735 169.220 ;
        RECT 163.340 165.965 163.720 166.345 ;
        RECT 163.340 164.895 163.710 165.965 ;
        RECT 163.340 164.515 163.720 164.895 ;
        RECT 162.315 162.840 162.695 163.220 ;
        RECT 162.320 160.220 162.690 162.840 ;
        RECT 162.315 159.840 162.695 160.220 ;
        RECT 162.320 157.220 162.690 159.840 ;
        RECT 162.315 156.840 162.695 157.220 ;
        RECT 162.320 154.220 162.690 156.840 ;
        RECT 162.315 153.840 162.695 154.220 ;
        RECT 162.320 151.220 162.690 153.840 ;
        RECT 162.315 150.840 162.695 151.220 ;
        RECT 162.320 148.220 162.690 150.840 ;
        RECT 162.315 147.840 162.695 148.220 ;
        RECT 162.320 146.585 162.690 147.840 ;
        RECT 163.340 146.585 163.710 164.515 ;
        RECT 164.360 163.220 164.730 168.840 ;
        RECT 164.355 162.840 164.735 163.220 ;
        RECT 164.360 160.220 164.730 162.840 ;
        RECT 164.355 159.840 164.735 160.220 ;
        RECT 164.360 157.220 164.730 159.840 ;
        RECT 164.355 156.840 164.735 157.220 ;
        RECT 164.360 154.220 164.730 156.840 ;
        RECT 164.355 153.840 164.735 154.220 ;
        RECT 164.360 151.220 164.730 153.840 ;
        RECT 164.355 150.840 164.735 151.220 ;
        RECT 164.360 148.220 164.730 150.840 ;
        RECT 164.355 147.840 164.735 148.220 ;
        RECT 164.360 146.585 164.730 147.840 ;
        RECT 165.380 146.585 165.760 184.855 ;
        RECT 166.110 146.595 166.550 184.845 ;
        RECT 128.150 146.335 128.770 146.520 ;
        RECT 159.750 146.335 160.370 146.520 ;
        RECT 31.650 145.885 62.170 146.265 ;
        RECT 64.100 145.885 94.620 146.265 ;
        RECT 96.550 145.885 127.070 146.265 ;
        RECT 129.000 145.885 159.520 146.265 ;
        RECT 31.650 145.165 62.170 145.545 ;
        RECT 64.100 145.165 94.620 145.545 ;
        RECT 96.550 145.165 127.070 145.545 ;
        RECT 129.000 145.165 159.520 145.545 ;
        RECT 30.800 144.910 31.420 145.095 ;
        RECT 62.400 144.910 63.020 145.095 ;
        RECT 30.800 144.680 63.020 144.910 ;
        RECT 30.800 144.495 31.420 144.680 ;
        RECT 62.400 144.495 63.020 144.680 ;
        RECT 63.250 144.910 63.870 145.095 ;
        RECT 94.850 144.910 95.470 145.095 ;
        RECT 63.250 144.680 95.470 144.910 ;
        RECT 63.250 144.495 63.870 144.680 ;
        RECT 94.850 144.495 95.470 144.680 ;
        RECT 95.700 144.910 96.320 145.095 ;
        RECT 127.300 144.910 127.920 145.095 ;
        RECT 95.700 144.680 127.920 144.910 ;
        RECT 95.700 144.495 96.320 144.680 ;
        RECT 127.300 144.495 127.920 144.680 ;
        RECT 128.150 144.910 128.770 145.095 ;
        RECT 159.750 144.910 160.370 145.095 ;
        RECT 128.150 144.680 160.370 144.910 ;
        RECT 128.150 144.495 128.770 144.680 ;
        RECT 159.750 144.495 160.370 144.680 ;
        RECT 58.400 144.415 60.020 144.425 ;
        RECT 90.850 144.415 92.470 144.425 ;
        RECT 123.300 144.415 124.920 144.425 ;
        RECT 155.750 144.415 157.370 144.425 ;
        RECT 31.650 144.045 62.170 144.415 ;
        RECT 64.100 144.045 94.620 144.415 ;
        RECT 96.550 144.045 127.070 144.415 ;
        RECT 129.000 144.045 159.520 144.415 ;
        RECT 31.650 143.325 62.170 143.705 ;
        RECT 64.100 143.325 94.620 143.705 ;
        RECT 96.550 143.325 127.070 143.705 ;
        RECT 129.000 143.325 159.520 143.705 ;
        RECT 30.800 143.070 31.420 143.255 ;
        RECT 62.400 143.070 63.020 143.255 ;
        RECT 30.800 142.840 63.020 143.070 ;
        RECT 30.800 142.655 31.420 142.840 ;
        RECT 62.400 142.655 63.020 142.840 ;
        RECT 63.250 143.070 63.870 143.255 ;
        RECT 94.850 143.070 95.470 143.255 ;
        RECT 63.250 142.840 95.470 143.070 ;
        RECT 63.250 142.655 63.870 142.840 ;
        RECT 94.850 142.655 95.470 142.840 ;
        RECT 95.700 143.070 96.320 143.255 ;
        RECT 127.300 143.070 127.920 143.255 ;
        RECT 95.700 142.840 127.920 143.070 ;
        RECT 95.700 142.655 96.320 142.840 ;
        RECT 127.300 142.655 127.920 142.840 ;
        RECT 128.150 143.070 128.770 143.255 ;
        RECT 159.750 143.070 160.370 143.255 ;
        RECT 128.150 142.840 160.370 143.070 ;
        RECT 128.150 142.655 128.770 142.840 ;
        RECT 159.750 142.655 160.370 142.840 ;
        RECT 54.560 142.575 56.180 142.585 ;
        RECT 87.010 142.575 88.630 142.585 ;
        RECT 119.460 142.575 121.080 142.585 ;
        RECT 151.910 142.575 153.530 142.585 ;
        RECT 31.650 142.205 62.170 142.575 ;
        RECT 64.100 142.205 94.620 142.575 ;
        RECT 96.550 142.205 127.070 142.575 ;
        RECT 129.000 142.205 159.520 142.575 ;
        RECT 31.660 141.410 62.160 141.850 ;
        RECT 64.110 141.410 94.610 141.850 ;
        RECT 96.560 141.410 127.060 141.850 ;
        RECT 129.010 141.410 159.510 141.850 ;
        RECT 31.650 140.680 62.170 141.060 ;
        RECT 64.100 140.680 94.620 141.060 ;
        RECT 96.550 140.680 127.070 141.060 ;
        RECT 129.000 140.680 159.520 141.060 ;
        RECT 30.800 140.425 31.420 140.610 ;
        RECT 62.400 140.425 63.020 140.610 ;
        RECT 30.800 140.195 63.020 140.425 ;
        RECT 30.800 140.010 31.420 140.195 ;
        RECT 62.400 140.010 63.020 140.195 ;
        RECT 63.250 140.425 63.870 140.610 ;
        RECT 94.850 140.425 95.470 140.610 ;
        RECT 63.250 140.195 95.470 140.425 ;
        RECT 63.250 140.010 63.870 140.195 ;
        RECT 94.850 140.010 95.470 140.195 ;
        RECT 95.700 140.425 96.320 140.610 ;
        RECT 127.300 140.425 127.920 140.610 ;
        RECT 95.700 140.195 127.920 140.425 ;
        RECT 95.700 140.010 96.320 140.195 ;
        RECT 127.300 140.010 127.920 140.195 ;
        RECT 128.150 140.425 128.770 140.610 ;
        RECT 159.750 140.425 160.370 140.610 ;
        RECT 128.150 140.195 160.370 140.425 ;
        RECT 128.150 140.010 128.770 140.195 ;
        RECT 159.750 140.010 160.370 140.195 ;
        RECT 50.720 139.930 52.340 139.940 ;
        RECT 83.170 139.930 84.790 139.940 ;
        RECT 115.620 139.930 117.240 139.940 ;
        RECT 148.070 139.930 149.690 139.940 ;
        RECT 31.650 139.560 62.170 139.930 ;
        RECT 64.100 139.560 94.620 139.930 ;
        RECT 96.550 139.560 127.070 139.930 ;
        RECT 129.000 139.560 159.520 139.930 ;
        RECT 31.650 138.840 62.170 139.220 ;
        RECT 64.100 138.840 94.620 139.220 ;
        RECT 96.550 138.840 127.070 139.220 ;
        RECT 129.000 138.840 159.520 139.220 ;
        RECT 30.800 138.585 31.420 138.770 ;
        RECT 62.400 138.585 63.020 138.770 ;
        RECT 30.800 138.355 63.020 138.585 ;
        RECT 30.800 138.170 31.420 138.355 ;
        RECT 62.400 138.170 63.020 138.355 ;
        RECT 63.250 138.585 63.870 138.770 ;
        RECT 94.850 138.585 95.470 138.770 ;
        RECT 63.250 138.355 95.470 138.585 ;
        RECT 63.250 138.170 63.870 138.355 ;
        RECT 94.850 138.170 95.470 138.355 ;
        RECT 95.700 138.585 96.320 138.770 ;
        RECT 127.300 138.585 127.920 138.770 ;
        RECT 95.700 138.355 127.920 138.585 ;
        RECT 95.700 138.170 96.320 138.355 ;
        RECT 127.300 138.170 127.920 138.355 ;
        RECT 128.150 138.585 128.770 138.770 ;
        RECT 159.750 138.585 160.370 138.770 ;
        RECT 128.150 138.355 160.370 138.585 ;
        RECT 128.150 138.170 128.770 138.355 ;
        RECT 159.750 138.170 160.370 138.355 ;
        RECT 46.880 138.090 48.500 138.100 ;
        RECT 79.330 138.090 80.950 138.100 ;
        RECT 111.780 138.090 113.400 138.100 ;
        RECT 144.230 138.090 145.850 138.100 ;
        RECT 31.650 137.720 62.170 138.090 ;
        RECT 64.100 137.720 94.620 138.090 ;
        RECT 96.550 137.720 127.070 138.090 ;
        RECT 129.000 137.720 159.520 138.090 ;
        RECT 31.650 137.000 62.170 137.380 ;
        RECT 64.100 137.000 94.620 137.380 ;
        RECT 96.550 137.000 127.070 137.380 ;
        RECT 129.000 137.000 159.520 137.380 ;
        RECT 30.800 136.745 31.420 136.930 ;
        RECT 62.400 136.745 63.020 136.930 ;
        RECT 30.800 136.515 63.020 136.745 ;
        RECT 30.800 136.330 31.420 136.515 ;
        RECT 62.400 136.330 63.020 136.515 ;
        RECT 63.250 136.745 63.870 136.930 ;
        RECT 94.850 136.745 95.470 136.930 ;
        RECT 63.250 136.515 95.470 136.745 ;
        RECT 63.250 136.330 63.870 136.515 ;
        RECT 94.850 136.330 95.470 136.515 ;
        RECT 95.700 136.745 96.320 136.930 ;
        RECT 127.300 136.745 127.920 136.930 ;
        RECT 95.700 136.515 127.920 136.745 ;
        RECT 95.700 136.330 96.320 136.515 ;
        RECT 127.300 136.330 127.920 136.515 ;
        RECT 128.150 136.745 128.770 136.930 ;
        RECT 159.750 136.745 160.370 136.930 ;
        RECT 128.150 136.515 160.370 136.745 ;
        RECT 128.150 136.330 128.770 136.515 ;
        RECT 159.750 136.330 160.370 136.515 ;
        RECT 43.040 136.250 44.660 136.260 ;
        RECT 75.490 136.250 77.110 136.260 ;
        RECT 107.940 136.250 109.560 136.260 ;
        RECT 140.390 136.250 142.010 136.260 ;
        RECT 31.650 135.880 62.170 136.250 ;
        RECT 64.100 135.880 94.620 136.250 ;
        RECT 96.550 135.880 127.070 136.250 ;
        RECT 129.000 135.880 159.520 136.250 ;
        RECT 31.660 135.085 62.160 135.525 ;
        RECT 64.110 135.085 94.610 135.525 ;
        RECT 96.560 135.085 127.060 135.525 ;
        RECT 129.010 135.085 159.510 135.525 ;
        RECT 31.650 134.355 62.170 134.735 ;
        RECT 64.100 134.355 94.620 134.735 ;
        RECT 96.550 134.355 127.070 134.735 ;
        RECT 129.000 134.355 159.520 134.735 ;
        RECT 30.800 134.100 31.420 134.285 ;
        RECT 62.400 134.100 63.020 134.285 ;
        RECT 30.800 133.870 63.020 134.100 ;
        RECT 30.800 133.685 31.420 133.870 ;
        RECT 62.400 133.685 63.020 133.870 ;
        RECT 63.250 134.100 63.870 134.285 ;
        RECT 94.850 134.100 95.470 134.285 ;
        RECT 63.250 133.870 95.470 134.100 ;
        RECT 63.250 133.685 63.870 133.870 ;
        RECT 94.850 133.685 95.470 133.870 ;
        RECT 95.700 134.100 96.320 134.285 ;
        RECT 127.300 134.100 127.920 134.285 ;
        RECT 95.700 133.870 127.920 134.100 ;
        RECT 95.700 133.685 96.320 133.870 ;
        RECT 127.300 133.685 127.920 133.870 ;
        RECT 128.150 134.100 128.770 134.285 ;
        RECT 159.750 134.100 160.370 134.285 ;
        RECT 128.150 133.870 160.370 134.100 ;
        RECT 128.150 133.685 128.770 133.870 ;
        RECT 159.750 133.685 160.370 133.870 ;
        RECT 39.200 133.605 40.820 133.615 ;
        RECT 71.650 133.605 73.270 133.615 ;
        RECT 104.100 133.605 105.720 133.615 ;
        RECT 136.550 133.605 138.170 133.615 ;
        RECT 31.650 133.235 62.170 133.605 ;
        RECT 64.100 133.235 94.620 133.605 ;
        RECT 96.550 133.235 127.070 133.605 ;
        RECT 129.000 133.235 159.520 133.605 ;
        RECT 31.650 132.515 62.170 132.895 ;
        RECT 64.100 132.515 94.620 132.895 ;
        RECT 96.550 132.515 127.070 132.895 ;
        RECT 129.000 132.515 159.520 132.895 ;
        RECT 30.800 132.260 31.420 132.445 ;
        RECT 62.400 132.260 63.020 132.445 ;
        RECT 30.800 132.030 63.020 132.260 ;
        RECT 30.800 131.845 31.420 132.030 ;
        RECT 62.400 131.845 63.020 132.030 ;
        RECT 63.250 132.260 63.870 132.445 ;
        RECT 94.850 132.260 95.470 132.445 ;
        RECT 63.250 132.030 95.470 132.260 ;
        RECT 63.250 131.845 63.870 132.030 ;
        RECT 94.850 131.845 95.470 132.030 ;
        RECT 95.700 132.260 96.320 132.445 ;
        RECT 127.300 132.260 127.920 132.445 ;
        RECT 95.700 132.030 127.920 132.260 ;
        RECT 95.700 131.845 96.320 132.030 ;
        RECT 127.300 131.845 127.920 132.030 ;
        RECT 128.150 132.260 128.770 132.445 ;
        RECT 159.750 132.260 160.370 132.445 ;
        RECT 128.150 132.030 160.370 132.260 ;
        RECT 128.150 131.845 128.770 132.030 ;
        RECT 159.750 131.845 160.370 132.030 ;
        RECT 35.360 131.765 36.980 131.775 ;
        RECT 67.810 131.765 69.430 131.775 ;
        RECT 100.260 131.765 101.880 131.775 ;
        RECT 132.710 131.765 134.330 131.775 ;
        RECT 31.650 131.395 62.170 131.765 ;
        RECT 64.100 131.395 94.620 131.765 ;
        RECT 96.550 131.395 127.070 131.765 ;
        RECT 129.000 131.395 159.520 131.765 ;
        RECT 31.650 130.675 62.170 131.055 ;
        RECT 64.100 130.675 94.620 131.055 ;
        RECT 96.550 130.675 127.070 131.055 ;
        RECT 129.000 130.675 159.520 131.055 ;
        RECT 30.800 130.420 31.420 130.605 ;
        RECT 62.400 130.420 63.020 130.605 ;
        RECT 30.800 130.190 63.020 130.420 ;
        RECT 30.800 130.005 31.420 130.190 ;
        RECT 62.400 130.005 63.020 130.190 ;
        RECT 63.250 130.420 63.870 130.605 ;
        RECT 94.850 130.420 95.470 130.605 ;
        RECT 63.250 130.190 95.470 130.420 ;
        RECT 63.250 130.005 63.870 130.190 ;
        RECT 94.850 130.005 95.470 130.190 ;
        RECT 95.700 130.420 96.320 130.605 ;
        RECT 127.300 130.420 127.920 130.605 ;
        RECT 95.700 130.190 127.920 130.420 ;
        RECT 95.700 130.005 96.320 130.190 ;
        RECT 127.300 130.005 127.920 130.190 ;
        RECT 128.150 130.420 128.770 130.605 ;
        RECT 159.750 130.420 160.370 130.605 ;
        RECT 128.150 130.190 160.370 130.420 ;
        RECT 128.150 130.005 128.770 130.190 ;
        RECT 159.750 130.005 160.370 130.190 ;
        RECT 31.650 129.555 62.170 129.925 ;
        RECT 64.100 129.555 94.620 129.925 ;
        RECT 96.550 129.555 127.070 129.925 ;
        RECT 129.000 129.555 159.520 129.925 ;
        RECT 25.090 127.205 27.380 127.545 ;
        RECT 28.125 127.205 29.610 127.545 ;
        RECT 25.090 126.570 25.690 127.205 ;
        RECT 25.090 126.340 26.670 126.570 ;
        RECT 25.090 124.300 25.690 126.340 ;
        RECT 27.100 126.110 27.460 126.195 ;
        RECT 25.970 125.880 27.460 126.110 ;
        RECT 25.970 125.730 26.330 125.880 ;
        RECT 25.920 125.095 26.870 125.500 ;
        RECT 25.090 124.070 26.380 124.300 ;
        RECT 25.090 123.110 25.690 124.070 ;
        RECT 26.610 123.750 26.870 125.095 ;
        RECT 27.100 124.445 27.460 125.880 ;
        RECT 27.690 124.545 28.040 125.745 ;
        RECT 28.400 125.135 28.780 126.780 ;
        RECT 27.480 123.750 27.830 123.810 ;
        RECT 28.400 123.750 28.740 124.355 ;
        RECT 26.610 123.490 28.740 123.750 ;
        RECT 27.480 123.430 27.830 123.490 ;
        RECT 29.010 123.210 29.610 127.205 ;
        RECT 31.455 126.770 33.205 129.555 ;
        RECT 33.845 126.770 34.655 127.770 ;
        RECT 35.295 126.770 37.045 129.065 ;
        RECT 37.685 126.770 38.495 127.770 ;
        RECT 39.135 126.770 40.885 129.065 ;
        RECT 41.525 126.770 42.335 127.770 ;
        RECT 42.975 126.770 44.725 129.065 ;
        RECT 45.365 126.770 46.175 127.770 ;
        RECT 46.815 126.770 48.565 129.065 ;
        RECT 49.205 126.770 50.015 127.770 ;
        RECT 50.655 126.770 52.405 129.065 ;
        RECT 53.045 126.770 53.855 127.770 ;
        RECT 54.495 126.770 56.245 129.065 ;
        RECT 56.885 126.770 57.695 127.770 ;
        RECT 58.335 126.770 60.085 129.065 ;
        RECT 60.725 126.770 61.535 127.770 ;
        RECT 63.905 126.770 65.655 129.555 ;
        RECT 66.295 126.770 67.105 127.770 ;
        RECT 67.745 126.770 69.495 129.065 ;
        RECT 70.135 126.770 70.945 127.770 ;
        RECT 71.585 126.770 73.335 129.065 ;
        RECT 73.975 126.770 74.785 127.770 ;
        RECT 75.425 126.770 77.175 129.065 ;
        RECT 77.815 126.770 78.625 127.770 ;
        RECT 79.265 126.770 81.015 129.065 ;
        RECT 81.655 126.770 82.465 127.770 ;
        RECT 83.105 126.770 84.855 129.065 ;
        RECT 85.495 126.770 86.305 127.770 ;
        RECT 86.945 126.770 88.695 129.065 ;
        RECT 89.335 126.770 90.145 127.770 ;
        RECT 90.785 126.770 92.535 129.065 ;
        RECT 93.175 126.770 93.985 127.770 ;
        RECT 96.355 126.770 98.105 129.555 ;
        RECT 98.745 126.770 99.555 127.770 ;
        RECT 100.195 126.770 101.945 129.065 ;
        RECT 102.585 126.770 103.395 127.770 ;
        RECT 104.035 126.770 105.785 129.065 ;
        RECT 106.425 126.770 107.235 127.770 ;
        RECT 107.875 126.770 109.625 129.065 ;
        RECT 110.265 126.770 111.075 127.770 ;
        RECT 111.715 126.770 113.465 129.065 ;
        RECT 114.105 126.770 114.915 127.770 ;
        RECT 115.555 126.770 117.305 129.065 ;
        RECT 117.945 126.770 118.755 127.770 ;
        RECT 119.395 126.770 121.145 129.065 ;
        RECT 121.785 126.770 122.595 127.770 ;
        RECT 123.235 126.770 124.985 129.065 ;
        RECT 125.625 126.770 126.435 127.770 ;
        RECT 128.805 126.770 130.555 129.555 ;
        RECT 131.195 126.770 132.005 127.770 ;
        RECT 132.645 126.770 134.395 129.065 ;
        RECT 135.035 126.770 135.845 127.770 ;
        RECT 136.485 126.770 138.235 129.065 ;
        RECT 138.875 126.770 139.685 127.770 ;
        RECT 140.325 126.770 142.075 129.065 ;
        RECT 142.715 126.770 143.525 127.770 ;
        RECT 144.165 126.770 145.915 129.065 ;
        RECT 146.555 126.770 147.365 127.770 ;
        RECT 148.005 126.770 149.755 129.065 ;
        RECT 150.395 126.770 151.205 127.770 ;
        RECT 151.845 126.770 153.595 129.065 ;
        RECT 154.235 126.770 155.045 127.770 ;
        RECT 155.685 126.770 157.435 129.065 ;
        RECT 158.075 126.770 158.885 127.770 ;
        RECT 161.300 126.960 161.670 145.470 ;
        RECT 162.320 141.835 162.690 145.470 ;
        RECT 162.315 141.455 162.695 141.835 ;
        RECT 162.320 138.835 162.690 141.455 ;
        RECT 162.315 138.455 162.695 138.835 ;
        RECT 162.320 135.835 162.690 138.455 ;
        RECT 162.315 135.455 162.695 135.835 ;
        RECT 162.320 132.835 162.690 135.455 ;
        RECT 162.315 132.455 162.695 132.835 ;
        RECT 162.320 129.835 162.690 132.455 ;
        RECT 162.315 129.455 162.695 129.835 ;
        RECT 161.300 126.580 161.680 126.960 ;
        RECT 161.300 125.510 161.670 126.580 ;
        RECT 31.925 124.320 32.735 125.320 ;
        RECT 25.090 122.880 26.780 123.110 ;
        RECT 28.150 122.980 29.610 123.210 ;
        RECT 25.090 120.870 25.690 122.880 ;
        RECT 27.110 122.420 28.110 122.745 ;
        RECT 25.920 121.860 28.780 122.190 ;
        RECT 25.090 120.640 26.780 120.870 ;
        RECT 25.090 118.630 25.690 120.640 ;
        RECT 27.495 120.505 27.760 121.860 ;
        RECT 29.010 120.970 29.610 122.980 ;
        RECT 33.375 122.490 35.125 125.320 ;
        RECT 35.765 124.320 36.575 125.320 ;
        RECT 37.215 123.025 38.965 125.320 ;
        RECT 39.605 124.320 40.415 125.320 ;
        RECT 41.055 123.025 42.805 125.320 ;
        RECT 43.445 124.320 44.255 125.320 ;
        RECT 44.895 123.025 46.645 125.320 ;
        RECT 47.285 124.320 48.095 125.320 ;
        RECT 48.735 123.025 50.485 125.320 ;
        RECT 51.125 124.320 51.935 125.320 ;
        RECT 52.575 123.025 54.325 125.320 ;
        RECT 54.965 124.320 55.775 125.320 ;
        RECT 56.415 123.025 58.165 125.320 ;
        RECT 58.805 124.320 59.615 125.320 ;
        RECT 60.255 123.025 62.005 125.320 ;
        RECT 64.375 124.320 65.185 125.320 ;
        RECT 65.825 122.490 67.575 125.320 ;
        RECT 68.215 124.320 69.025 125.320 ;
        RECT 69.665 123.025 71.415 125.320 ;
        RECT 72.055 124.320 72.865 125.320 ;
        RECT 73.505 123.025 75.255 125.320 ;
        RECT 75.895 124.320 76.705 125.320 ;
        RECT 77.345 123.025 79.095 125.320 ;
        RECT 79.735 124.320 80.545 125.320 ;
        RECT 81.185 123.025 82.935 125.320 ;
        RECT 83.575 124.320 84.385 125.320 ;
        RECT 85.025 123.025 86.775 125.320 ;
        RECT 87.415 124.320 88.225 125.320 ;
        RECT 88.865 123.025 90.615 125.320 ;
        RECT 91.255 124.320 92.065 125.320 ;
        RECT 92.705 123.025 94.455 125.320 ;
        RECT 96.825 124.320 97.635 125.320 ;
        RECT 98.275 122.490 100.025 125.320 ;
        RECT 100.665 124.320 101.475 125.320 ;
        RECT 102.115 123.025 103.865 125.320 ;
        RECT 104.505 124.320 105.315 125.320 ;
        RECT 105.955 123.025 107.705 125.320 ;
        RECT 108.345 124.320 109.155 125.320 ;
        RECT 109.795 123.025 111.545 125.320 ;
        RECT 112.185 124.320 112.995 125.320 ;
        RECT 113.635 123.025 115.385 125.320 ;
        RECT 116.025 124.320 116.835 125.320 ;
        RECT 117.475 123.025 119.225 125.320 ;
        RECT 119.865 124.320 120.675 125.320 ;
        RECT 121.315 123.025 123.065 125.320 ;
        RECT 123.705 124.320 124.515 125.320 ;
        RECT 125.155 123.025 126.905 125.320 ;
        RECT 129.275 124.320 130.085 125.320 ;
        RECT 130.725 122.490 132.475 125.320 ;
        RECT 133.115 124.320 133.925 125.320 ;
        RECT 134.565 123.025 136.315 125.320 ;
        RECT 136.955 124.320 137.765 125.320 ;
        RECT 138.405 123.025 140.155 125.320 ;
        RECT 140.795 124.320 141.605 125.320 ;
        RECT 142.245 123.025 143.995 125.320 ;
        RECT 144.635 124.320 145.445 125.320 ;
        RECT 146.085 123.025 147.835 125.320 ;
        RECT 148.475 124.320 149.285 125.320 ;
        RECT 149.925 123.025 151.675 125.320 ;
        RECT 152.315 124.320 153.125 125.320 ;
        RECT 153.765 123.025 155.515 125.320 ;
        RECT 156.155 124.320 156.965 125.320 ;
        RECT 157.605 123.025 159.355 125.320 ;
        RECT 161.300 125.130 161.680 125.510 ;
        RECT 31.650 122.120 62.170 122.490 ;
        RECT 64.100 122.120 94.620 122.490 ;
        RECT 96.550 122.120 127.070 122.490 ;
        RECT 129.000 122.120 159.520 122.490 ;
        RECT 30.800 121.855 31.420 122.040 ;
        RECT 62.400 121.855 63.020 122.040 ;
        RECT 30.800 121.625 63.020 121.855 ;
        RECT 30.800 121.440 31.420 121.625 ;
        RECT 62.400 121.440 63.020 121.625 ;
        RECT 63.250 121.855 63.870 122.040 ;
        RECT 94.850 121.855 95.470 122.040 ;
        RECT 63.250 121.625 95.470 121.855 ;
        RECT 63.250 121.440 63.870 121.625 ;
        RECT 94.850 121.440 95.470 121.625 ;
        RECT 95.700 121.855 96.320 122.040 ;
        RECT 127.300 121.855 127.920 122.040 ;
        RECT 95.700 121.625 127.920 121.855 ;
        RECT 95.700 121.440 96.320 121.625 ;
        RECT 127.300 121.440 127.920 121.625 ;
        RECT 128.150 121.855 128.770 122.040 ;
        RECT 159.750 121.855 160.370 122.040 ;
        RECT 128.150 121.625 160.370 121.855 ;
        RECT 128.150 121.440 128.770 121.625 ;
        RECT 159.750 121.440 160.370 121.625 ;
        RECT 31.650 120.990 62.170 121.370 ;
        RECT 64.100 120.990 94.620 121.370 ;
        RECT 96.550 120.990 127.070 121.370 ;
        RECT 129.000 120.990 159.520 121.370 ;
        RECT 28.150 120.740 29.610 120.970 ;
        RECT 27.110 120.180 28.110 120.505 ;
        RECT 25.920 119.620 28.780 119.950 ;
        RECT 29.010 118.730 29.610 120.740 ;
        RECT 31.650 120.280 62.170 120.650 ;
        RECT 64.100 120.280 94.620 120.650 ;
        RECT 96.550 120.280 127.070 120.650 ;
        RECT 129.000 120.280 159.520 120.650 ;
        RECT 37.280 120.270 38.900 120.280 ;
        RECT 69.730 120.270 71.350 120.280 ;
        RECT 102.180 120.270 103.800 120.280 ;
        RECT 134.630 120.270 136.250 120.280 ;
        RECT 30.800 120.015 31.420 120.200 ;
        RECT 62.400 120.015 63.020 120.200 ;
        RECT 30.800 119.785 63.020 120.015 ;
        RECT 30.800 119.600 31.420 119.785 ;
        RECT 62.400 119.600 63.020 119.785 ;
        RECT 63.250 120.015 63.870 120.200 ;
        RECT 94.850 120.015 95.470 120.200 ;
        RECT 63.250 119.785 95.470 120.015 ;
        RECT 63.250 119.600 63.870 119.785 ;
        RECT 94.850 119.600 95.470 119.785 ;
        RECT 95.700 120.015 96.320 120.200 ;
        RECT 127.300 120.015 127.920 120.200 ;
        RECT 95.700 119.785 127.920 120.015 ;
        RECT 95.700 119.600 96.320 119.785 ;
        RECT 127.300 119.600 127.920 119.785 ;
        RECT 128.150 120.015 128.770 120.200 ;
        RECT 159.750 120.015 160.370 120.200 ;
        RECT 128.150 119.785 160.370 120.015 ;
        RECT 128.150 119.600 128.770 119.785 ;
        RECT 159.750 119.600 160.370 119.785 ;
        RECT 31.650 119.150 62.170 119.530 ;
        RECT 64.100 119.150 94.620 119.530 ;
        RECT 96.550 119.150 127.070 119.530 ;
        RECT 129.000 119.150 159.520 119.530 ;
        RECT 25.090 118.400 26.780 118.630 ;
        RECT 28.150 118.500 29.610 118.730 ;
        RECT 25.090 116.345 25.690 118.400 ;
        RECT 27.110 117.940 28.110 118.265 ;
        RECT 29.010 116.345 29.610 118.500 ;
        RECT 31.650 118.435 62.170 118.805 ;
        RECT 64.100 118.435 94.620 118.805 ;
        RECT 96.550 118.435 127.070 118.805 ;
        RECT 129.000 118.435 159.520 118.805 ;
        RECT 41.120 118.425 42.740 118.435 ;
        RECT 73.570 118.425 75.190 118.435 ;
        RECT 106.020 118.425 107.640 118.435 ;
        RECT 138.470 118.425 140.090 118.435 ;
        RECT 30.800 118.170 31.420 118.355 ;
        RECT 62.400 118.170 63.020 118.355 ;
        RECT 30.800 117.940 63.020 118.170 ;
        RECT 30.800 117.755 31.420 117.940 ;
        RECT 62.400 117.755 63.020 117.940 ;
        RECT 63.250 118.170 63.870 118.355 ;
        RECT 94.850 118.170 95.470 118.355 ;
        RECT 63.250 117.940 95.470 118.170 ;
        RECT 63.250 117.755 63.870 117.940 ;
        RECT 94.850 117.755 95.470 117.940 ;
        RECT 95.700 118.170 96.320 118.355 ;
        RECT 127.300 118.170 127.920 118.355 ;
        RECT 95.700 117.940 127.920 118.170 ;
        RECT 95.700 117.755 96.320 117.940 ;
        RECT 127.300 117.755 127.920 117.940 ;
        RECT 128.150 118.170 128.770 118.355 ;
        RECT 159.750 118.170 160.370 118.355 ;
        RECT 128.150 117.940 160.370 118.170 ;
        RECT 128.150 117.755 128.770 117.940 ;
        RECT 159.750 117.755 160.370 117.940 ;
        RECT 31.650 117.305 62.170 117.685 ;
        RECT 64.100 117.305 94.620 117.685 ;
        RECT 96.550 117.305 127.070 117.685 ;
        RECT 129.000 117.305 159.520 117.685 ;
        RECT 31.660 116.515 62.160 116.955 ;
        RECT 64.110 116.515 94.610 116.955 ;
        RECT 96.560 116.515 127.060 116.955 ;
        RECT 129.010 116.515 159.510 116.955 ;
        RECT 25.090 116.005 27.380 116.345 ;
        RECT 28.125 116.005 29.610 116.345 ;
        RECT 25.090 88.160 25.690 116.005 ;
        RECT 29.010 88.160 29.610 116.005 ;
        RECT 31.650 115.795 62.170 116.165 ;
        RECT 64.100 115.795 94.620 116.165 ;
        RECT 96.550 115.795 127.070 116.165 ;
        RECT 129.000 115.795 159.520 116.165 ;
        RECT 44.960 115.785 46.580 115.795 ;
        RECT 77.410 115.785 79.030 115.795 ;
        RECT 109.860 115.785 111.480 115.795 ;
        RECT 142.310 115.785 143.930 115.795 ;
        RECT 30.800 115.530 31.420 115.715 ;
        RECT 62.400 115.530 63.020 115.715 ;
        RECT 30.800 115.300 63.020 115.530 ;
        RECT 30.800 115.115 31.420 115.300 ;
        RECT 62.400 115.115 63.020 115.300 ;
        RECT 63.250 115.530 63.870 115.715 ;
        RECT 94.850 115.530 95.470 115.715 ;
        RECT 63.250 115.300 95.470 115.530 ;
        RECT 63.250 115.115 63.870 115.300 ;
        RECT 94.850 115.115 95.470 115.300 ;
        RECT 95.700 115.530 96.320 115.715 ;
        RECT 127.300 115.530 127.920 115.715 ;
        RECT 95.700 115.300 127.920 115.530 ;
        RECT 95.700 115.115 96.320 115.300 ;
        RECT 127.300 115.115 127.920 115.300 ;
        RECT 128.150 115.530 128.770 115.715 ;
        RECT 159.750 115.530 160.370 115.715 ;
        RECT 128.150 115.300 160.370 115.530 ;
        RECT 128.150 115.115 128.770 115.300 ;
        RECT 159.750 115.115 160.370 115.300 ;
        RECT 31.650 114.665 62.170 115.045 ;
        RECT 64.100 114.665 94.620 115.045 ;
        RECT 96.550 114.665 127.070 115.045 ;
        RECT 129.000 114.665 159.520 115.045 ;
        RECT 31.650 113.955 62.170 114.325 ;
        RECT 64.100 113.955 94.620 114.325 ;
        RECT 96.550 113.955 127.070 114.325 ;
        RECT 129.000 113.955 159.520 114.325 ;
        RECT 48.800 113.945 50.420 113.955 ;
        RECT 81.250 113.945 82.870 113.955 ;
        RECT 113.700 113.945 115.320 113.955 ;
        RECT 146.150 113.945 147.770 113.955 ;
        RECT 30.800 113.690 31.420 113.875 ;
        RECT 62.400 113.690 63.020 113.875 ;
        RECT 30.800 113.460 63.020 113.690 ;
        RECT 30.800 113.275 31.420 113.460 ;
        RECT 62.400 113.275 63.020 113.460 ;
        RECT 63.250 113.690 63.870 113.875 ;
        RECT 94.850 113.690 95.470 113.875 ;
        RECT 63.250 113.460 95.470 113.690 ;
        RECT 63.250 113.275 63.870 113.460 ;
        RECT 94.850 113.275 95.470 113.460 ;
        RECT 95.700 113.690 96.320 113.875 ;
        RECT 127.300 113.690 127.920 113.875 ;
        RECT 95.700 113.460 127.920 113.690 ;
        RECT 95.700 113.275 96.320 113.460 ;
        RECT 127.300 113.275 127.920 113.460 ;
        RECT 128.150 113.690 128.770 113.875 ;
        RECT 159.750 113.690 160.370 113.875 ;
        RECT 128.150 113.460 160.370 113.690 ;
        RECT 128.150 113.275 128.770 113.460 ;
        RECT 159.750 113.275 160.370 113.460 ;
        RECT 31.650 112.825 62.170 113.205 ;
        RECT 64.100 112.825 94.620 113.205 ;
        RECT 96.550 112.825 127.070 113.205 ;
        RECT 129.000 112.825 159.520 113.205 ;
        RECT 31.650 112.110 62.170 112.480 ;
        RECT 64.100 112.110 94.620 112.480 ;
        RECT 96.550 112.110 127.070 112.480 ;
        RECT 129.000 112.110 159.520 112.480 ;
        RECT 52.640 112.100 54.260 112.110 ;
        RECT 85.090 112.100 86.710 112.110 ;
        RECT 117.540 112.100 119.160 112.110 ;
        RECT 149.990 112.100 151.610 112.110 ;
        RECT 30.800 111.845 31.420 112.030 ;
        RECT 62.400 111.845 63.020 112.030 ;
        RECT 30.800 111.615 63.020 111.845 ;
        RECT 30.800 111.430 31.420 111.615 ;
        RECT 62.400 111.430 63.020 111.615 ;
        RECT 63.250 111.845 63.870 112.030 ;
        RECT 94.850 111.845 95.470 112.030 ;
        RECT 63.250 111.615 95.470 111.845 ;
        RECT 63.250 111.430 63.870 111.615 ;
        RECT 94.850 111.430 95.470 111.615 ;
        RECT 95.700 111.845 96.320 112.030 ;
        RECT 127.300 111.845 127.920 112.030 ;
        RECT 95.700 111.615 127.920 111.845 ;
        RECT 95.700 111.430 96.320 111.615 ;
        RECT 127.300 111.430 127.920 111.615 ;
        RECT 128.150 111.845 128.770 112.030 ;
        RECT 159.750 111.845 160.370 112.030 ;
        RECT 128.150 111.615 160.370 111.845 ;
        RECT 128.150 111.430 128.770 111.615 ;
        RECT 159.750 111.430 160.370 111.615 ;
        RECT 31.650 110.980 62.170 111.360 ;
        RECT 64.100 110.980 94.620 111.360 ;
        RECT 96.550 110.980 127.070 111.360 ;
        RECT 129.000 110.980 159.520 111.360 ;
        RECT 31.660 110.190 62.160 110.630 ;
        RECT 64.110 110.190 94.610 110.630 ;
        RECT 96.560 110.190 127.060 110.630 ;
        RECT 129.010 110.190 159.510 110.630 ;
        RECT 31.650 109.470 62.170 109.840 ;
        RECT 64.100 109.470 94.620 109.840 ;
        RECT 96.550 109.470 127.070 109.840 ;
        RECT 129.000 109.470 159.520 109.840 ;
        RECT 56.480 109.460 58.100 109.470 ;
        RECT 88.930 109.460 90.550 109.470 ;
        RECT 121.380 109.460 123.000 109.470 ;
        RECT 153.830 109.460 155.450 109.470 ;
        RECT 30.800 109.205 31.420 109.390 ;
        RECT 62.400 109.205 63.020 109.390 ;
        RECT 30.800 108.975 63.020 109.205 ;
        RECT 30.800 108.790 31.420 108.975 ;
        RECT 62.400 108.790 63.020 108.975 ;
        RECT 63.250 109.205 63.870 109.390 ;
        RECT 94.850 109.205 95.470 109.390 ;
        RECT 63.250 108.975 95.470 109.205 ;
        RECT 63.250 108.790 63.870 108.975 ;
        RECT 94.850 108.790 95.470 108.975 ;
        RECT 95.700 109.205 96.320 109.390 ;
        RECT 127.300 109.205 127.920 109.390 ;
        RECT 95.700 108.975 127.920 109.205 ;
        RECT 95.700 108.790 96.320 108.975 ;
        RECT 127.300 108.790 127.920 108.975 ;
        RECT 128.150 109.205 128.770 109.390 ;
        RECT 159.750 109.205 160.370 109.390 ;
        RECT 128.150 108.975 160.370 109.205 ;
        RECT 128.150 108.790 128.770 108.975 ;
        RECT 159.750 108.790 160.370 108.975 ;
        RECT 31.650 108.340 62.170 108.720 ;
        RECT 64.100 108.340 94.620 108.720 ;
        RECT 96.550 108.340 127.070 108.720 ;
        RECT 129.000 108.340 159.520 108.720 ;
        RECT 31.650 107.630 62.170 108.000 ;
        RECT 64.100 107.630 94.620 108.000 ;
        RECT 96.550 107.630 127.070 108.000 ;
        RECT 129.000 107.630 159.520 108.000 ;
        RECT 60.320 107.620 61.940 107.630 ;
        RECT 92.770 107.620 94.390 107.630 ;
        RECT 125.220 107.620 126.840 107.630 ;
        RECT 157.670 107.620 159.290 107.630 ;
        RECT 30.800 107.365 31.420 107.550 ;
        RECT 62.400 107.365 63.020 107.550 ;
        RECT 30.800 107.135 63.020 107.365 ;
        RECT 30.800 106.950 31.420 107.135 ;
        RECT 62.400 106.950 63.020 107.135 ;
        RECT 63.250 107.365 63.870 107.550 ;
        RECT 94.850 107.365 95.470 107.550 ;
        RECT 63.250 107.135 95.470 107.365 ;
        RECT 63.250 106.950 63.870 107.135 ;
        RECT 94.850 106.950 95.470 107.135 ;
        RECT 95.700 107.365 96.320 107.550 ;
        RECT 127.300 107.365 127.920 107.550 ;
        RECT 95.700 107.135 127.920 107.365 ;
        RECT 95.700 106.950 96.320 107.135 ;
        RECT 127.300 106.950 127.920 107.135 ;
        RECT 128.150 107.365 128.770 107.550 ;
        RECT 159.750 107.365 160.370 107.550 ;
        RECT 128.150 107.135 160.370 107.365 ;
        RECT 161.300 107.200 161.670 125.130 ;
        RECT 162.320 123.835 162.690 129.455 ;
        RECT 163.340 126.960 163.710 145.470 ;
        RECT 164.360 141.835 164.730 145.470 ;
        RECT 164.355 141.455 164.735 141.835 ;
        RECT 164.360 138.835 164.730 141.455 ;
        RECT 164.355 138.455 164.735 138.835 ;
        RECT 164.360 135.835 164.730 138.455 ;
        RECT 164.355 135.455 164.735 135.835 ;
        RECT 164.360 132.835 164.730 135.455 ;
        RECT 164.355 132.455 164.735 132.835 ;
        RECT 164.360 129.835 164.730 132.455 ;
        RECT 164.355 129.455 164.735 129.835 ;
        RECT 163.340 126.580 163.720 126.960 ;
        RECT 163.340 125.510 163.710 126.580 ;
        RECT 163.340 125.130 163.720 125.510 ;
        RECT 162.315 123.455 162.695 123.835 ;
        RECT 162.320 120.835 162.690 123.455 ;
        RECT 162.315 120.455 162.695 120.835 ;
        RECT 162.320 117.835 162.690 120.455 ;
        RECT 162.315 117.455 162.695 117.835 ;
        RECT 162.320 114.835 162.690 117.455 ;
        RECT 162.315 114.455 162.695 114.835 ;
        RECT 162.320 111.835 162.690 114.455 ;
        RECT 162.315 111.455 162.695 111.835 ;
        RECT 162.320 108.835 162.690 111.455 ;
        RECT 162.315 108.455 162.695 108.835 ;
        RECT 162.320 107.200 162.690 108.455 ;
        RECT 163.340 107.200 163.710 125.130 ;
        RECT 164.360 123.835 164.730 129.455 ;
        RECT 164.355 123.455 164.735 123.835 ;
        RECT 164.360 120.835 164.730 123.455 ;
        RECT 164.355 120.455 164.735 120.835 ;
        RECT 164.360 117.835 164.730 120.455 ;
        RECT 164.355 117.455 164.735 117.835 ;
        RECT 164.360 114.835 164.730 117.455 ;
        RECT 164.355 114.455 164.735 114.835 ;
        RECT 164.360 111.835 164.730 114.455 ;
        RECT 164.355 111.455 164.735 111.835 ;
        RECT 164.360 108.835 164.730 111.455 ;
        RECT 164.355 108.455 164.735 108.835 ;
        RECT 164.360 107.200 164.730 108.455 ;
        RECT 165.380 107.200 165.760 145.470 ;
        RECT 166.110 107.210 166.550 145.460 ;
        RECT 128.150 106.950 128.770 107.135 ;
        RECT 159.750 106.950 160.370 107.135 ;
        RECT 31.650 106.500 62.170 106.880 ;
        RECT 64.100 106.500 94.620 106.880 ;
        RECT 96.550 106.500 127.070 106.880 ;
        RECT 129.000 106.500 159.520 106.880 ;
        RECT 31.650 105.780 62.170 106.160 ;
        RECT 64.100 105.780 94.620 106.160 ;
        RECT 96.550 105.780 127.070 106.160 ;
        RECT 129.000 105.780 159.520 106.160 ;
        RECT 30.800 105.525 31.420 105.710 ;
        RECT 62.400 105.525 63.020 105.710 ;
        RECT 30.800 105.295 63.020 105.525 ;
        RECT 30.800 105.110 31.420 105.295 ;
        RECT 62.400 105.110 63.020 105.295 ;
        RECT 63.250 105.525 63.870 105.710 ;
        RECT 94.850 105.525 95.470 105.710 ;
        RECT 63.250 105.295 95.470 105.525 ;
        RECT 63.250 105.110 63.870 105.295 ;
        RECT 94.850 105.110 95.470 105.295 ;
        RECT 95.700 105.525 96.320 105.710 ;
        RECT 127.300 105.525 127.920 105.710 ;
        RECT 95.700 105.295 127.920 105.525 ;
        RECT 95.700 105.110 96.320 105.295 ;
        RECT 127.300 105.110 127.920 105.295 ;
        RECT 128.150 105.525 128.770 105.710 ;
        RECT 159.750 105.525 160.370 105.710 ;
        RECT 128.150 105.295 160.370 105.525 ;
        RECT 128.150 105.110 128.770 105.295 ;
        RECT 159.750 105.110 160.370 105.295 ;
        RECT 58.400 105.030 60.020 105.040 ;
        RECT 90.850 105.030 92.470 105.040 ;
        RECT 123.300 105.030 124.920 105.040 ;
        RECT 155.750 105.030 157.370 105.040 ;
        RECT 31.650 104.660 62.170 105.030 ;
        RECT 64.100 104.660 94.620 105.030 ;
        RECT 96.550 104.660 127.070 105.030 ;
        RECT 129.000 104.660 159.520 105.030 ;
        RECT 31.650 103.940 62.170 104.320 ;
        RECT 64.100 103.940 94.620 104.320 ;
        RECT 96.550 103.940 127.070 104.320 ;
        RECT 129.000 103.940 159.520 104.320 ;
        RECT 30.800 103.685 31.420 103.870 ;
        RECT 62.400 103.685 63.020 103.870 ;
        RECT 30.800 103.455 63.020 103.685 ;
        RECT 30.800 103.270 31.420 103.455 ;
        RECT 62.400 103.270 63.020 103.455 ;
        RECT 63.250 103.685 63.870 103.870 ;
        RECT 94.850 103.685 95.470 103.870 ;
        RECT 63.250 103.455 95.470 103.685 ;
        RECT 63.250 103.270 63.870 103.455 ;
        RECT 94.850 103.270 95.470 103.455 ;
        RECT 95.700 103.685 96.320 103.870 ;
        RECT 127.300 103.685 127.920 103.870 ;
        RECT 95.700 103.455 127.920 103.685 ;
        RECT 95.700 103.270 96.320 103.455 ;
        RECT 127.300 103.270 127.920 103.455 ;
        RECT 128.150 103.685 128.770 103.870 ;
        RECT 159.750 103.685 160.370 103.870 ;
        RECT 128.150 103.455 160.370 103.685 ;
        RECT 128.150 103.270 128.770 103.455 ;
        RECT 159.750 103.270 160.370 103.455 ;
        RECT 54.560 103.190 56.180 103.200 ;
        RECT 87.010 103.190 88.630 103.200 ;
        RECT 119.460 103.190 121.080 103.200 ;
        RECT 151.910 103.190 153.530 103.200 ;
        RECT 31.650 102.820 62.170 103.190 ;
        RECT 64.100 102.820 94.620 103.190 ;
        RECT 96.550 102.820 127.070 103.190 ;
        RECT 129.000 102.820 159.520 103.190 ;
        RECT 31.660 102.025 62.160 102.465 ;
        RECT 64.110 102.025 94.610 102.465 ;
        RECT 96.560 102.025 127.060 102.465 ;
        RECT 129.010 102.025 159.510 102.465 ;
        RECT 31.650 101.295 62.170 101.675 ;
        RECT 64.100 101.295 94.620 101.675 ;
        RECT 96.550 101.295 127.070 101.675 ;
        RECT 129.000 101.295 159.520 101.675 ;
        RECT 30.800 101.040 31.420 101.225 ;
        RECT 62.400 101.040 63.020 101.225 ;
        RECT 30.800 100.810 63.020 101.040 ;
        RECT 30.800 100.625 31.420 100.810 ;
        RECT 62.400 100.625 63.020 100.810 ;
        RECT 63.250 101.040 63.870 101.225 ;
        RECT 94.850 101.040 95.470 101.225 ;
        RECT 63.250 100.810 95.470 101.040 ;
        RECT 63.250 100.625 63.870 100.810 ;
        RECT 94.850 100.625 95.470 100.810 ;
        RECT 95.700 101.040 96.320 101.225 ;
        RECT 127.300 101.040 127.920 101.225 ;
        RECT 95.700 100.810 127.920 101.040 ;
        RECT 95.700 100.625 96.320 100.810 ;
        RECT 127.300 100.625 127.920 100.810 ;
        RECT 128.150 101.040 128.770 101.225 ;
        RECT 159.750 101.040 160.370 101.225 ;
        RECT 128.150 100.810 160.370 101.040 ;
        RECT 128.150 100.625 128.770 100.810 ;
        RECT 159.750 100.625 160.370 100.810 ;
        RECT 50.720 100.545 52.340 100.555 ;
        RECT 83.170 100.545 84.790 100.555 ;
        RECT 115.620 100.545 117.240 100.555 ;
        RECT 148.070 100.545 149.690 100.555 ;
        RECT 31.650 100.175 62.170 100.545 ;
        RECT 64.100 100.175 94.620 100.545 ;
        RECT 96.550 100.175 127.070 100.545 ;
        RECT 129.000 100.175 159.520 100.545 ;
        RECT 31.650 99.455 62.170 99.835 ;
        RECT 64.100 99.455 94.620 99.835 ;
        RECT 96.550 99.455 127.070 99.835 ;
        RECT 129.000 99.455 159.520 99.835 ;
        RECT 30.800 99.200 31.420 99.385 ;
        RECT 62.400 99.200 63.020 99.385 ;
        RECT 30.800 98.970 63.020 99.200 ;
        RECT 30.800 98.785 31.420 98.970 ;
        RECT 62.400 98.785 63.020 98.970 ;
        RECT 63.250 99.200 63.870 99.385 ;
        RECT 94.850 99.200 95.470 99.385 ;
        RECT 63.250 98.970 95.470 99.200 ;
        RECT 63.250 98.785 63.870 98.970 ;
        RECT 94.850 98.785 95.470 98.970 ;
        RECT 95.700 99.200 96.320 99.385 ;
        RECT 127.300 99.200 127.920 99.385 ;
        RECT 95.700 98.970 127.920 99.200 ;
        RECT 95.700 98.785 96.320 98.970 ;
        RECT 127.300 98.785 127.920 98.970 ;
        RECT 128.150 99.200 128.770 99.385 ;
        RECT 159.750 99.200 160.370 99.385 ;
        RECT 128.150 98.970 160.370 99.200 ;
        RECT 128.150 98.785 128.770 98.970 ;
        RECT 159.750 98.785 160.370 98.970 ;
        RECT 46.880 98.705 48.500 98.715 ;
        RECT 79.330 98.705 80.950 98.715 ;
        RECT 111.780 98.705 113.400 98.715 ;
        RECT 144.230 98.705 145.850 98.715 ;
        RECT 31.650 98.335 62.170 98.705 ;
        RECT 64.100 98.335 94.620 98.705 ;
        RECT 96.550 98.335 127.070 98.705 ;
        RECT 129.000 98.335 159.520 98.705 ;
        RECT 31.650 97.615 62.170 97.995 ;
        RECT 64.100 97.615 94.620 97.995 ;
        RECT 96.550 97.615 127.070 97.995 ;
        RECT 129.000 97.615 159.520 97.995 ;
        RECT 30.800 97.360 31.420 97.545 ;
        RECT 62.400 97.360 63.020 97.545 ;
        RECT 30.800 97.130 63.020 97.360 ;
        RECT 30.800 96.945 31.420 97.130 ;
        RECT 62.400 96.945 63.020 97.130 ;
        RECT 63.250 97.360 63.870 97.545 ;
        RECT 94.850 97.360 95.470 97.545 ;
        RECT 63.250 97.130 95.470 97.360 ;
        RECT 63.250 96.945 63.870 97.130 ;
        RECT 94.850 96.945 95.470 97.130 ;
        RECT 95.700 97.360 96.320 97.545 ;
        RECT 127.300 97.360 127.920 97.545 ;
        RECT 95.700 97.130 127.920 97.360 ;
        RECT 95.700 96.945 96.320 97.130 ;
        RECT 127.300 96.945 127.920 97.130 ;
        RECT 128.150 97.360 128.770 97.545 ;
        RECT 159.750 97.360 160.370 97.545 ;
        RECT 128.150 97.130 160.370 97.360 ;
        RECT 128.150 96.945 128.770 97.130 ;
        RECT 159.750 96.945 160.370 97.130 ;
        RECT 43.040 96.865 44.660 96.875 ;
        RECT 75.490 96.865 77.110 96.875 ;
        RECT 107.940 96.865 109.560 96.875 ;
        RECT 140.390 96.865 142.010 96.875 ;
        RECT 31.650 96.495 62.170 96.865 ;
        RECT 64.100 96.495 94.620 96.865 ;
        RECT 96.550 96.495 127.070 96.865 ;
        RECT 129.000 96.495 159.520 96.865 ;
        RECT 31.660 95.700 62.160 96.140 ;
        RECT 64.110 95.700 94.610 96.140 ;
        RECT 96.560 95.700 127.060 96.140 ;
        RECT 129.010 95.700 159.510 96.140 ;
        RECT 31.650 94.970 62.170 95.350 ;
        RECT 64.100 94.970 94.620 95.350 ;
        RECT 96.550 94.970 127.070 95.350 ;
        RECT 129.000 94.970 159.520 95.350 ;
        RECT 30.800 94.715 31.420 94.900 ;
        RECT 62.400 94.715 63.020 94.900 ;
        RECT 30.800 94.485 63.020 94.715 ;
        RECT 30.800 94.300 31.420 94.485 ;
        RECT 62.400 94.300 63.020 94.485 ;
        RECT 63.250 94.715 63.870 94.900 ;
        RECT 94.850 94.715 95.470 94.900 ;
        RECT 63.250 94.485 95.470 94.715 ;
        RECT 63.250 94.300 63.870 94.485 ;
        RECT 94.850 94.300 95.470 94.485 ;
        RECT 95.700 94.715 96.320 94.900 ;
        RECT 127.300 94.715 127.920 94.900 ;
        RECT 95.700 94.485 127.920 94.715 ;
        RECT 95.700 94.300 96.320 94.485 ;
        RECT 127.300 94.300 127.920 94.485 ;
        RECT 128.150 94.715 128.770 94.900 ;
        RECT 159.750 94.715 160.370 94.900 ;
        RECT 128.150 94.485 160.370 94.715 ;
        RECT 128.150 94.300 128.770 94.485 ;
        RECT 159.750 94.300 160.370 94.485 ;
        RECT 39.200 94.220 40.820 94.230 ;
        RECT 71.650 94.220 73.270 94.230 ;
        RECT 104.100 94.220 105.720 94.230 ;
        RECT 136.550 94.220 138.170 94.230 ;
        RECT 31.650 93.850 62.170 94.220 ;
        RECT 64.100 93.850 94.620 94.220 ;
        RECT 96.550 93.850 127.070 94.220 ;
        RECT 129.000 93.850 159.520 94.220 ;
        RECT 31.650 93.130 62.170 93.510 ;
        RECT 64.100 93.130 94.620 93.510 ;
        RECT 96.550 93.130 127.070 93.510 ;
        RECT 129.000 93.130 159.520 93.510 ;
        RECT 30.800 92.875 31.420 93.060 ;
        RECT 62.400 92.875 63.020 93.060 ;
        RECT 30.800 92.645 63.020 92.875 ;
        RECT 30.800 92.460 31.420 92.645 ;
        RECT 62.400 92.460 63.020 92.645 ;
        RECT 63.250 92.875 63.870 93.060 ;
        RECT 94.850 92.875 95.470 93.060 ;
        RECT 63.250 92.645 95.470 92.875 ;
        RECT 63.250 92.460 63.870 92.645 ;
        RECT 94.850 92.460 95.470 92.645 ;
        RECT 95.700 92.875 96.320 93.060 ;
        RECT 127.300 92.875 127.920 93.060 ;
        RECT 95.700 92.645 127.920 92.875 ;
        RECT 95.700 92.460 96.320 92.645 ;
        RECT 127.300 92.460 127.920 92.645 ;
        RECT 128.150 92.875 128.770 93.060 ;
        RECT 159.750 92.875 160.370 93.060 ;
        RECT 128.150 92.645 160.370 92.875 ;
        RECT 128.150 92.460 128.770 92.645 ;
        RECT 159.750 92.460 160.370 92.645 ;
        RECT 35.360 92.380 36.980 92.390 ;
        RECT 67.810 92.380 69.430 92.390 ;
        RECT 100.260 92.380 101.880 92.390 ;
        RECT 132.710 92.380 134.330 92.390 ;
        RECT 31.650 92.010 62.170 92.380 ;
        RECT 64.100 92.010 94.620 92.380 ;
        RECT 96.550 92.010 127.070 92.380 ;
        RECT 129.000 92.010 159.520 92.380 ;
        RECT 31.650 91.290 62.170 91.670 ;
        RECT 64.100 91.290 94.620 91.670 ;
        RECT 96.550 91.290 127.070 91.670 ;
        RECT 129.000 91.290 159.520 91.670 ;
        RECT 30.800 91.035 31.420 91.220 ;
        RECT 62.400 91.035 63.020 91.220 ;
        RECT 30.800 90.805 63.020 91.035 ;
        RECT 30.800 90.620 31.420 90.805 ;
        RECT 62.400 90.620 63.020 90.805 ;
        RECT 63.250 91.035 63.870 91.220 ;
        RECT 94.850 91.035 95.470 91.220 ;
        RECT 63.250 90.805 95.470 91.035 ;
        RECT 63.250 90.620 63.870 90.805 ;
        RECT 94.850 90.620 95.470 90.805 ;
        RECT 95.700 91.035 96.320 91.220 ;
        RECT 127.300 91.035 127.920 91.220 ;
        RECT 95.700 90.805 127.920 91.035 ;
        RECT 95.700 90.620 96.320 90.805 ;
        RECT 127.300 90.620 127.920 90.805 ;
        RECT 128.150 91.035 128.770 91.220 ;
        RECT 159.750 91.035 160.370 91.220 ;
        RECT 128.150 90.805 160.370 91.035 ;
        RECT 128.150 90.620 128.770 90.805 ;
        RECT 159.750 90.620 160.370 90.805 ;
        RECT 31.650 90.170 62.170 90.540 ;
        RECT 64.100 90.170 94.620 90.540 ;
        RECT 96.550 90.170 127.070 90.540 ;
        RECT 129.000 90.170 159.520 90.540 ;
        RECT 25.090 87.820 27.380 88.160 ;
        RECT 28.125 87.820 29.610 88.160 ;
        RECT 25.090 87.185 25.690 87.820 ;
        RECT 25.090 86.955 26.670 87.185 ;
        RECT 25.090 84.915 25.690 86.955 ;
        RECT 27.100 86.725 27.460 86.810 ;
        RECT 25.970 86.495 27.460 86.725 ;
        RECT 25.970 86.345 26.330 86.495 ;
        RECT 25.920 85.710 26.870 86.115 ;
        RECT 25.090 84.685 26.380 84.915 ;
        RECT 25.090 83.725 25.690 84.685 ;
        RECT 26.610 84.365 26.870 85.710 ;
        RECT 27.100 85.060 27.460 86.495 ;
        RECT 27.690 85.160 28.040 86.360 ;
        RECT 28.400 85.750 28.780 87.395 ;
        RECT 27.480 84.365 27.830 84.425 ;
        RECT 28.400 84.365 28.740 84.970 ;
        RECT 26.610 84.105 28.740 84.365 ;
        RECT 27.480 84.045 27.830 84.105 ;
        RECT 29.010 83.825 29.610 87.820 ;
        RECT 31.455 87.385 33.205 90.170 ;
        RECT 33.845 87.385 34.655 88.385 ;
        RECT 35.295 87.385 37.045 89.680 ;
        RECT 37.685 87.385 38.495 88.385 ;
        RECT 39.135 87.385 40.885 89.680 ;
        RECT 41.525 87.385 42.335 88.385 ;
        RECT 42.975 87.385 44.725 89.680 ;
        RECT 45.365 87.385 46.175 88.385 ;
        RECT 46.815 87.385 48.565 89.680 ;
        RECT 49.205 87.385 50.015 88.385 ;
        RECT 50.655 87.385 52.405 89.680 ;
        RECT 53.045 87.385 53.855 88.385 ;
        RECT 54.495 87.385 56.245 89.680 ;
        RECT 56.885 87.385 57.695 88.385 ;
        RECT 58.335 87.385 60.085 89.680 ;
        RECT 60.725 87.385 61.535 88.385 ;
        RECT 63.905 87.385 65.655 90.170 ;
        RECT 66.295 87.385 67.105 88.385 ;
        RECT 67.745 87.385 69.495 89.680 ;
        RECT 70.135 87.385 70.945 88.385 ;
        RECT 71.585 87.385 73.335 89.680 ;
        RECT 73.975 87.385 74.785 88.385 ;
        RECT 75.425 87.385 77.175 89.680 ;
        RECT 77.815 87.385 78.625 88.385 ;
        RECT 79.265 87.385 81.015 89.680 ;
        RECT 81.655 87.385 82.465 88.385 ;
        RECT 83.105 87.385 84.855 89.680 ;
        RECT 85.495 87.385 86.305 88.385 ;
        RECT 86.945 87.385 88.695 89.680 ;
        RECT 89.335 87.385 90.145 88.385 ;
        RECT 90.785 87.385 92.535 89.680 ;
        RECT 93.175 87.385 93.985 88.385 ;
        RECT 96.355 87.385 98.105 90.170 ;
        RECT 98.745 87.385 99.555 88.385 ;
        RECT 100.195 87.385 101.945 89.680 ;
        RECT 102.585 87.385 103.395 88.385 ;
        RECT 104.035 87.385 105.785 89.680 ;
        RECT 106.425 87.385 107.235 88.385 ;
        RECT 107.875 87.385 109.625 89.680 ;
        RECT 110.265 87.385 111.075 88.385 ;
        RECT 111.715 87.385 113.465 89.680 ;
        RECT 114.105 87.385 114.915 88.385 ;
        RECT 115.555 87.385 117.305 89.680 ;
        RECT 117.945 87.385 118.755 88.385 ;
        RECT 119.395 87.385 121.145 89.680 ;
        RECT 121.785 87.385 122.595 88.385 ;
        RECT 123.235 87.385 124.985 89.680 ;
        RECT 125.625 87.385 126.435 88.385 ;
        RECT 128.805 87.385 130.555 90.170 ;
        RECT 131.195 87.385 132.005 88.385 ;
        RECT 132.645 87.385 134.395 89.680 ;
        RECT 135.035 87.385 135.845 88.385 ;
        RECT 136.485 87.385 138.235 89.680 ;
        RECT 138.875 87.385 139.685 88.385 ;
        RECT 140.325 87.385 142.075 89.680 ;
        RECT 142.715 87.385 143.525 88.385 ;
        RECT 144.165 87.385 145.915 89.680 ;
        RECT 146.555 87.385 147.365 88.385 ;
        RECT 148.005 87.385 149.755 89.680 ;
        RECT 150.395 87.385 151.205 88.385 ;
        RECT 151.845 87.385 153.595 89.680 ;
        RECT 154.235 87.385 155.045 88.385 ;
        RECT 155.685 87.385 157.435 89.680 ;
        RECT 158.075 87.385 158.885 88.385 ;
        RECT 161.300 87.575 161.670 106.085 ;
        RECT 162.320 102.450 162.690 106.085 ;
        RECT 162.315 102.070 162.695 102.450 ;
        RECT 162.320 99.450 162.690 102.070 ;
        RECT 162.315 99.070 162.695 99.450 ;
        RECT 162.320 96.450 162.690 99.070 ;
        RECT 162.315 96.070 162.695 96.450 ;
        RECT 162.320 93.450 162.690 96.070 ;
        RECT 162.315 93.070 162.695 93.450 ;
        RECT 162.320 90.450 162.690 93.070 ;
        RECT 162.315 90.070 162.695 90.450 ;
        RECT 161.300 87.195 161.680 87.575 ;
        RECT 161.300 86.125 161.670 87.195 ;
        RECT 31.925 84.935 32.735 85.935 ;
        RECT 25.090 83.495 26.780 83.725 ;
        RECT 28.150 83.595 29.610 83.825 ;
        RECT 25.090 81.485 25.690 83.495 ;
        RECT 27.110 83.035 28.110 83.360 ;
        RECT 25.920 82.475 28.780 82.805 ;
        RECT 25.090 81.255 26.780 81.485 ;
        RECT 25.090 79.245 25.690 81.255 ;
        RECT 27.495 81.120 27.760 82.475 ;
        RECT 29.010 81.585 29.610 83.595 ;
        RECT 33.375 83.105 35.125 85.935 ;
        RECT 35.765 84.935 36.575 85.935 ;
        RECT 37.215 83.640 38.965 85.935 ;
        RECT 39.605 84.935 40.415 85.935 ;
        RECT 41.055 83.640 42.805 85.935 ;
        RECT 43.445 84.935 44.255 85.935 ;
        RECT 44.895 83.640 46.645 85.935 ;
        RECT 47.285 84.935 48.095 85.935 ;
        RECT 48.735 83.640 50.485 85.935 ;
        RECT 51.125 84.935 51.935 85.935 ;
        RECT 52.575 83.640 54.325 85.935 ;
        RECT 54.965 84.935 55.775 85.935 ;
        RECT 56.415 83.640 58.165 85.935 ;
        RECT 58.805 84.935 59.615 85.935 ;
        RECT 60.255 83.640 62.005 85.935 ;
        RECT 64.375 84.935 65.185 85.935 ;
        RECT 65.825 83.105 67.575 85.935 ;
        RECT 68.215 84.935 69.025 85.935 ;
        RECT 69.665 83.640 71.415 85.935 ;
        RECT 72.055 84.935 72.865 85.935 ;
        RECT 73.505 83.640 75.255 85.935 ;
        RECT 75.895 84.935 76.705 85.935 ;
        RECT 77.345 83.640 79.095 85.935 ;
        RECT 79.735 84.935 80.545 85.935 ;
        RECT 81.185 83.640 82.935 85.935 ;
        RECT 83.575 84.935 84.385 85.935 ;
        RECT 85.025 83.640 86.775 85.935 ;
        RECT 87.415 84.935 88.225 85.935 ;
        RECT 88.865 83.640 90.615 85.935 ;
        RECT 91.255 84.935 92.065 85.935 ;
        RECT 92.705 83.640 94.455 85.935 ;
        RECT 96.825 84.935 97.635 85.935 ;
        RECT 98.275 83.105 100.025 85.935 ;
        RECT 100.665 84.935 101.475 85.935 ;
        RECT 102.115 83.640 103.865 85.935 ;
        RECT 104.505 84.935 105.315 85.935 ;
        RECT 105.955 83.640 107.705 85.935 ;
        RECT 108.345 84.935 109.155 85.935 ;
        RECT 109.795 83.640 111.545 85.935 ;
        RECT 112.185 84.935 112.995 85.935 ;
        RECT 113.635 83.640 115.385 85.935 ;
        RECT 116.025 84.935 116.835 85.935 ;
        RECT 117.475 83.640 119.225 85.935 ;
        RECT 119.865 84.935 120.675 85.935 ;
        RECT 121.315 83.640 123.065 85.935 ;
        RECT 123.705 84.935 124.515 85.935 ;
        RECT 125.155 83.640 126.905 85.935 ;
        RECT 129.275 84.935 130.085 85.935 ;
        RECT 130.725 83.105 132.475 85.935 ;
        RECT 133.115 84.935 133.925 85.935 ;
        RECT 134.565 83.640 136.315 85.935 ;
        RECT 136.955 84.935 137.765 85.935 ;
        RECT 138.405 83.640 140.155 85.935 ;
        RECT 140.795 84.935 141.605 85.935 ;
        RECT 142.245 83.640 143.995 85.935 ;
        RECT 144.635 84.935 145.445 85.935 ;
        RECT 146.085 83.640 147.835 85.935 ;
        RECT 148.475 84.935 149.285 85.935 ;
        RECT 149.925 83.640 151.675 85.935 ;
        RECT 152.315 84.935 153.125 85.935 ;
        RECT 153.765 83.640 155.515 85.935 ;
        RECT 156.155 84.935 156.965 85.935 ;
        RECT 157.605 83.640 159.355 85.935 ;
        RECT 161.300 85.745 161.680 86.125 ;
        RECT 31.650 82.735 62.170 83.105 ;
        RECT 64.100 82.735 94.620 83.105 ;
        RECT 96.550 82.735 127.070 83.105 ;
        RECT 129.000 82.735 159.520 83.105 ;
        RECT 30.800 82.470 31.420 82.655 ;
        RECT 62.400 82.470 63.020 82.655 ;
        RECT 30.800 82.240 63.020 82.470 ;
        RECT 30.800 82.055 31.420 82.240 ;
        RECT 62.400 82.055 63.020 82.240 ;
        RECT 63.250 82.470 63.870 82.655 ;
        RECT 94.850 82.470 95.470 82.655 ;
        RECT 63.250 82.240 95.470 82.470 ;
        RECT 63.250 82.055 63.870 82.240 ;
        RECT 94.850 82.055 95.470 82.240 ;
        RECT 95.700 82.470 96.320 82.655 ;
        RECT 127.300 82.470 127.920 82.655 ;
        RECT 95.700 82.240 127.920 82.470 ;
        RECT 95.700 82.055 96.320 82.240 ;
        RECT 127.300 82.055 127.920 82.240 ;
        RECT 128.150 82.470 128.770 82.655 ;
        RECT 159.750 82.470 160.370 82.655 ;
        RECT 128.150 82.240 160.370 82.470 ;
        RECT 128.150 82.055 128.770 82.240 ;
        RECT 159.750 82.055 160.370 82.240 ;
        RECT 31.650 81.605 62.170 81.985 ;
        RECT 64.100 81.605 94.620 81.985 ;
        RECT 96.550 81.605 127.070 81.985 ;
        RECT 129.000 81.605 159.520 81.985 ;
        RECT 28.150 81.355 29.610 81.585 ;
        RECT 27.110 80.795 28.110 81.120 ;
        RECT 25.920 80.235 28.780 80.565 ;
        RECT 29.010 79.345 29.610 81.355 ;
        RECT 31.650 80.895 62.170 81.265 ;
        RECT 64.100 80.895 94.620 81.265 ;
        RECT 96.550 80.895 127.070 81.265 ;
        RECT 129.000 80.895 159.520 81.265 ;
        RECT 37.280 80.885 38.900 80.895 ;
        RECT 69.730 80.885 71.350 80.895 ;
        RECT 102.180 80.885 103.800 80.895 ;
        RECT 134.630 80.885 136.250 80.895 ;
        RECT 30.800 80.630 31.420 80.815 ;
        RECT 62.400 80.630 63.020 80.815 ;
        RECT 30.800 80.400 63.020 80.630 ;
        RECT 30.800 80.215 31.420 80.400 ;
        RECT 62.400 80.215 63.020 80.400 ;
        RECT 63.250 80.630 63.870 80.815 ;
        RECT 94.850 80.630 95.470 80.815 ;
        RECT 63.250 80.400 95.470 80.630 ;
        RECT 63.250 80.215 63.870 80.400 ;
        RECT 94.850 80.215 95.470 80.400 ;
        RECT 95.700 80.630 96.320 80.815 ;
        RECT 127.300 80.630 127.920 80.815 ;
        RECT 95.700 80.400 127.920 80.630 ;
        RECT 95.700 80.215 96.320 80.400 ;
        RECT 127.300 80.215 127.920 80.400 ;
        RECT 128.150 80.630 128.770 80.815 ;
        RECT 159.750 80.630 160.370 80.815 ;
        RECT 128.150 80.400 160.370 80.630 ;
        RECT 128.150 80.215 128.770 80.400 ;
        RECT 159.750 80.215 160.370 80.400 ;
        RECT 31.650 79.765 62.170 80.145 ;
        RECT 64.100 79.765 94.620 80.145 ;
        RECT 96.550 79.765 127.070 80.145 ;
        RECT 129.000 79.765 159.520 80.145 ;
        RECT 25.090 79.015 26.780 79.245 ;
        RECT 28.150 79.115 29.610 79.345 ;
        RECT 25.090 76.960 25.690 79.015 ;
        RECT 27.110 78.555 28.110 78.880 ;
        RECT 29.010 76.960 29.610 79.115 ;
        RECT 31.650 79.050 62.170 79.420 ;
        RECT 64.100 79.050 94.620 79.420 ;
        RECT 96.550 79.050 127.070 79.420 ;
        RECT 129.000 79.050 159.520 79.420 ;
        RECT 41.120 79.040 42.740 79.050 ;
        RECT 73.570 79.040 75.190 79.050 ;
        RECT 106.020 79.040 107.640 79.050 ;
        RECT 138.470 79.040 140.090 79.050 ;
        RECT 30.800 78.785 31.420 78.970 ;
        RECT 62.400 78.785 63.020 78.970 ;
        RECT 30.800 78.555 63.020 78.785 ;
        RECT 30.800 78.370 31.420 78.555 ;
        RECT 62.400 78.370 63.020 78.555 ;
        RECT 63.250 78.785 63.870 78.970 ;
        RECT 94.850 78.785 95.470 78.970 ;
        RECT 63.250 78.555 95.470 78.785 ;
        RECT 63.250 78.370 63.870 78.555 ;
        RECT 94.850 78.370 95.470 78.555 ;
        RECT 95.700 78.785 96.320 78.970 ;
        RECT 127.300 78.785 127.920 78.970 ;
        RECT 95.700 78.555 127.920 78.785 ;
        RECT 95.700 78.370 96.320 78.555 ;
        RECT 127.300 78.370 127.920 78.555 ;
        RECT 128.150 78.785 128.770 78.970 ;
        RECT 159.750 78.785 160.370 78.970 ;
        RECT 128.150 78.555 160.370 78.785 ;
        RECT 128.150 78.370 128.770 78.555 ;
        RECT 159.750 78.370 160.370 78.555 ;
        RECT 31.650 77.920 62.170 78.300 ;
        RECT 64.100 77.920 94.620 78.300 ;
        RECT 96.550 77.920 127.070 78.300 ;
        RECT 129.000 77.920 159.520 78.300 ;
        RECT 31.660 77.130 62.160 77.570 ;
        RECT 64.110 77.130 94.610 77.570 ;
        RECT 96.560 77.130 127.060 77.570 ;
        RECT 129.010 77.130 159.510 77.570 ;
        RECT 25.090 76.620 27.380 76.960 ;
        RECT 28.125 76.620 29.610 76.960 ;
        RECT 25.090 66.885 25.690 76.620 ;
        RECT 29.010 66.885 29.610 76.620 ;
        RECT 31.650 76.410 62.170 76.780 ;
        RECT 64.100 76.410 94.620 76.780 ;
        RECT 96.550 76.410 127.070 76.780 ;
        RECT 129.000 76.410 159.520 76.780 ;
        RECT 44.960 76.400 46.580 76.410 ;
        RECT 77.410 76.400 79.030 76.410 ;
        RECT 109.860 76.400 111.480 76.410 ;
        RECT 142.310 76.400 143.930 76.410 ;
        RECT 30.800 76.145 31.420 76.330 ;
        RECT 62.400 76.145 63.020 76.330 ;
        RECT 30.800 75.915 63.020 76.145 ;
        RECT 30.800 75.730 31.420 75.915 ;
        RECT 62.400 75.730 63.020 75.915 ;
        RECT 63.250 76.145 63.870 76.330 ;
        RECT 94.850 76.145 95.470 76.330 ;
        RECT 63.250 75.915 95.470 76.145 ;
        RECT 63.250 75.730 63.870 75.915 ;
        RECT 94.850 75.730 95.470 75.915 ;
        RECT 95.700 76.145 96.320 76.330 ;
        RECT 127.300 76.145 127.920 76.330 ;
        RECT 95.700 75.915 127.920 76.145 ;
        RECT 95.700 75.730 96.320 75.915 ;
        RECT 127.300 75.730 127.920 75.915 ;
        RECT 128.150 76.145 128.770 76.330 ;
        RECT 159.750 76.145 160.370 76.330 ;
        RECT 128.150 75.915 160.370 76.145 ;
        RECT 128.150 75.730 128.770 75.915 ;
        RECT 159.750 75.730 160.370 75.915 ;
        RECT 31.650 75.280 62.170 75.660 ;
        RECT 64.100 75.280 94.620 75.660 ;
        RECT 96.550 75.280 127.070 75.660 ;
        RECT 129.000 75.280 159.520 75.660 ;
        RECT 31.650 74.570 62.170 74.940 ;
        RECT 64.100 74.570 94.620 74.940 ;
        RECT 96.550 74.570 127.070 74.940 ;
        RECT 129.000 74.570 159.520 74.940 ;
        RECT 48.800 74.560 50.420 74.570 ;
        RECT 81.250 74.560 82.870 74.570 ;
        RECT 113.700 74.560 115.320 74.570 ;
        RECT 146.150 74.560 147.770 74.570 ;
        RECT 30.800 74.305 31.420 74.490 ;
        RECT 62.400 74.305 63.020 74.490 ;
        RECT 30.800 74.075 63.020 74.305 ;
        RECT 30.800 73.890 31.420 74.075 ;
        RECT 62.400 73.890 63.020 74.075 ;
        RECT 63.250 74.305 63.870 74.490 ;
        RECT 94.850 74.305 95.470 74.490 ;
        RECT 63.250 74.075 95.470 74.305 ;
        RECT 63.250 73.890 63.870 74.075 ;
        RECT 94.850 73.890 95.470 74.075 ;
        RECT 95.700 74.305 96.320 74.490 ;
        RECT 127.300 74.305 127.920 74.490 ;
        RECT 95.700 74.075 127.920 74.305 ;
        RECT 95.700 73.890 96.320 74.075 ;
        RECT 127.300 73.890 127.920 74.075 ;
        RECT 128.150 74.305 128.770 74.490 ;
        RECT 159.750 74.305 160.370 74.490 ;
        RECT 128.150 74.075 160.370 74.305 ;
        RECT 128.150 73.890 128.770 74.075 ;
        RECT 159.750 73.890 160.370 74.075 ;
        RECT 31.650 73.440 62.170 73.820 ;
        RECT 64.100 73.440 94.620 73.820 ;
        RECT 96.550 73.440 127.070 73.820 ;
        RECT 129.000 73.440 159.520 73.820 ;
        RECT 31.650 72.725 62.170 73.095 ;
        RECT 64.100 72.725 94.620 73.095 ;
        RECT 96.550 72.725 127.070 73.095 ;
        RECT 129.000 72.725 159.520 73.095 ;
        RECT 52.640 72.715 54.260 72.725 ;
        RECT 85.090 72.715 86.710 72.725 ;
        RECT 117.540 72.715 119.160 72.725 ;
        RECT 149.990 72.715 151.610 72.725 ;
        RECT 30.800 72.460 31.420 72.645 ;
        RECT 62.400 72.460 63.020 72.645 ;
        RECT 30.800 72.230 63.020 72.460 ;
        RECT 30.800 72.045 31.420 72.230 ;
        RECT 62.400 72.045 63.020 72.230 ;
        RECT 63.250 72.460 63.870 72.645 ;
        RECT 94.850 72.460 95.470 72.645 ;
        RECT 63.250 72.230 95.470 72.460 ;
        RECT 63.250 72.045 63.870 72.230 ;
        RECT 94.850 72.045 95.470 72.230 ;
        RECT 95.700 72.460 96.320 72.645 ;
        RECT 127.300 72.460 127.920 72.645 ;
        RECT 95.700 72.230 127.920 72.460 ;
        RECT 95.700 72.045 96.320 72.230 ;
        RECT 127.300 72.045 127.920 72.230 ;
        RECT 128.150 72.460 128.770 72.645 ;
        RECT 159.750 72.460 160.370 72.645 ;
        RECT 128.150 72.230 160.370 72.460 ;
        RECT 128.150 72.045 128.770 72.230 ;
        RECT 159.750 72.045 160.370 72.230 ;
        RECT 31.650 71.595 62.170 71.975 ;
        RECT 64.100 71.595 94.620 71.975 ;
        RECT 96.550 71.595 127.070 71.975 ;
        RECT 129.000 71.595 159.520 71.975 ;
        RECT 31.660 70.805 62.160 71.245 ;
        RECT 64.110 70.805 94.610 71.245 ;
        RECT 96.560 70.805 127.060 71.245 ;
        RECT 129.010 70.805 159.510 71.245 ;
        RECT 31.650 70.085 62.170 70.455 ;
        RECT 64.100 70.085 94.620 70.455 ;
        RECT 96.550 70.085 127.070 70.455 ;
        RECT 129.000 70.085 159.520 70.455 ;
        RECT 56.480 70.075 58.100 70.085 ;
        RECT 88.930 70.075 90.550 70.085 ;
        RECT 121.380 70.075 123.000 70.085 ;
        RECT 153.830 70.075 155.450 70.085 ;
        RECT 30.800 69.820 31.420 70.005 ;
        RECT 62.400 69.820 63.020 70.005 ;
        RECT 30.800 69.590 63.020 69.820 ;
        RECT 30.800 69.405 31.420 69.590 ;
        RECT 62.400 69.405 63.020 69.590 ;
        RECT 63.250 69.820 63.870 70.005 ;
        RECT 94.850 69.820 95.470 70.005 ;
        RECT 63.250 69.590 95.470 69.820 ;
        RECT 63.250 69.405 63.870 69.590 ;
        RECT 94.850 69.405 95.470 69.590 ;
        RECT 95.700 69.820 96.320 70.005 ;
        RECT 127.300 69.820 127.920 70.005 ;
        RECT 95.700 69.590 127.920 69.820 ;
        RECT 95.700 69.405 96.320 69.590 ;
        RECT 127.300 69.405 127.920 69.590 ;
        RECT 128.150 69.820 128.770 70.005 ;
        RECT 159.750 69.820 160.370 70.005 ;
        RECT 128.150 69.590 160.370 69.820 ;
        RECT 128.150 69.405 128.770 69.590 ;
        RECT 159.750 69.405 160.370 69.590 ;
        RECT 31.650 68.955 62.170 69.335 ;
        RECT 64.100 68.955 94.620 69.335 ;
        RECT 96.550 68.955 127.070 69.335 ;
        RECT 129.000 68.955 159.520 69.335 ;
        RECT 31.650 68.245 62.170 68.615 ;
        RECT 64.100 68.245 94.620 68.615 ;
        RECT 96.550 68.245 127.070 68.615 ;
        RECT 129.000 68.245 159.520 68.615 ;
        RECT 60.320 68.235 61.940 68.245 ;
        RECT 92.770 68.235 94.390 68.245 ;
        RECT 125.220 68.235 126.840 68.245 ;
        RECT 157.670 68.235 159.290 68.245 ;
        RECT 30.800 67.980 31.420 68.165 ;
        RECT 62.400 67.980 63.020 68.165 ;
        RECT 30.800 67.750 63.020 67.980 ;
        RECT 30.800 67.565 31.420 67.750 ;
        RECT 62.400 67.565 63.020 67.750 ;
        RECT 63.250 67.980 63.870 68.165 ;
        RECT 94.850 67.980 95.470 68.165 ;
        RECT 63.250 67.750 95.470 67.980 ;
        RECT 63.250 67.565 63.870 67.750 ;
        RECT 94.850 67.565 95.470 67.750 ;
        RECT 95.700 67.980 96.320 68.165 ;
        RECT 127.300 67.980 127.920 68.165 ;
        RECT 95.700 67.750 127.920 67.980 ;
        RECT 95.700 67.565 96.320 67.750 ;
        RECT 127.300 67.565 127.920 67.750 ;
        RECT 128.150 67.980 128.770 68.165 ;
        RECT 159.750 67.980 160.370 68.165 ;
        RECT 128.150 67.750 160.370 67.980 ;
        RECT 161.300 67.815 161.670 85.745 ;
        RECT 162.320 84.450 162.690 90.070 ;
        RECT 163.340 87.575 163.710 106.085 ;
        RECT 164.360 102.450 164.730 106.085 ;
        RECT 164.355 102.070 164.735 102.450 ;
        RECT 164.360 99.450 164.730 102.070 ;
        RECT 164.355 99.070 164.735 99.450 ;
        RECT 164.360 96.450 164.730 99.070 ;
        RECT 164.355 96.070 164.735 96.450 ;
        RECT 164.360 93.450 164.730 96.070 ;
        RECT 164.355 93.070 164.735 93.450 ;
        RECT 164.360 90.450 164.730 93.070 ;
        RECT 164.355 90.070 164.735 90.450 ;
        RECT 163.340 87.195 163.720 87.575 ;
        RECT 163.340 86.125 163.710 87.195 ;
        RECT 163.340 85.745 163.720 86.125 ;
        RECT 162.315 84.070 162.695 84.450 ;
        RECT 162.320 81.450 162.690 84.070 ;
        RECT 162.315 81.070 162.695 81.450 ;
        RECT 162.320 78.450 162.690 81.070 ;
        RECT 162.315 78.070 162.695 78.450 ;
        RECT 162.320 75.450 162.690 78.070 ;
        RECT 162.315 75.070 162.695 75.450 ;
        RECT 162.320 72.450 162.690 75.070 ;
        RECT 162.315 72.070 162.695 72.450 ;
        RECT 162.320 69.450 162.690 72.070 ;
        RECT 162.315 69.070 162.695 69.450 ;
        RECT 162.320 67.815 162.690 69.070 ;
        RECT 163.340 67.815 163.710 85.745 ;
        RECT 164.360 84.450 164.730 90.070 ;
        RECT 164.355 84.070 164.735 84.450 ;
        RECT 164.360 81.450 164.730 84.070 ;
        RECT 164.355 81.070 164.735 81.450 ;
        RECT 164.360 78.450 164.730 81.070 ;
        RECT 164.355 78.070 164.735 78.450 ;
        RECT 164.360 75.450 164.730 78.070 ;
        RECT 164.355 75.070 164.735 75.450 ;
        RECT 164.360 72.450 164.730 75.070 ;
        RECT 164.355 72.070 164.735 72.450 ;
        RECT 164.360 69.450 164.730 72.070 ;
        RECT 164.355 69.070 164.735 69.450 ;
        RECT 164.360 67.815 164.730 69.070 ;
        RECT 165.380 67.815 165.760 106.085 ;
        RECT 166.110 67.825 166.550 106.075 ;
        RECT 128.150 67.565 128.770 67.750 ;
        RECT 159.750 67.565 160.370 67.750 ;
        RECT 31.650 67.115 62.170 67.495 ;
        RECT 64.100 67.115 94.620 67.495 ;
        RECT 96.550 67.115 127.070 67.495 ;
        RECT 129.000 67.115 159.520 67.495 ;
      LAYER Metal2 ;
        RECT 31.920 381.475 34.160 381.855 ;
        RECT 64.370 381.475 66.610 381.855 ;
        RECT 96.820 381.475 99.060 381.855 ;
        RECT 129.270 381.475 131.510 381.855 ;
        RECT 62.520 380.915 62.900 381.295 ;
        RECT 94.970 380.915 95.350 381.295 ;
        RECT 127.420 380.915 127.800 381.295 ;
        RECT 159.870 380.915 160.250 381.295 ;
        RECT 25.200 379.265 25.580 379.645 ;
        RECT 29.120 379.265 29.500 379.645 ;
        RECT 31.920 379.635 34.160 380.015 ;
        RECT 31.925 377.750 34.165 378.130 ;
        RECT 31.920 376.990 34.160 377.370 ;
        RECT 25.200 376.265 25.580 376.645 ;
        RECT 29.120 376.265 29.500 376.645 ;
        RECT 31.920 375.150 34.160 375.530 ;
        RECT 25.200 373.265 25.580 373.645 ;
        RECT 29.120 373.265 29.500 373.645 ;
        RECT 31.920 373.310 34.160 373.690 ;
        RECT 31.925 371.425 34.165 371.805 ;
        RECT 31.920 370.665 34.160 371.045 ;
        RECT 25.200 370.265 25.580 370.645 ;
        RECT 29.120 370.265 29.500 370.645 ;
        RECT 31.920 368.825 34.160 369.205 ;
        RECT 25.200 367.265 25.580 367.645 ;
        RECT 29.120 367.265 29.500 367.645 ;
        RECT 31.920 366.985 34.160 367.365 ;
        RECT 25.200 364.265 25.580 364.645 ;
        RECT 29.120 364.265 29.500 364.645 ;
        RECT 35.295 364.275 37.045 368.085 ;
        RECT 39.135 364.275 40.885 369.925 ;
        RECT 42.975 364.275 44.725 372.570 ;
        RECT 46.815 364.275 48.565 374.410 ;
        RECT 50.655 364.275 52.405 376.250 ;
        RECT 54.495 364.275 56.245 378.895 ;
        RECT 58.335 364.275 60.085 380.735 ;
        RECT 64.370 379.635 66.610 380.015 ;
        RECT 62.520 379.075 62.900 379.455 ;
        RECT 64.375 377.750 66.615 378.130 ;
        RECT 64.370 376.990 66.610 377.370 ;
        RECT 62.520 376.430 62.900 376.810 ;
        RECT 64.370 375.150 66.610 375.530 ;
        RECT 62.520 374.590 62.900 374.970 ;
        RECT 64.370 373.310 66.610 373.690 ;
        RECT 62.520 372.750 62.900 373.130 ;
        RECT 64.375 371.425 66.615 371.805 ;
        RECT 64.370 370.665 66.610 371.045 ;
        RECT 62.520 370.105 62.900 370.485 ;
        RECT 64.370 368.825 66.610 369.205 ;
        RECT 62.520 368.265 62.900 368.645 ;
        RECT 64.370 366.985 66.610 367.365 ;
        RECT 62.520 366.425 62.900 366.805 ;
        RECT 67.745 364.275 69.495 368.085 ;
        RECT 71.585 364.275 73.335 369.925 ;
        RECT 75.425 364.275 77.175 372.570 ;
        RECT 79.265 364.275 81.015 374.410 ;
        RECT 83.105 364.275 84.855 376.250 ;
        RECT 86.945 364.275 88.695 378.895 ;
        RECT 90.785 364.275 92.535 380.735 ;
        RECT 96.820 379.635 99.060 380.015 ;
        RECT 94.970 379.075 95.350 379.455 ;
        RECT 96.825 377.750 99.065 378.130 ;
        RECT 96.820 376.990 99.060 377.370 ;
        RECT 94.970 376.430 95.350 376.810 ;
        RECT 96.820 375.150 99.060 375.530 ;
        RECT 94.970 374.590 95.350 374.970 ;
        RECT 96.820 373.310 99.060 373.690 ;
        RECT 94.970 372.750 95.350 373.130 ;
        RECT 96.825 371.425 99.065 371.805 ;
        RECT 96.820 370.665 99.060 371.045 ;
        RECT 94.970 370.105 95.350 370.485 ;
        RECT 96.820 368.825 99.060 369.205 ;
        RECT 94.970 368.265 95.350 368.645 ;
        RECT 96.820 366.985 99.060 367.365 ;
        RECT 94.970 366.425 95.350 366.805 ;
        RECT 100.195 364.275 101.945 368.085 ;
        RECT 104.035 364.275 105.785 369.925 ;
        RECT 107.875 364.275 109.625 372.570 ;
        RECT 111.715 364.275 113.465 374.410 ;
        RECT 115.555 364.275 117.305 376.250 ;
        RECT 119.395 364.275 121.145 378.895 ;
        RECT 123.235 364.275 124.985 380.735 ;
        RECT 129.270 379.635 131.510 380.015 ;
        RECT 127.420 379.075 127.800 379.455 ;
        RECT 129.275 377.750 131.515 378.130 ;
        RECT 129.270 376.990 131.510 377.370 ;
        RECT 127.420 376.430 127.800 376.810 ;
        RECT 129.270 375.150 131.510 375.530 ;
        RECT 127.420 374.590 127.800 374.970 ;
        RECT 129.270 373.310 131.510 373.690 ;
        RECT 127.420 372.750 127.800 373.130 ;
        RECT 129.275 371.425 131.515 371.805 ;
        RECT 129.270 370.665 131.510 371.045 ;
        RECT 127.420 370.105 127.800 370.485 ;
        RECT 129.270 368.825 131.510 369.205 ;
        RECT 127.420 368.265 127.800 368.645 ;
        RECT 129.270 366.985 131.510 367.365 ;
        RECT 127.420 366.425 127.800 366.805 ;
        RECT 132.645 364.275 134.395 368.085 ;
        RECT 136.485 364.275 138.235 369.925 ;
        RECT 140.325 364.275 142.075 372.570 ;
        RECT 144.165 364.275 145.915 374.410 ;
        RECT 148.005 364.275 149.755 376.250 ;
        RECT 151.845 364.275 153.595 378.895 ;
        RECT 155.685 364.275 157.435 380.735 ;
        RECT 159.870 379.075 160.250 379.455 ;
        RECT 162.315 377.765 162.695 378.145 ;
        RECT 164.355 377.765 164.735 378.145 ;
        RECT 166.140 377.765 166.520 378.145 ;
        RECT 159.870 376.430 160.250 376.810 ;
        RECT 159.870 374.590 160.250 374.970 ;
        RECT 162.315 374.765 162.695 375.145 ;
        RECT 164.355 374.765 164.735 375.145 ;
        RECT 166.140 374.765 166.520 375.145 ;
        RECT 159.870 372.750 160.250 373.130 ;
        RECT 162.315 371.765 162.695 372.145 ;
        RECT 164.355 371.765 164.735 372.145 ;
        RECT 166.140 371.765 166.520 372.145 ;
        RECT 159.870 370.105 160.250 370.485 ;
        RECT 162.315 368.765 162.695 369.145 ;
        RECT 164.355 368.765 164.735 369.145 ;
        RECT 166.140 368.765 166.520 369.145 ;
        RECT 159.870 368.265 160.250 368.645 ;
        RECT 159.870 366.425 160.250 366.805 ;
        RECT 162.315 365.765 162.695 366.145 ;
        RECT 164.355 365.765 164.735 366.145 ;
        RECT 166.140 365.765 166.520 366.145 ;
        RECT 34.060 363.890 34.440 364.080 ;
        RECT 37.900 363.890 38.280 364.080 ;
        RECT 41.740 363.890 42.120 364.080 ;
        RECT 45.580 363.890 45.960 364.080 ;
        RECT 49.420 363.890 49.800 364.080 ;
        RECT 53.260 363.890 53.640 364.080 ;
        RECT 57.100 363.890 57.480 364.080 ;
        RECT 60.940 363.890 61.320 364.080 ;
        RECT 66.510 363.890 66.890 364.080 ;
        RECT 70.350 363.890 70.730 364.080 ;
        RECT 74.190 363.890 74.570 364.080 ;
        RECT 78.030 363.890 78.410 364.080 ;
        RECT 81.870 363.890 82.250 364.080 ;
        RECT 85.710 363.890 86.090 364.080 ;
        RECT 89.550 363.890 89.930 364.080 ;
        RECT 93.390 363.890 93.770 364.080 ;
        RECT 98.960 363.890 99.340 364.080 ;
        RECT 102.800 363.890 103.180 364.080 ;
        RECT 106.640 363.890 107.020 364.080 ;
        RECT 110.480 363.890 110.860 364.080 ;
        RECT 114.320 363.890 114.700 364.080 ;
        RECT 118.160 363.890 118.540 364.080 ;
        RECT 122.000 363.890 122.380 364.080 ;
        RECT 125.840 363.890 126.220 364.080 ;
        RECT 131.410 363.890 131.790 364.080 ;
        RECT 135.250 363.890 135.630 364.080 ;
        RECT 139.090 363.890 139.470 364.080 ;
        RECT 142.930 363.890 143.310 364.080 ;
        RECT 146.770 363.890 147.150 364.080 ;
        RECT 150.610 363.890 150.990 364.080 ;
        RECT 154.450 363.890 154.830 364.080 ;
        RECT 158.290 363.890 158.670 364.080 ;
        RECT 28.390 363.080 166.790 363.890 ;
        RECT 25.200 361.265 25.580 361.645 ;
        RECT 28.390 361.630 29.200 363.080 ;
        RECT 161.300 362.890 161.680 363.080 ;
        RECT 163.340 362.890 163.720 363.080 ;
        RECT 165.380 362.890 165.760 363.080 ;
        RECT 161.300 361.630 161.680 361.820 ;
        RECT 163.340 361.630 163.720 361.820 ;
        RECT 165.380 361.630 165.760 361.820 ;
        RECT 28.390 360.820 166.790 361.630 ;
        RECT 32.140 360.630 32.520 360.820 ;
        RECT 35.980 360.630 36.360 360.820 ;
        RECT 39.820 360.630 40.200 360.820 ;
        RECT 43.660 360.630 44.040 360.820 ;
        RECT 47.500 360.630 47.880 360.820 ;
        RECT 51.340 360.630 51.720 360.820 ;
        RECT 55.180 360.630 55.560 360.820 ;
        RECT 59.020 360.630 59.400 360.820 ;
        RECT 64.590 360.630 64.970 360.820 ;
        RECT 68.430 360.630 68.810 360.820 ;
        RECT 72.270 360.630 72.650 360.820 ;
        RECT 76.110 360.630 76.490 360.820 ;
        RECT 79.950 360.630 80.330 360.820 ;
        RECT 83.790 360.630 84.170 360.820 ;
        RECT 87.630 360.630 88.010 360.820 ;
        RECT 91.470 360.630 91.850 360.820 ;
        RECT 97.040 360.630 97.420 360.820 ;
        RECT 100.880 360.630 101.260 360.820 ;
        RECT 104.720 360.630 105.100 360.820 ;
        RECT 108.560 360.630 108.940 360.820 ;
        RECT 112.400 360.630 112.780 360.820 ;
        RECT 116.240 360.630 116.620 360.820 ;
        RECT 120.080 360.630 120.460 360.820 ;
        RECT 123.920 360.630 124.300 360.820 ;
        RECT 129.490 360.630 129.870 360.820 ;
        RECT 133.330 360.630 133.710 360.820 ;
        RECT 137.170 360.630 137.550 360.820 ;
        RECT 141.010 360.630 141.390 360.820 ;
        RECT 144.850 360.630 145.230 360.820 ;
        RECT 148.690 360.630 149.070 360.820 ;
        RECT 152.530 360.630 152.910 360.820 ;
        RECT 156.370 360.630 156.750 360.820 ;
        RECT 25.200 358.265 25.580 358.645 ;
        RECT 27.480 355.930 27.830 360.120 ;
        RECT 25.200 355.265 25.580 355.645 ;
        RECT 28.110 354.575 28.460 358.490 ;
        RECT 29.120 358.265 29.500 358.645 ;
        RECT 31.920 357.300 34.160 357.680 ;
        RECT 37.215 356.580 38.965 360.435 ;
        RECT 29.120 355.265 29.500 355.645 ;
        RECT 31.920 355.460 34.160 355.840 ;
        RECT 41.055 354.735 42.805 360.435 ;
        RECT 27.705 354.250 28.460 354.575 ;
        RECT 28.110 354.245 28.460 354.250 ;
        RECT 31.920 353.615 34.160 353.995 ;
        RECT 31.925 352.855 34.165 353.235 ;
        RECT 25.200 352.265 25.580 352.645 ;
        RECT 29.120 352.265 29.500 352.645 ;
        RECT 44.895 352.095 46.645 360.435 ;
        RECT 31.920 350.975 34.160 351.355 ;
        RECT 48.735 350.255 50.485 360.435 ;
        RECT 25.200 349.265 25.580 349.645 ;
        RECT 29.120 349.265 29.500 349.645 ;
        RECT 31.920 349.135 34.160 349.515 ;
        RECT 52.575 348.410 54.325 360.435 ;
        RECT 31.920 347.290 34.160 347.670 ;
        RECT 25.200 346.265 25.580 346.645 ;
        RECT 29.120 346.265 29.500 346.645 ;
        RECT 31.925 346.530 34.165 346.910 ;
        RECT 56.415 345.770 58.165 360.435 ;
        RECT 31.920 344.650 34.160 345.030 ;
        RECT 60.255 343.930 62.005 360.435 ;
        RECT 62.520 357.860 62.900 358.240 ;
        RECT 64.370 357.300 66.610 357.680 ;
        RECT 69.665 356.580 71.415 360.435 ;
        RECT 62.520 356.020 62.900 356.400 ;
        RECT 64.370 355.460 66.610 355.840 ;
        RECT 73.505 354.735 75.255 360.435 ;
        RECT 62.520 354.175 62.900 354.555 ;
        RECT 64.370 353.615 66.610 353.995 ;
        RECT 64.375 352.855 66.615 353.235 ;
        RECT 77.345 352.095 79.095 360.435 ;
        RECT 62.520 351.535 62.900 351.915 ;
        RECT 64.370 350.975 66.610 351.355 ;
        RECT 81.185 350.255 82.935 360.435 ;
        RECT 62.520 349.695 62.900 350.075 ;
        RECT 64.370 349.135 66.610 349.515 ;
        RECT 85.025 348.410 86.775 360.435 ;
        RECT 62.520 347.850 62.900 348.230 ;
        RECT 64.370 347.290 66.610 347.670 ;
        RECT 64.375 346.530 66.615 346.910 ;
        RECT 88.865 345.770 90.615 360.435 ;
        RECT 62.520 345.210 62.900 345.590 ;
        RECT 64.370 344.650 66.610 345.030 ;
        RECT 92.705 343.930 94.455 360.435 ;
        RECT 94.970 357.860 95.350 358.240 ;
        RECT 96.820 357.300 99.060 357.680 ;
        RECT 102.115 356.580 103.865 360.435 ;
        RECT 94.970 356.020 95.350 356.400 ;
        RECT 96.820 355.460 99.060 355.840 ;
        RECT 105.955 354.735 107.705 360.435 ;
        RECT 94.970 354.175 95.350 354.555 ;
        RECT 96.820 353.615 99.060 353.995 ;
        RECT 96.825 352.855 99.065 353.235 ;
        RECT 109.795 352.095 111.545 360.435 ;
        RECT 94.970 351.535 95.350 351.915 ;
        RECT 96.820 350.975 99.060 351.355 ;
        RECT 113.635 350.255 115.385 360.435 ;
        RECT 94.970 349.695 95.350 350.075 ;
        RECT 96.820 349.135 99.060 349.515 ;
        RECT 117.475 348.410 119.225 360.435 ;
        RECT 94.970 347.850 95.350 348.230 ;
        RECT 96.820 347.290 99.060 347.670 ;
        RECT 96.825 346.530 99.065 346.910 ;
        RECT 121.315 345.770 123.065 360.435 ;
        RECT 94.970 345.210 95.350 345.590 ;
        RECT 96.820 344.650 99.060 345.030 ;
        RECT 125.155 343.930 126.905 360.435 ;
        RECT 127.420 357.860 127.800 358.240 ;
        RECT 129.270 357.300 131.510 357.680 ;
        RECT 134.565 356.580 136.315 360.435 ;
        RECT 127.420 356.020 127.800 356.400 ;
        RECT 129.270 355.460 131.510 355.840 ;
        RECT 138.405 354.735 140.155 360.435 ;
        RECT 127.420 354.175 127.800 354.555 ;
        RECT 129.270 353.615 131.510 353.995 ;
        RECT 129.275 352.855 131.515 353.235 ;
        RECT 142.245 352.095 143.995 360.435 ;
        RECT 127.420 351.535 127.800 351.915 ;
        RECT 129.270 350.975 131.510 351.355 ;
        RECT 146.085 350.255 147.835 360.435 ;
        RECT 127.420 349.695 127.800 350.075 ;
        RECT 129.270 349.135 131.510 349.515 ;
        RECT 149.925 348.410 151.675 360.435 ;
        RECT 127.420 347.850 127.800 348.230 ;
        RECT 129.270 347.290 131.510 347.670 ;
        RECT 129.275 346.530 131.515 346.910 ;
        RECT 153.765 345.770 155.515 360.435 ;
        RECT 127.420 345.210 127.800 345.590 ;
        RECT 129.270 344.650 131.510 345.030 ;
        RECT 157.605 343.930 159.355 360.435 ;
        RECT 162.315 359.765 162.695 360.145 ;
        RECT 164.355 359.765 164.735 360.145 ;
        RECT 166.140 359.765 166.520 360.145 ;
        RECT 159.870 357.860 160.250 358.240 ;
        RECT 162.315 356.765 162.695 357.145 ;
        RECT 164.355 356.765 164.735 357.145 ;
        RECT 166.140 356.765 166.520 357.145 ;
        RECT 159.870 356.020 160.250 356.400 ;
        RECT 159.870 354.175 160.250 354.555 ;
        RECT 162.315 353.765 162.695 354.145 ;
        RECT 164.355 353.765 164.735 354.145 ;
        RECT 166.140 353.765 166.520 354.145 ;
        RECT 159.870 351.535 160.250 351.915 ;
        RECT 162.315 350.765 162.695 351.145 ;
        RECT 164.355 350.765 164.735 351.145 ;
        RECT 166.140 350.765 166.520 351.145 ;
        RECT 159.870 349.695 160.250 350.075 ;
        RECT 159.870 347.850 160.250 348.230 ;
        RECT 162.315 347.765 162.695 348.145 ;
        RECT 164.355 347.765 164.735 348.145 ;
        RECT 166.140 347.765 166.520 348.145 ;
        RECT 159.870 345.210 160.250 345.590 ;
        RECT 162.315 344.765 162.695 345.145 ;
        RECT 164.355 344.765 164.735 345.145 ;
        RECT 166.140 344.765 166.520 345.145 ;
        RECT 25.200 343.265 25.580 343.645 ;
        RECT 29.120 343.265 29.500 343.645 ;
        RECT 62.520 343.370 62.900 343.750 ;
        RECT 94.970 343.370 95.350 343.750 ;
        RECT 127.420 343.370 127.800 343.750 ;
        RECT 159.870 343.370 160.250 343.750 ;
        RECT 31.920 342.810 34.160 343.190 ;
        RECT 64.370 342.810 66.610 343.190 ;
        RECT 96.820 342.810 99.060 343.190 ;
        RECT 129.270 342.810 131.510 343.190 ;
        RECT 31.920 342.090 34.160 342.470 ;
        RECT 64.370 342.090 66.610 342.470 ;
        RECT 96.820 342.090 99.060 342.470 ;
        RECT 129.270 342.090 131.510 342.470 ;
        RECT 62.520 341.530 62.900 341.910 ;
        RECT 94.970 341.530 95.350 341.910 ;
        RECT 127.420 341.530 127.800 341.910 ;
        RECT 159.870 341.530 160.250 341.910 ;
        RECT 25.200 339.880 25.580 340.260 ;
        RECT 29.120 339.880 29.500 340.260 ;
        RECT 31.920 340.250 34.160 340.630 ;
        RECT 31.925 338.365 34.165 338.745 ;
        RECT 31.920 337.605 34.160 337.985 ;
        RECT 25.200 336.880 25.580 337.260 ;
        RECT 29.120 336.880 29.500 337.260 ;
        RECT 31.920 335.765 34.160 336.145 ;
        RECT 25.200 333.880 25.580 334.260 ;
        RECT 29.120 333.880 29.500 334.260 ;
        RECT 31.920 333.925 34.160 334.305 ;
        RECT 31.925 332.040 34.165 332.420 ;
        RECT 31.920 331.280 34.160 331.660 ;
        RECT 25.200 330.880 25.580 331.260 ;
        RECT 29.120 330.880 29.500 331.260 ;
        RECT 31.920 329.440 34.160 329.820 ;
        RECT 25.200 327.880 25.580 328.260 ;
        RECT 29.120 327.880 29.500 328.260 ;
        RECT 31.920 327.600 34.160 327.980 ;
        RECT 25.200 324.880 25.580 325.260 ;
        RECT 29.120 324.880 29.500 325.260 ;
        RECT 35.295 324.890 37.045 328.700 ;
        RECT 39.135 324.890 40.885 330.540 ;
        RECT 42.975 324.890 44.725 333.185 ;
        RECT 46.815 324.890 48.565 335.025 ;
        RECT 50.655 324.890 52.405 336.865 ;
        RECT 54.495 324.890 56.245 339.510 ;
        RECT 58.335 324.890 60.085 341.350 ;
        RECT 64.370 340.250 66.610 340.630 ;
        RECT 62.520 339.690 62.900 340.070 ;
        RECT 64.375 338.365 66.615 338.745 ;
        RECT 64.370 337.605 66.610 337.985 ;
        RECT 62.520 337.045 62.900 337.425 ;
        RECT 64.370 335.765 66.610 336.145 ;
        RECT 62.520 335.205 62.900 335.585 ;
        RECT 64.370 333.925 66.610 334.305 ;
        RECT 62.520 333.365 62.900 333.745 ;
        RECT 64.375 332.040 66.615 332.420 ;
        RECT 64.370 331.280 66.610 331.660 ;
        RECT 62.520 330.720 62.900 331.100 ;
        RECT 64.370 329.440 66.610 329.820 ;
        RECT 62.520 328.880 62.900 329.260 ;
        RECT 64.370 327.600 66.610 327.980 ;
        RECT 62.520 327.040 62.900 327.420 ;
        RECT 67.745 324.890 69.495 328.700 ;
        RECT 71.585 324.890 73.335 330.540 ;
        RECT 75.425 324.890 77.175 333.185 ;
        RECT 79.265 324.890 81.015 335.025 ;
        RECT 83.105 324.890 84.855 336.865 ;
        RECT 86.945 324.890 88.695 339.510 ;
        RECT 90.785 324.890 92.535 341.350 ;
        RECT 96.820 340.250 99.060 340.630 ;
        RECT 94.970 339.690 95.350 340.070 ;
        RECT 96.825 338.365 99.065 338.745 ;
        RECT 96.820 337.605 99.060 337.985 ;
        RECT 94.970 337.045 95.350 337.425 ;
        RECT 96.820 335.765 99.060 336.145 ;
        RECT 94.970 335.205 95.350 335.585 ;
        RECT 96.820 333.925 99.060 334.305 ;
        RECT 94.970 333.365 95.350 333.745 ;
        RECT 96.825 332.040 99.065 332.420 ;
        RECT 96.820 331.280 99.060 331.660 ;
        RECT 94.970 330.720 95.350 331.100 ;
        RECT 96.820 329.440 99.060 329.820 ;
        RECT 94.970 328.880 95.350 329.260 ;
        RECT 96.820 327.600 99.060 327.980 ;
        RECT 94.970 327.040 95.350 327.420 ;
        RECT 100.195 324.890 101.945 328.700 ;
        RECT 104.035 324.890 105.785 330.540 ;
        RECT 107.875 324.890 109.625 333.185 ;
        RECT 111.715 324.890 113.465 335.025 ;
        RECT 115.555 324.890 117.305 336.865 ;
        RECT 119.395 324.890 121.145 339.510 ;
        RECT 123.235 324.890 124.985 341.350 ;
        RECT 129.270 340.250 131.510 340.630 ;
        RECT 127.420 339.690 127.800 340.070 ;
        RECT 129.275 338.365 131.515 338.745 ;
        RECT 129.270 337.605 131.510 337.985 ;
        RECT 127.420 337.045 127.800 337.425 ;
        RECT 129.270 335.765 131.510 336.145 ;
        RECT 127.420 335.205 127.800 335.585 ;
        RECT 129.270 333.925 131.510 334.305 ;
        RECT 127.420 333.365 127.800 333.745 ;
        RECT 129.275 332.040 131.515 332.420 ;
        RECT 129.270 331.280 131.510 331.660 ;
        RECT 127.420 330.720 127.800 331.100 ;
        RECT 129.270 329.440 131.510 329.820 ;
        RECT 127.420 328.880 127.800 329.260 ;
        RECT 129.270 327.600 131.510 327.980 ;
        RECT 127.420 327.040 127.800 327.420 ;
        RECT 132.645 324.890 134.395 328.700 ;
        RECT 136.485 324.890 138.235 330.540 ;
        RECT 140.325 324.890 142.075 333.185 ;
        RECT 144.165 324.890 145.915 335.025 ;
        RECT 148.005 324.890 149.755 336.865 ;
        RECT 151.845 324.890 153.595 339.510 ;
        RECT 155.685 324.890 157.435 341.350 ;
        RECT 159.870 339.690 160.250 340.070 ;
        RECT 162.315 338.380 162.695 338.760 ;
        RECT 164.355 338.380 164.735 338.760 ;
        RECT 166.140 338.380 166.520 338.760 ;
        RECT 159.870 337.045 160.250 337.425 ;
        RECT 159.870 335.205 160.250 335.585 ;
        RECT 162.315 335.380 162.695 335.760 ;
        RECT 164.355 335.380 164.735 335.760 ;
        RECT 166.140 335.380 166.520 335.760 ;
        RECT 159.870 333.365 160.250 333.745 ;
        RECT 162.315 332.380 162.695 332.760 ;
        RECT 164.355 332.380 164.735 332.760 ;
        RECT 166.140 332.380 166.520 332.760 ;
        RECT 159.870 330.720 160.250 331.100 ;
        RECT 162.315 329.380 162.695 329.760 ;
        RECT 164.355 329.380 164.735 329.760 ;
        RECT 166.140 329.380 166.520 329.760 ;
        RECT 159.870 328.880 160.250 329.260 ;
        RECT 159.870 327.040 160.250 327.420 ;
        RECT 162.315 326.380 162.695 326.760 ;
        RECT 164.355 326.380 164.735 326.760 ;
        RECT 166.140 326.380 166.520 326.760 ;
        RECT 34.060 324.505 34.440 324.695 ;
        RECT 37.900 324.505 38.280 324.695 ;
        RECT 41.740 324.505 42.120 324.695 ;
        RECT 45.580 324.505 45.960 324.695 ;
        RECT 49.420 324.505 49.800 324.695 ;
        RECT 53.260 324.505 53.640 324.695 ;
        RECT 57.100 324.505 57.480 324.695 ;
        RECT 60.940 324.505 61.320 324.695 ;
        RECT 66.510 324.505 66.890 324.695 ;
        RECT 70.350 324.505 70.730 324.695 ;
        RECT 74.190 324.505 74.570 324.695 ;
        RECT 78.030 324.505 78.410 324.695 ;
        RECT 81.870 324.505 82.250 324.695 ;
        RECT 85.710 324.505 86.090 324.695 ;
        RECT 89.550 324.505 89.930 324.695 ;
        RECT 93.390 324.505 93.770 324.695 ;
        RECT 98.960 324.505 99.340 324.695 ;
        RECT 102.800 324.505 103.180 324.695 ;
        RECT 106.640 324.505 107.020 324.695 ;
        RECT 110.480 324.505 110.860 324.695 ;
        RECT 114.320 324.505 114.700 324.695 ;
        RECT 118.160 324.505 118.540 324.695 ;
        RECT 122.000 324.505 122.380 324.695 ;
        RECT 125.840 324.505 126.220 324.695 ;
        RECT 131.410 324.505 131.790 324.695 ;
        RECT 135.250 324.505 135.630 324.695 ;
        RECT 139.090 324.505 139.470 324.695 ;
        RECT 142.930 324.505 143.310 324.695 ;
        RECT 146.770 324.505 147.150 324.695 ;
        RECT 150.610 324.505 150.990 324.695 ;
        RECT 154.450 324.505 154.830 324.695 ;
        RECT 158.290 324.505 158.670 324.695 ;
        RECT 28.390 323.695 166.790 324.505 ;
        RECT 25.200 321.880 25.580 322.260 ;
        RECT 28.390 322.245 29.200 323.695 ;
        RECT 161.300 323.505 161.680 323.695 ;
        RECT 163.340 323.505 163.720 323.695 ;
        RECT 165.380 323.505 165.760 323.695 ;
        RECT 161.300 322.245 161.680 322.435 ;
        RECT 163.340 322.245 163.720 322.435 ;
        RECT 165.380 322.245 165.760 322.435 ;
        RECT 28.390 321.435 166.790 322.245 ;
        RECT 32.140 321.245 32.520 321.435 ;
        RECT 35.980 321.245 36.360 321.435 ;
        RECT 39.820 321.245 40.200 321.435 ;
        RECT 43.660 321.245 44.040 321.435 ;
        RECT 47.500 321.245 47.880 321.435 ;
        RECT 51.340 321.245 51.720 321.435 ;
        RECT 55.180 321.245 55.560 321.435 ;
        RECT 59.020 321.245 59.400 321.435 ;
        RECT 64.590 321.245 64.970 321.435 ;
        RECT 68.430 321.245 68.810 321.435 ;
        RECT 72.270 321.245 72.650 321.435 ;
        RECT 76.110 321.245 76.490 321.435 ;
        RECT 79.950 321.245 80.330 321.435 ;
        RECT 83.790 321.245 84.170 321.435 ;
        RECT 87.630 321.245 88.010 321.435 ;
        RECT 91.470 321.245 91.850 321.435 ;
        RECT 97.040 321.245 97.420 321.435 ;
        RECT 100.880 321.245 101.260 321.435 ;
        RECT 104.720 321.245 105.100 321.435 ;
        RECT 108.560 321.245 108.940 321.435 ;
        RECT 112.400 321.245 112.780 321.435 ;
        RECT 116.240 321.245 116.620 321.435 ;
        RECT 120.080 321.245 120.460 321.435 ;
        RECT 123.920 321.245 124.300 321.435 ;
        RECT 129.490 321.245 129.870 321.435 ;
        RECT 133.330 321.245 133.710 321.435 ;
        RECT 137.170 321.245 137.550 321.435 ;
        RECT 141.010 321.245 141.390 321.435 ;
        RECT 144.850 321.245 145.230 321.435 ;
        RECT 148.690 321.245 149.070 321.435 ;
        RECT 152.530 321.245 152.910 321.435 ;
        RECT 156.370 321.245 156.750 321.435 ;
        RECT 25.200 318.880 25.580 319.260 ;
        RECT 27.480 316.545 27.830 320.735 ;
        RECT 25.200 315.880 25.580 316.260 ;
        RECT 28.110 315.190 28.460 319.105 ;
        RECT 29.120 318.880 29.500 319.260 ;
        RECT 31.920 317.915 34.160 318.295 ;
        RECT 37.215 317.195 38.965 321.050 ;
        RECT 29.120 315.880 29.500 316.260 ;
        RECT 31.920 316.075 34.160 316.455 ;
        RECT 41.055 315.350 42.805 321.050 ;
        RECT 27.705 314.865 28.460 315.190 ;
        RECT 28.110 314.860 28.460 314.865 ;
        RECT 31.920 314.230 34.160 314.610 ;
        RECT 31.925 313.470 34.165 313.850 ;
        RECT 25.200 312.880 25.580 313.260 ;
        RECT 29.120 312.880 29.500 313.260 ;
        RECT 44.895 312.710 46.645 321.050 ;
        RECT 31.920 311.590 34.160 311.970 ;
        RECT 48.735 310.870 50.485 321.050 ;
        RECT 25.200 309.880 25.580 310.260 ;
        RECT 29.120 309.880 29.500 310.260 ;
        RECT 31.920 309.750 34.160 310.130 ;
        RECT 52.575 309.025 54.325 321.050 ;
        RECT 31.920 307.905 34.160 308.285 ;
        RECT 25.200 306.880 25.580 307.260 ;
        RECT 29.120 306.880 29.500 307.260 ;
        RECT 31.925 307.145 34.165 307.525 ;
        RECT 56.415 306.385 58.165 321.050 ;
        RECT 31.920 305.265 34.160 305.645 ;
        RECT 60.255 304.545 62.005 321.050 ;
        RECT 62.520 318.475 62.900 318.855 ;
        RECT 64.370 317.915 66.610 318.295 ;
        RECT 69.665 317.195 71.415 321.050 ;
        RECT 62.520 316.635 62.900 317.015 ;
        RECT 64.370 316.075 66.610 316.455 ;
        RECT 73.505 315.350 75.255 321.050 ;
        RECT 62.520 314.790 62.900 315.170 ;
        RECT 64.370 314.230 66.610 314.610 ;
        RECT 64.375 313.470 66.615 313.850 ;
        RECT 77.345 312.710 79.095 321.050 ;
        RECT 62.520 312.150 62.900 312.530 ;
        RECT 64.370 311.590 66.610 311.970 ;
        RECT 81.185 310.870 82.935 321.050 ;
        RECT 62.520 310.310 62.900 310.690 ;
        RECT 64.370 309.750 66.610 310.130 ;
        RECT 85.025 309.025 86.775 321.050 ;
        RECT 62.520 308.465 62.900 308.845 ;
        RECT 64.370 307.905 66.610 308.285 ;
        RECT 64.375 307.145 66.615 307.525 ;
        RECT 88.865 306.385 90.615 321.050 ;
        RECT 62.520 305.825 62.900 306.205 ;
        RECT 64.370 305.265 66.610 305.645 ;
        RECT 92.705 304.545 94.455 321.050 ;
        RECT 94.970 318.475 95.350 318.855 ;
        RECT 96.820 317.915 99.060 318.295 ;
        RECT 102.115 317.195 103.865 321.050 ;
        RECT 94.970 316.635 95.350 317.015 ;
        RECT 96.820 316.075 99.060 316.455 ;
        RECT 105.955 315.350 107.705 321.050 ;
        RECT 94.970 314.790 95.350 315.170 ;
        RECT 96.820 314.230 99.060 314.610 ;
        RECT 96.825 313.470 99.065 313.850 ;
        RECT 109.795 312.710 111.545 321.050 ;
        RECT 94.970 312.150 95.350 312.530 ;
        RECT 96.820 311.590 99.060 311.970 ;
        RECT 113.635 310.870 115.385 321.050 ;
        RECT 94.970 310.310 95.350 310.690 ;
        RECT 96.820 309.750 99.060 310.130 ;
        RECT 117.475 309.025 119.225 321.050 ;
        RECT 94.970 308.465 95.350 308.845 ;
        RECT 96.820 307.905 99.060 308.285 ;
        RECT 96.825 307.145 99.065 307.525 ;
        RECT 121.315 306.385 123.065 321.050 ;
        RECT 94.970 305.825 95.350 306.205 ;
        RECT 96.820 305.265 99.060 305.645 ;
        RECT 125.155 304.545 126.905 321.050 ;
        RECT 127.420 318.475 127.800 318.855 ;
        RECT 129.270 317.915 131.510 318.295 ;
        RECT 134.565 317.195 136.315 321.050 ;
        RECT 127.420 316.635 127.800 317.015 ;
        RECT 129.270 316.075 131.510 316.455 ;
        RECT 138.405 315.350 140.155 321.050 ;
        RECT 127.420 314.790 127.800 315.170 ;
        RECT 129.270 314.230 131.510 314.610 ;
        RECT 129.275 313.470 131.515 313.850 ;
        RECT 142.245 312.710 143.995 321.050 ;
        RECT 127.420 312.150 127.800 312.530 ;
        RECT 129.270 311.590 131.510 311.970 ;
        RECT 146.085 310.870 147.835 321.050 ;
        RECT 127.420 310.310 127.800 310.690 ;
        RECT 129.270 309.750 131.510 310.130 ;
        RECT 149.925 309.025 151.675 321.050 ;
        RECT 127.420 308.465 127.800 308.845 ;
        RECT 129.270 307.905 131.510 308.285 ;
        RECT 129.275 307.145 131.515 307.525 ;
        RECT 153.765 306.385 155.515 321.050 ;
        RECT 127.420 305.825 127.800 306.205 ;
        RECT 129.270 305.265 131.510 305.645 ;
        RECT 157.605 304.545 159.355 321.050 ;
        RECT 162.315 320.380 162.695 320.760 ;
        RECT 164.355 320.380 164.735 320.760 ;
        RECT 166.140 320.380 166.520 320.760 ;
        RECT 159.870 318.475 160.250 318.855 ;
        RECT 162.315 317.380 162.695 317.760 ;
        RECT 164.355 317.380 164.735 317.760 ;
        RECT 166.140 317.380 166.520 317.760 ;
        RECT 159.870 316.635 160.250 317.015 ;
        RECT 159.870 314.790 160.250 315.170 ;
        RECT 162.315 314.380 162.695 314.760 ;
        RECT 164.355 314.380 164.735 314.760 ;
        RECT 166.140 314.380 166.520 314.760 ;
        RECT 159.870 312.150 160.250 312.530 ;
        RECT 162.315 311.380 162.695 311.760 ;
        RECT 164.355 311.380 164.735 311.760 ;
        RECT 166.140 311.380 166.520 311.760 ;
        RECT 159.870 310.310 160.250 310.690 ;
        RECT 159.870 308.465 160.250 308.845 ;
        RECT 162.315 308.380 162.695 308.760 ;
        RECT 164.355 308.380 164.735 308.760 ;
        RECT 166.140 308.380 166.520 308.760 ;
        RECT 159.870 305.825 160.250 306.205 ;
        RECT 162.315 305.380 162.695 305.760 ;
        RECT 164.355 305.380 164.735 305.760 ;
        RECT 166.140 305.380 166.520 305.760 ;
        RECT 25.200 303.880 25.580 304.260 ;
        RECT 29.120 303.880 29.500 304.260 ;
        RECT 62.520 303.985 62.900 304.365 ;
        RECT 94.970 303.985 95.350 304.365 ;
        RECT 127.420 303.985 127.800 304.365 ;
        RECT 159.870 303.985 160.250 304.365 ;
        RECT 31.920 303.425 34.160 303.805 ;
        RECT 64.370 303.425 66.610 303.805 ;
        RECT 96.820 303.425 99.060 303.805 ;
        RECT 129.270 303.425 131.510 303.805 ;
        RECT 31.920 302.705 34.160 303.085 ;
        RECT 64.370 302.705 66.610 303.085 ;
        RECT 96.820 302.705 99.060 303.085 ;
        RECT 129.270 302.705 131.510 303.085 ;
        RECT 62.520 302.145 62.900 302.525 ;
        RECT 94.970 302.145 95.350 302.525 ;
        RECT 127.420 302.145 127.800 302.525 ;
        RECT 159.870 302.145 160.250 302.525 ;
        RECT 25.200 300.495 25.580 300.875 ;
        RECT 29.120 300.495 29.500 300.875 ;
        RECT 31.920 300.865 34.160 301.245 ;
        RECT 31.925 298.980 34.165 299.360 ;
        RECT 31.920 298.220 34.160 298.600 ;
        RECT 25.200 297.495 25.580 297.875 ;
        RECT 29.120 297.495 29.500 297.875 ;
        RECT 31.920 296.380 34.160 296.760 ;
        RECT 25.200 294.495 25.580 294.875 ;
        RECT 29.120 294.495 29.500 294.875 ;
        RECT 31.920 294.540 34.160 294.920 ;
        RECT 31.925 292.655 34.165 293.035 ;
        RECT 31.920 291.895 34.160 292.275 ;
        RECT 25.200 291.495 25.580 291.875 ;
        RECT 29.120 291.495 29.500 291.875 ;
        RECT 31.920 290.055 34.160 290.435 ;
        RECT 25.200 288.495 25.580 288.875 ;
        RECT 29.120 288.495 29.500 288.875 ;
        RECT 31.920 288.215 34.160 288.595 ;
        RECT 25.200 285.495 25.580 285.875 ;
        RECT 29.120 285.495 29.500 285.875 ;
        RECT 35.295 285.505 37.045 289.315 ;
        RECT 39.135 285.505 40.885 291.155 ;
        RECT 42.975 285.505 44.725 293.800 ;
        RECT 46.815 285.505 48.565 295.640 ;
        RECT 50.655 285.505 52.405 297.480 ;
        RECT 54.495 285.505 56.245 300.125 ;
        RECT 58.335 285.505 60.085 301.965 ;
        RECT 64.370 300.865 66.610 301.245 ;
        RECT 62.520 300.305 62.900 300.685 ;
        RECT 64.375 298.980 66.615 299.360 ;
        RECT 64.370 298.220 66.610 298.600 ;
        RECT 62.520 297.660 62.900 298.040 ;
        RECT 64.370 296.380 66.610 296.760 ;
        RECT 62.520 295.820 62.900 296.200 ;
        RECT 64.370 294.540 66.610 294.920 ;
        RECT 62.520 293.980 62.900 294.360 ;
        RECT 64.375 292.655 66.615 293.035 ;
        RECT 64.370 291.895 66.610 292.275 ;
        RECT 62.520 291.335 62.900 291.715 ;
        RECT 64.370 290.055 66.610 290.435 ;
        RECT 62.520 289.495 62.900 289.875 ;
        RECT 64.370 288.215 66.610 288.595 ;
        RECT 62.520 287.655 62.900 288.035 ;
        RECT 67.745 285.505 69.495 289.315 ;
        RECT 71.585 285.505 73.335 291.155 ;
        RECT 75.425 285.505 77.175 293.800 ;
        RECT 79.265 285.505 81.015 295.640 ;
        RECT 83.105 285.505 84.855 297.480 ;
        RECT 86.945 285.505 88.695 300.125 ;
        RECT 90.785 285.505 92.535 301.965 ;
        RECT 96.820 300.865 99.060 301.245 ;
        RECT 94.970 300.305 95.350 300.685 ;
        RECT 96.825 298.980 99.065 299.360 ;
        RECT 96.820 298.220 99.060 298.600 ;
        RECT 94.970 297.660 95.350 298.040 ;
        RECT 96.820 296.380 99.060 296.760 ;
        RECT 94.970 295.820 95.350 296.200 ;
        RECT 96.820 294.540 99.060 294.920 ;
        RECT 94.970 293.980 95.350 294.360 ;
        RECT 96.825 292.655 99.065 293.035 ;
        RECT 96.820 291.895 99.060 292.275 ;
        RECT 94.970 291.335 95.350 291.715 ;
        RECT 96.820 290.055 99.060 290.435 ;
        RECT 94.970 289.495 95.350 289.875 ;
        RECT 96.820 288.215 99.060 288.595 ;
        RECT 94.970 287.655 95.350 288.035 ;
        RECT 100.195 285.505 101.945 289.315 ;
        RECT 104.035 285.505 105.785 291.155 ;
        RECT 107.875 285.505 109.625 293.800 ;
        RECT 111.715 285.505 113.465 295.640 ;
        RECT 115.555 285.505 117.305 297.480 ;
        RECT 119.395 285.505 121.145 300.125 ;
        RECT 123.235 285.505 124.985 301.965 ;
        RECT 129.270 300.865 131.510 301.245 ;
        RECT 127.420 300.305 127.800 300.685 ;
        RECT 129.275 298.980 131.515 299.360 ;
        RECT 129.270 298.220 131.510 298.600 ;
        RECT 127.420 297.660 127.800 298.040 ;
        RECT 129.270 296.380 131.510 296.760 ;
        RECT 127.420 295.820 127.800 296.200 ;
        RECT 129.270 294.540 131.510 294.920 ;
        RECT 127.420 293.980 127.800 294.360 ;
        RECT 129.275 292.655 131.515 293.035 ;
        RECT 129.270 291.895 131.510 292.275 ;
        RECT 127.420 291.335 127.800 291.715 ;
        RECT 129.270 290.055 131.510 290.435 ;
        RECT 127.420 289.495 127.800 289.875 ;
        RECT 129.270 288.215 131.510 288.595 ;
        RECT 127.420 287.655 127.800 288.035 ;
        RECT 132.645 285.505 134.395 289.315 ;
        RECT 136.485 285.505 138.235 291.155 ;
        RECT 140.325 285.505 142.075 293.800 ;
        RECT 144.165 285.505 145.915 295.640 ;
        RECT 148.005 285.505 149.755 297.480 ;
        RECT 151.845 285.505 153.595 300.125 ;
        RECT 155.685 285.505 157.435 301.965 ;
        RECT 159.870 300.305 160.250 300.685 ;
        RECT 162.315 298.995 162.695 299.375 ;
        RECT 164.355 298.995 164.735 299.375 ;
        RECT 166.140 298.995 166.520 299.375 ;
        RECT 159.870 297.660 160.250 298.040 ;
        RECT 159.870 295.820 160.250 296.200 ;
        RECT 162.315 295.995 162.695 296.375 ;
        RECT 164.355 295.995 164.735 296.375 ;
        RECT 166.140 295.995 166.520 296.375 ;
        RECT 159.870 293.980 160.250 294.360 ;
        RECT 162.315 292.995 162.695 293.375 ;
        RECT 164.355 292.995 164.735 293.375 ;
        RECT 166.140 292.995 166.520 293.375 ;
        RECT 159.870 291.335 160.250 291.715 ;
        RECT 162.315 289.995 162.695 290.375 ;
        RECT 164.355 289.995 164.735 290.375 ;
        RECT 166.140 289.995 166.520 290.375 ;
        RECT 159.870 289.495 160.250 289.875 ;
        RECT 159.870 287.655 160.250 288.035 ;
        RECT 162.315 286.995 162.695 287.375 ;
        RECT 164.355 286.995 164.735 287.375 ;
        RECT 166.140 286.995 166.520 287.375 ;
        RECT 34.060 285.120 34.440 285.310 ;
        RECT 37.900 285.120 38.280 285.310 ;
        RECT 41.740 285.120 42.120 285.310 ;
        RECT 45.580 285.120 45.960 285.310 ;
        RECT 49.420 285.120 49.800 285.310 ;
        RECT 53.260 285.120 53.640 285.310 ;
        RECT 57.100 285.120 57.480 285.310 ;
        RECT 60.940 285.120 61.320 285.310 ;
        RECT 66.510 285.120 66.890 285.310 ;
        RECT 70.350 285.120 70.730 285.310 ;
        RECT 74.190 285.120 74.570 285.310 ;
        RECT 78.030 285.120 78.410 285.310 ;
        RECT 81.870 285.120 82.250 285.310 ;
        RECT 85.710 285.120 86.090 285.310 ;
        RECT 89.550 285.120 89.930 285.310 ;
        RECT 93.390 285.120 93.770 285.310 ;
        RECT 98.960 285.120 99.340 285.310 ;
        RECT 102.800 285.120 103.180 285.310 ;
        RECT 106.640 285.120 107.020 285.310 ;
        RECT 110.480 285.120 110.860 285.310 ;
        RECT 114.320 285.120 114.700 285.310 ;
        RECT 118.160 285.120 118.540 285.310 ;
        RECT 122.000 285.120 122.380 285.310 ;
        RECT 125.840 285.120 126.220 285.310 ;
        RECT 131.410 285.120 131.790 285.310 ;
        RECT 135.250 285.120 135.630 285.310 ;
        RECT 139.090 285.120 139.470 285.310 ;
        RECT 142.930 285.120 143.310 285.310 ;
        RECT 146.770 285.120 147.150 285.310 ;
        RECT 150.610 285.120 150.990 285.310 ;
        RECT 154.450 285.120 154.830 285.310 ;
        RECT 158.290 285.120 158.670 285.310 ;
        RECT 28.390 284.310 166.790 285.120 ;
        RECT 25.200 282.495 25.580 282.875 ;
        RECT 28.390 282.860 29.200 284.310 ;
        RECT 161.300 284.120 161.680 284.310 ;
        RECT 163.340 284.120 163.720 284.310 ;
        RECT 165.380 284.120 165.760 284.310 ;
        RECT 161.300 282.860 161.680 283.050 ;
        RECT 163.340 282.860 163.720 283.050 ;
        RECT 165.380 282.860 165.760 283.050 ;
        RECT 28.390 282.050 166.790 282.860 ;
        RECT 32.140 281.860 32.520 282.050 ;
        RECT 35.980 281.860 36.360 282.050 ;
        RECT 39.820 281.860 40.200 282.050 ;
        RECT 43.660 281.860 44.040 282.050 ;
        RECT 47.500 281.860 47.880 282.050 ;
        RECT 51.340 281.860 51.720 282.050 ;
        RECT 55.180 281.860 55.560 282.050 ;
        RECT 59.020 281.860 59.400 282.050 ;
        RECT 64.590 281.860 64.970 282.050 ;
        RECT 68.430 281.860 68.810 282.050 ;
        RECT 72.270 281.860 72.650 282.050 ;
        RECT 76.110 281.860 76.490 282.050 ;
        RECT 79.950 281.860 80.330 282.050 ;
        RECT 83.790 281.860 84.170 282.050 ;
        RECT 87.630 281.860 88.010 282.050 ;
        RECT 91.470 281.860 91.850 282.050 ;
        RECT 97.040 281.860 97.420 282.050 ;
        RECT 100.880 281.860 101.260 282.050 ;
        RECT 104.720 281.860 105.100 282.050 ;
        RECT 108.560 281.860 108.940 282.050 ;
        RECT 112.400 281.860 112.780 282.050 ;
        RECT 116.240 281.860 116.620 282.050 ;
        RECT 120.080 281.860 120.460 282.050 ;
        RECT 123.920 281.860 124.300 282.050 ;
        RECT 129.490 281.860 129.870 282.050 ;
        RECT 133.330 281.860 133.710 282.050 ;
        RECT 137.170 281.860 137.550 282.050 ;
        RECT 141.010 281.860 141.390 282.050 ;
        RECT 144.850 281.860 145.230 282.050 ;
        RECT 148.690 281.860 149.070 282.050 ;
        RECT 152.530 281.860 152.910 282.050 ;
        RECT 156.370 281.860 156.750 282.050 ;
        RECT 25.200 279.495 25.580 279.875 ;
        RECT 27.480 277.160 27.830 281.350 ;
        RECT 25.200 276.495 25.580 276.875 ;
        RECT 28.110 275.805 28.460 279.720 ;
        RECT 29.120 279.495 29.500 279.875 ;
        RECT 31.920 278.530 34.160 278.910 ;
        RECT 37.215 277.810 38.965 281.665 ;
        RECT 29.120 276.495 29.500 276.875 ;
        RECT 31.920 276.690 34.160 277.070 ;
        RECT 41.055 275.965 42.805 281.665 ;
        RECT 27.705 275.480 28.460 275.805 ;
        RECT 28.110 275.475 28.460 275.480 ;
        RECT 31.920 274.845 34.160 275.225 ;
        RECT 31.925 274.085 34.165 274.465 ;
        RECT 25.200 273.495 25.580 273.875 ;
        RECT 29.120 273.495 29.500 273.875 ;
        RECT 44.895 273.325 46.645 281.665 ;
        RECT 31.920 272.205 34.160 272.585 ;
        RECT 48.735 271.485 50.485 281.665 ;
        RECT 25.200 270.495 25.580 270.875 ;
        RECT 29.120 270.495 29.500 270.875 ;
        RECT 31.920 270.365 34.160 270.745 ;
        RECT 52.575 269.640 54.325 281.665 ;
        RECT 31.920 268.520 34.160 268.900 ;
        RECT 25.200 267.495 25.580 267.875 ;
        RECT 29.120 267.495 29.500 267.875 ;
        RECT 31.925 267.760 34.165 268.140 ;
        RECT 56.415 267.000 58.165 281.665 ;
        RECT 31.920 265.880 34.160 266.260 ;
        RECT 60.255 265.160 62.005 281.665 ;
        RECT 62.520 279.090 62.900 279.470 ;
        RECT 64.370 278.530 66.610 278.910 ;
        RECT 69.665 277.810 71.415 281.665 ;
        RECT 62.520 277.250 62.900 277.630 ;
        RECT 64.370 276.690 66.610 277.070 ;
        RECT 73.505 275.965 75.255 281.665 ;
        RECT 62.520 275.405 62.900 275.785 ;
        RECT 64.370 274.845 66.610 275.225 ;
        RECT 64.375 274.085 66.615 274.465 ;
        RECT 77.345 273.325 79.095 281.665 ;
        RECT 62.520 272.765 62.900 273.145 ;
        RECT 64.370 272.205 66.610 272.585 ;
        RECT 81.185 271.485 82.935 281.665 ;
        RECT 62.520 270.925 62.900 271.305 ;
        RECT 64.370 270.365 66.610 270.745 ;
        RECT 85.025 269.640 86.775 281.665 ;
        RECT 62.520 269.080 62.900 269.460 ;
        RECT 64.370 268.520 66.610 268.900 ;
        RECT 64.375 267.760 66.615 268.140 ;
        RECT 88.865 267.000 90.615 281.665 ;
        RECT 62.520 266.440 62.900 266.820 ;
        RECT 64.370 265.880 66.610 266.260 ;
        RECT 92.705 265.160 94.455 281.665 ;
        RECT 94.970 279.090 95.350 279.470 ;
        RECT 96.820 278.530 99.060 278.910 ;
        RECT 102.115 277.810 103.865 281.665 ;
        RECT 94.970 277.250 95.350 277.630 ;
        RECT 96.820 276.690 99.060 277.070 ;
        RECT 105.955 275.965 107.705 281.665 ;
        RECT 94.970 275.405 95.350 275.785 ;
        RECT 96.820 274.845 99.060 275.225 ;
        RECT 96.825 274.085 99.065 274.465 ;
        RECT 109.795 273.325 111.545 281.665 ;
        RECT 94.970 272.765 95.350 273.145 ;
        RECT 96.820 272.205 99.060 272.585 ;
        RECT 113.635 271.485 115.385 281.665 ;
        RECT 94.970 270.925 95.350 271.305 ;
        RECT 96.820 270.365 99.060 270.745 ;
        RECT 117.475 269.640 119.225 281.665 ;
        RECT 94.970 269.080 95.350 269.460 ;
        RECT 96.820 268.520 99.060 268.900 ;
        RECT 96.825 267.760 99.065 268.140 ;
        RECT 121.315 267.000 123.065 281.665 ;
        RECT 94.970 266.440 95.350 266.820 ;
        RECT 96.820 265.880 99.060 266.260 ;
        RECT 125.155 265.160 126.905 281.665 ;
        RECT 127.420 279.090 127.800 279.470 ;
        RECT 129.270 278.530 131.510 278.910 ;
        RECT 134.565 277.810 136.315 281.665 ;
        RECT 127.420 277.250 127.800 277.630 ;
        RECT 129.270 276.690 131.510 277.070 ;
        RECT 138.405 275.965 140.155 281.665 ;
        RECT 127.420 275.405 127.800 275.785 ;
        RECT 129.270 274.845 131.510 275.225 ;
        RECT 129.275 274.085 131.515 274.465 ;
        RECT 142.245 273.325 143.995 281.665 ;
        RECT 127.420 272.765 127.800 273.145 ;
        RECT 129.270 272.205 131.510 272.585 ;
        RECT 146.085 271.485 147.835 281.665 ;
        RECT 127.420 270.925 127.800 271.305 ;
        RECT 129.270 270.365 131.510 270.745 ;
        RECT 149.925 269.640 151.675 281.665 ;
        RECT 127.420 269.080 127.800 269.460 ;
        RECT 129.270 268.520 131.510 268.900 ;
        RECT 129.275 267.760 131.515 268.140 ;
        RECT 153.765 267.000 155.515 281.665 ;
        RECT 127.420 266.440 127.800 266.820 ;
        RECT 129.270 265.880 131.510 266.260 ;
        RECT 157.605 265.160 159.355 281.665 ;
        RECT 162.315 280.995 162.695 281.375 ;
        RECT 164.355 280.995 164.735 281.375 ;
        RECT 166.140 280.995 166.520 281.375 ;
        RECT 159.870 279.090 160.250 279.470 ;
        RECT 162.315 277.995 162.695 278.375 ;
        RECT 164.355 277.995 164.735 278.375 ;
        RECT 166.140 277.995 166.520 278.375 ;
        RECT 159.870 277.250 160.250 277.630 ;
        RECT 159.870 275.405 160.250 275.785 ;
        RECT 162.315 274.995 162.695 275.375 ;
        RECT 164.355 274.995 164.735 275.375 ;
        RECT 166.140 274.995 166.520 275.375 ;
        RECT 159.870 272.765 160.250 273.145 ;
        RECT 162.315 271.995 162.695 272.375 ;
        RECT 164.355 271.995 164.735 272.375 ;
        RECT 166.140 271.995 166.520 272.375 ;
        RECT 159.870 270.925 160.250 271.305 ;
        RECT 159.870 269.080 160.250 269.460 ;
        RECT 162.315 268.995 162.695 269.375 ;
        RECT 164.355 268.995 164.735 269.375 ;
        RECT 166.140 268.995 166.520 269.375 ;
        RECT 159.870 266.440 160.250 266.820 ;
        RECT 162.315 265.995 162.695 266.375 ;
        RECT 164.355 265.995 164.735 266.375 ;
        RECT 166.140 265.995 166.520 266.375 ;
        RECT 25.200 264.495 25.580 264.875 ;
        RECT 29.120 264.495 29.500 264.875 ;
        RECT 62.520 264.600 62.900 264.980 ;
        RECT 94.970 264.600 95.350 264.980 ;
        RECT 127.420 264.600 127.800 264.980 ;
        RECT 159.870 264.600 160.250 264.980 ;
        RECT 31.920 264.040 34.160 264.420 ;
        RECT 64.370 264.040 66.610 264.420 ;
        RECT 96.820 264.040 99.060 264.420 ;
        RECT 129.270 264.040 131.510 264.420 ;
        RECT 31.920 263.320 34.160 263.700 ;
        RECT 64.370 263.320 66.610 263.700 ;
        RECT 96.820 263.320 99.060 263.700 ;
        RECT 129.270 263.320 131.510 263.700 ;
        RECT 62.520 262.760 62.900 263.140 ;
        RECT 94.970 262.760 95.350 263.140 ;
        RECT 127.420 262.760 127.800 263.140 ;
        RECT 159.870 262.760 160.250 263.140 ;
        RECT 25.200 261.110 25.580 261.490 ;
        RECT 29.120 261.110 29.500 261.490 ;
        RECT 31.920 261.480 34.160 261.860 ;
        RECT 31.925 259.595 34.165 259.975 ;
        RECT 31.920 258.835 34.160 259.215 ;
        RECT 25.200 258.110 25.580 258.490 ;
        RECT 29.120 258.110 29.500 258.490 ;
        RECT 31.920 256.995 34.160 257.375 ;
        RECT 25.200 255.110 25.580 255.490 ;
        RECT 29.120 255.110 29.500 255.490 ;
        RECT 31.920 255.155 34.160 255.535 ;
        RECT 31.925 253.270 34.165 253.650 ;
        RECT 31.920 252.510 34.160 252.890 ;
        RECT 25.200 252.110 25.580 252.490 ;
        RECT 29.120 252.110 29.500 252.490 ;
        RECT 31.920 250.670 34.160 251.050 ;
        RECT 25.200 249.110 25.580 249.490 ;
        RECT 29.120 249.110 29.500 249.490 ;
        RECT 31.920 248.830 34.160 249.210 ;
        RECT 25.200 246.110 25.580 246.490 ;
        RECT 29.120 246.110 29.500 246.490 ;
        RECT 35.295 246.120 37.045 249.930 ;
        RECT 39.135 246.120 40.885 251.770 ;
        RECT 42.975 246.120 44.725 254.415 ;
        RECT 46.815 246.120 48.565 256.255 ;
        RECT 50.655 246.120 52.405 258.095 ;
        RECT 54.495 246.120 56.245 260.740 ;
        RECT 58.335 246.120 60.085 262.580 ;
        RECT 64.370 261.480 66.610 261.860 ;
        RECT 62.520 260.920 62.900 261.300 ;
        RECT 64.375 259.595 66.615 259.975 ;
        RECT 64.370 258.835 66.610 259.215 ;
        RECT 62.520 258.275 62.900 258.655 ;
        RECT 64.370 256.995 66.610 257.375 ;
        RECT 62.520 256.435 62.900 256.815 ;
        RECT 64.370 255.155 66.610 255.535 ;
        RECT 62.520 254.595 62.900 254.975 ;
        RECT 64.375 253.270 66.615 253.650 ;
        RECT 64.370 252.510 66.610 252.890 ;
        RECT 62.520 251.950 62.900 252.330 ;
        RECT 64.370 250.670 66.610 251.050 ;
        RECT 62.520 250.110 62.900 250.490 ;
        RECT 64.370 248.830 66.610 249.210 ;
        RECT 62.520 248.270 62.900 248.650 ;
        RECT 67.745 246.120 69.495 249.930 ;
        RECT 71.585 246.120 73.335 251.770 ;
        RECT 75.425 246.120 77.175 254.415 ;
        RECT 79.265 246.120 81.015 256.255 ;
        RECT 83.105 246.120 84.855 258.095 ;
        RECT 86.945 246.120 88.695 260.740 ;
        RECT 90.785 246.120 92.535 262.580 ;
        RECT 96.820 261.480 99.060 261.860 ;
        RECT 94.970 260.920 95.350 261.300 ;
        RECT 96.825 259.595 99.065 259.975 ;
        RECT 96.820 258.835 99.060 259.215 ;
        RECT 94.970 258.275 95.350 258.655 ;
        RECT 96.820 256.995 99.060 257.375 ;
        RECT 94.970 256.435 95.350 256.815 ;
        RECT 96.820 255.155 99.060 255.535 ;
        RECT 94.970 254.595 95.350 254.975 ;
        RECT 96.825 253.270 99.065 253.650 ;
        RECT 96.820 252.510 99.060 252.890 ;
        RECT 94.970 251.950 95.350 252.330 ;
        RECT 96.820 250.670 99.060 251.050 ;
        RECT 94.970 250.110 95.350 250.490 ;
        RECT 96.820 248.830 99.060 249.210 ;
        RECT 94.970 248.270 95.350 248.650 ;
        RECT 100.195 246.120 101.945 249.930 ;
        RECT 104.035 246.120 105.785 251.770 ;
        RECT 107.875 246.120 109.625 254.415 ;
        RECT 111.715 246.120 113.465 256.255 ;
        RECT 115.555 246.120 117.305 258.095 ;
        RECT 119.395 246.120 121.145 260.740 ;
        RECT 123.235 246.120 124.985 262.580 ;
        RECT 129.270 261.480 131.510 261.860 ;
        RECT 127.420 260.920 127.800 261.300 ;
        RECT 129.275 259.595 131.515 259.975 ;
        RECT 129.270 258.835 131.510 259.215 ;
        RECT 127.420 258.275 127.800 258.655 ;
        RECT 129.270 256.995 131.510 257.375 ;
        RECT 127.420 256.435 127.800 256.815 ;
        RECT 129.270 255.155 131.510 255.535 ;
        RECT 127.420 254.595 127.800 254.975 ;
        RECT 129.275 253.270 131.515 253.650 ;
        RECT 129.270 252.510 131.510 252.890 ;
        RECT 127.420 251.950 127.800 252.330 ;
        RECT 129.270 250.670 131.510 251.050 ;
        RECT 127.420 250.110 127.800 250.490 ;
        RECT 129.270 248.830 131.510 249.210 ;
        RECT 127.420 248.270 127.800 248.650 ;
        RECT 132.645 246.120 134.395 249.930 ;
        RECT 136.485 246.120 138.235 251.770 ;
        RECT 140.325 246.120 142.075 254.415 ;
        RECT 144.165 246.120 145.915 256.255 ;
        RECT 148.005 246.120 149.755 258.095 ;
        RECT 151.845 246.120 153.595 260.740 ;
        RECT 155.685 246.120 157.435 262.580 ;
        RECT 159.870 260.920 160.250 261.300 ;
        RECT 162.315 259.610 162.695 259.990 ;
        RECT 164.355 259.610 164.735 259.990 ;
        RECT 166.140 259.610 166.520 259.990 ;
        RECT 159.870 258.275 160.250 258.655 ;
        RECT 159.870 256.435 160.250 256.815 ;
        RECT 162.315 256.610 162.695 256.990 ;
        RECT 164.355 256.610 164.735 256.990 ;
        RECT 166.140 256.610 166.520 256.990 ;
        RECT 159.870 254.595 160.250 254.975 ;
        RECT 162.315 253.610 162.695 253.990 ;
        RECT 164.355 253.610 164.735 253.990 ;
        RECT 166.140 253.610 166.520 253.990 ;
        RECT 159.870 251.950 160.250 252.330 ;
        RECT 162.315 250.610 162.695 250.990 ;
        RECT 164.355 250.610 164.735 250.990 ;
        RECT 166.140 250.610 166.520 250.990 ;
        RECT 159.870 250.110 160.250 250.490 ;
        RECT 159.870 248.270 160.250 248.650 ;
        RECT 162.315 247.610 162.695 247.990 ;
        RECT 164.355 247.610 164.735 247.990 ;
        RECT 166.140 247.610 166.520 247.990 ;
        RECT 34.060 245.735 34.440 245.925 ;
        RECT 37.900 245.735 38.280 245.925 ;
        RECT 41.740 245.735 42.120 245.925 ;
        RECT 45.580 245.735 45.960 245.925 ;
        RECT 49.420 245.735 49.800 245.925 ;
        RECT 53.260 245.735 53.640 245.925 ;
        RECT 57.100 245.735 57.480 245.925 ;
        RECT 60.940 245.735 61.320 245.925 ;
        RECT 66.510 245.735 66.890 245.925 ;
        RECT 70.350 245.735 70.730 245.925 ;
        RECT 74.190 245.735 74.570 245.925 ;
        RECT 78.030 245.735 78.410 245.925 ;
        RECT 81.870 245.735 82.250 245.925 ;
        RECT 85.710 245.735 86.090 245.925 ;
        RECT 89.550 245.735 89.930 245.925 ;
        RECT 93.390 245.735 93.770 245.925 ;
        RECT 98.960 245.735 99.340 245.925 ;
        RECT 102.800 245.735 103.180 245.925 ;
        RECT 106.640 245.735 107.020 245.925 ;
        RECT 110.480 245.735 110.860 245.925 ;
        RECT 114.320 245.735 114.700 245.925 ;
        RECT 118.160 245.735 118.540 245.925 ;
        RECT 122.000 245.735 122.380 245.925 ;
        RECT 125.840 245.735 126.220 245.925 ;
        RECT 131.410 245.735 131.790 245.925 ;
        RECT 135.250 245.735 135.630 245.925 ;
        RECT 139.090 245.735 139.470 245.925 ;
        RECT 142.930 245.735 143.310 245.925 ;
        RECT 146.770 245.735 147.150 245.925 ;
        RECT 150.610 245.735 150.990 245.925 ;
        RECT 154.450 245.735 154.830 245.925 ;
        RECT 158.290 245.735 158.670 245.925 ;
        RECT 28.390 244.925 166.790 245.735 ;
        RECT 25.200 243.110 25.580 243.490 ;
        RECT 28.390 243.475 29.200 244.925 ;
        RECT 161.300 244.735 161.680 244.925 ;
        RECT 163.340 244.735 163.720 244.925 ;
        RECT 165.380 244.735 165.760 244.925 ;
        RECT 161.300 243.475 161.680 243.665 ;
        RECT 163.340 243.475 163.720 243.665 ;
        RECT 165.380 243.475 165.760 243.665 ;
        RECT 28.390 242.665 166.790 243.475 ;
        RECT 32.140 242.475 32.520 242.665 ;
        RECT 35.980 242.475 36.360 242.665 ;
        RECT 39.820 242.475 40.200 242.665 ;
        RECT 43.660 242.475 44.040 242.665 ;
        RECT 47.500 242.475 47.880 242.665 ;
        RECT 51.340 242.475 51.720 242.665 ;
        RECT 55.180 242.475 55.560 242.665 ;
        RECT 59.020 242.475 59.400 242.665 ;
        RECT 64.590 242.475 64.970 242.665 ;
        RECT 68.430 242.475 68.810 242.665 ;
        RECT 72.270 242.475 72.650 242.665 ;
        RECT 76.110 242.475 76.490 242.665 ;
        RECT 79.950 242.475 80.330 242.665 ;
        RECT 83.790 242.475 84.170 242.665 ;
        RECT 87.630 242.475 88.010 242.665 ;
        RECT 91.470 242.475 91.850 242.665 ;
        RECT 97.040 242.475 97.420 242.665 ;
        RECT 100.880 242.475 101.260 242.665 ;
        RECT 104.720 242.475 105.100 242.665 ;
        RECT 108.560 242.475 108.940 242.665 ;
        RECT 112.400 242.475 112.780 242.665 ;
        RECT 116.240 242.475 116.620 242.665 ;
        RECT 120.080 242.475 120.460 242.665 ;
        RECT 123.920 242.475 124.300 242.665 ;
        RECT 129.490 242.475 129.870 242.665 ;
        RECT 133.330 242.475 133.710 242.665 ;
        RECT 137.170 242.475 137.550 242.665 ;
        RECT 141.010 242.475 141.390 242.665 ;
        RECT 144.850 242.475 145.230 242.665 ;
        RECT 148.690 242.475 149.070 242.665 ;
        RECT 152.530 242.475 152.910 242.665 ;
        RECT 156.370 242.475 156.750 242.665 ;
        RECT 25.200 240.110 25.580 240.490 ;
        RECT 27.480 237.775 27.830 241.965 ;
        RECT 25.200 237.110 25.580 237.490 ;
        RECT 28.110 236.420 28.460 240.335 ;
        RECT 29.120 240.110 29.500 240.490 ;
        RECT 31.920 239.145 34.160 239.525 ;
        RECT 37.215 238.425 38.965 242.280 ;
        RECT 29.120 237.110 29.500 237.490 ;
        RECT 31.920 237.305 34.160 237.685 ;
        RECT 41.055 236.580 42.805 242.280 ;
        RECT 27.705 236.095 28.460 236.420 ;
        RECT 28.110 236.090 28.460 236.095 ;
        RECT 31.920 235.460 34.160 235.840 ;
        RECT 31.925 234.700 34.165 235.080 ;
        RECT 25.200 234.110 25.580 234.490 ;
        RECT 29.120 234.110 29.500 234.490 ;
        RECT 44.895 233.940 46.645 242.280 ;
        RECT 31.920 232.820 34.160 233.200 ;
        RECT 48.735 232.100 50.485 242.280 ;
        RECT 25.200 231.110 25.580 231.490 ;
        RECT 29.120 231.110 29.500 231.490 ;
        RECT 31.920 230.980 34.160 231.360 ;
        RECT 52.575 230.255 54.325 242.280 ;
        RECT 31.920 229.135 34.160 229.515 ;
        RECT 25.200 228.110 25.580 228.490 ;
        RECT 29.120 228.110 29.500 228.490 ;
        RECT 31.925 228.375 34.165 228.755 ;
        RECT 56.415 227.615 58.165 242.280 ;
        RECT 31.920 226.495 34.160 226.875 ;
        RECT 60.255 225.775 62.005 242.280 ;
        RECT 62.520 239.705 62.900 240.085 ;
        RECT 64.370 239.145 66.610 239.525 ;
        RECT 69.665 238.425 71.415 242.280 ;
        RECT 62.520 237.865 62.900 238.245 ;
        RECT 64.370 237.305 66.610 237.685 ;
        RECT 73.505 236.580 75.255 242.280 ;
        RECT 62.520 236.020 62.900 236.400 ;
        RECT 64.370 235.460 66.610 235.840 ;
        RECT 64.375 234.700 66.615 235.080 ;
        RECT 77.345 233.940 79.095 242.280 ;
        RECT 62.520 233.380 62.900 233.760 ;
        RECT 64.370 232.820 66.610 233.200 ;
        RECT 81.185 232.100 82.935 242.280 ;
        RECT 62.520 231.540 62.900 231.920 ;
        RECT 64.370 230.980 66.610 231.360 ;
        RECT 85.025 230.255 86.775 242.280 ;
        RECT 62.520 229.695 62.900 230.075 ;
        RECT 64.370 229.135 66.610 229.515 ;
        RECT 64.375 228.375 66.615 228.755 ;
        RECT 88.865 227.615 90.615 242.280 ;
        RECT 62.520 227.055 62.900 227.435 ;
        RECT 64.370 226.495 66.610 226.875 ;
        RECT 92.705 225.775 94.455 242.280 ;
        RECT 94.970 239.705 95.350 240.085 ;
        RECT 96.820 239.145 99.060 239.525 ;
        RECT 102.115 238.425 103.865 242.280 ;
        RECT 94.970 237.865 95.350 238.245 ;
        RECT 96.820 237.305 99.060 237.685 ;
        RECT 105.955 236.580 107.705 242.280 ;
        RECT 94.970 236.020 95.350 236.400 ;
        RECT 96.820 235.460 99.060 235.840 ;
        RECT 96.825 234.700 99.065 235.080 ;
        RECT 109.795 233.940 111.545 242.280 ;
        RECT 94.970 233.380 95.350 233.760 ;
        RECT 96.820 232.820 99.060 233.200 ;
        RECT 113.635 232.100 115.385 242.280 ;
        RECT 94.970 231.540 95.350 231.920 ;
        RECT 96.820 230.980 99.060 231.360 ;
        RECT 117.475 230.255 119.225 242.280 ;
        RECT 94.970 229.695 95.350 230.075 ;
        RECT 96.820 229.135 99.060 229.515 ;
        RECT 96.825 228.375 99.065 228.755 ;
        RECT 121.315 227.615 123.065 242.280 ;
        RECT 94.970 227.055 95.350 227.435 ;
        RECT 96.820 226.495 99.060 226.875 ;
        RECT 125.155 225.775 126.905 242.280 ;
        RECT 127.420 239.705 127.800 240.085 ;
        RECT 129.270 239.145 131.510 239.525 ;
        RECT 134.565 238.425 136.315 242.280 ;
        RECT 127.420 237.865 127.800 238.245 ;
        RECT 129.270 237.305 131.510 237.685 ;
        RECT 138.405 236.580 140.155 242.280 ;
        RECT 127.420 236.020 127.800 236.400 ;
        RECT 129.270 235.460 131.510 235.840 ;
        RECT 129.275 234.700 131.515 235.080 ;
        RECT 142.245 233.940 143.995 242.280 ;
        RECT 127.420 233.380 127.800 233.760 ;
        RECT 129.270 232.820 131.510 233.200 ;
        RECT 146.085 232.100 147.835 242.280 ;
        RECT 127.420 231.540 127.800 231.920 ;
        RECT 129.270 230.980 131.510 231.360 ;
        RECT 149.925 230.255 151.675 242.280 ;
        RECT 127.420 229.695 127.800 230.075 ;
        RECT 129.270 229.135 131.510 229.515 ;
        RECT 129.275 228.375 131.515 228.755 ;
        RECT 153.765 227.615 155.515 242.280 ;
        RECT 127.420 227.055 127.800 227.435 ;
        RECT 129.270 226.495 131.510 226.875 ;
        RECT 157.605 225.775 159.355 242.280 ;
        RECT 162.315 241.610 162.695 241.990 ;
        RECT 164.355 241.610 164.735 241.990 ;
        RECT 166.140 241.610 166.520 241.990 ;
        RECT 159.870 239.705 160.250 240.085 ;
        RECT 162.315 238.610 162.695 238.990 ;
        RECT 164.355 238.610 164.735 238.990 ;
        RECT 166.140 238.610 166.520 238.990 ;
        RECT 159.870 237.865 160.250 238.245 ;
        RECT 159.870 236.020 160.250 236.400 ;
        RECT 162.315 235.610 162.695 235.990 ;
        RECT 164.355 235.610 164.735 235.990 ;
        RECT 166.140 235.610 166.520 235.990 ;
        RECT 159.870 233.380 160.250 233.760 ;
        RECT 162.315 232.610 162.695 232.990 ;
        RECT 164.355 232.610 164.735 232.990 ;
        RECT 166.140 232.610 166.520 232.990 ;
        RECT 159.870 231.540 160.250 231.920 ;
        RECT 159.870 229.695 160.250 230.075 ;
        RECT 162.315 229.610 162.695 229.990 ;
        RECT 164.355 229.610 164.735 229.990 ;
        RECT 166.140 229.610 166.520 229.990 ;
        RECT 159.870 227.055 160.250 227.435 ;
        RECT 162.315 226.610 162.695 226.990 ;
        RECT 164.355 226.610 164.735 226.990 ;
        RECT 166.140 226.610 166.520 226.990 ;
        RECT 25.200 225.110 25.580 225.490 ;
        RECT 29.120 225.110 29.500 225.490 ;
        RECT 62.520 225.215 62.900 225.595 ;
        RECT 94.970 225.215 95.350 225.595 ;
        RECT 127.420 225.215 127.800 225.595 ;
        RECT 159.870 225.215 160.250 225.595 ;
        RECT 31.920 224.655 34.160 225.035 ;
        RECT 64.370 224.655 66.610 225.035 ;
        RECT 96.820 224.655 99.060 225.035 ;
        RECT 129.270 224.655 131.510 225.035 ;
        RECT 31.920 223.935 34.160 224.315 ;
        RECT 64.370 223.935 66.610 224.315 ;
        RECT 96.820 223.935 99.060 224.315 ;
        RECT 129.270 223.935 131.510 224.315 ;
        RECT 62.520 223.375 62.900 223.755 ;
        RECT 94.970 223.375 95.350 223.755 ;
        RECT 127.420 223.375 127.800 223.755 ;
        RECT 159.870 223.375 160.250 223.755 ;
        RECT 25.200 221.725 25.580 222.105 ;
        RECT 29.120 221.725 29.500 222.105 ;
        RECT 31.920 222.095 34.160 222.475 ;
        RECT 31.925 220.210 34.165 220.590 ;
        RECT 31.920 219.450 34.160 219.830 ;
        RECT 25.200 218.725 25.580 219.105 ;
        RECT 29.120 218.725 29.500 219.105 ;
        RECT 31.920 217.610 34.160 217.990 ;
        RECT 25.200 215.725 25.580 216.105 ;
        RECT 29.120 215.725 29.500 216.105 ;
        RECT 31.920 215.770 34.160 216.150 ;
        RECT 31.925 213.885 34.165 214.265 ;
        RECT 31.920 213.125 34.160 213.505 ;
        RECT 25.200 212.725 25.580 213.105 ;
        RECT 29.120 212.725 29.500 213.105 ;
        RECT 31.920 211.285 34.160 211.665 ;
        RECT 25.200 209.725 25.580 210.105 ;
        RECT 29.120 209.725 29.500 210.105 ;
        RECT 31.920 209.445 34.160 209.825 ;
        RECT 25.200 206.725 25.580 207.105 ;
        RECT 29.120 206.725 29.500 207.105 ;
        RECT 35.295 206.735 37.045 210.545 ;
        RECT 39.135 206.735 40.885 212.385 ;
        RECT 42.975 206.735 44.725 215.030 ;
        RECT 46.815 206.735 48.565 216.870 ;
        RECT 50.655 206.735 52.405 218.710 ;
        RECT 54.495 206.735 56.245 221.355 ;
        RECT 58.335 206.735 60.085 223.195 ;
        RECT 64.370 222.095 66.610 222.475 ;
        RECT 62.520 221.535 62.900 221.915 ;
        RECT 64.375 220.210 66.615 220.590 ;
        RECT 64.370 219.450 66.610 219.830 ;
        RECT 62.520 218.890 62.900 219.270 ;
        RECT 64.370 217.610 66.610 217.990 ;
        RECT 62.520 217.050 62.900 217.430 ;
        RECT 64.370 215.770 66.610 216.150 ;
        RECT 62.520 215.210 62.900 215.590 ;
        RECT 64.375 213.885 66.615 214.265 ;
        RECT 64.370 213.125 66.610 213.505 ;
        RECT 62.520 212.565 62.900 212.945 ;
        RECT 64.370 211.285 66.610 211.665 ;
        RECT 62.520 210.725 62.900 211.105 ;
        RECT 64.370 209.445 66.610 209.825 ;
        RECT 62.520 208.885 62.900 209.265 ;
        RECT 67.745 206.735 69.495 210.545 ;
        RECT 71.585 206.735 73.335 212.385 ;
        RECT 75.425 206.735 77.175 215.030 ;
        RECT 79.265 206.735 81.015 216.870 ;
        RECT 83.105 206.735 84.855 218.710 ;
        RECT 86.945 206.735 88.695 221.355 ;
        RECT 90.785 206.735 92.535 223.195 ;
        RECT 96.820 222.095 99.060 222.475 ;
        RECT 94.970 221.535 95.350 221.915 ;
        RECT 96.825 220.210 99.065 220.590 ;
        RECT 96.820 219.450 99.060 219.830 ;
        RECT 94.970 218.890 95.350 219.270 ;
        RECT 96.820 217.610 99.060 217.990 ;
        RECT 94.970 217.050 95.350 217.430 ;
        RECT 96.820 215.770 99.060 216.150 ;
        RECT 94.970 215.210 95.350 215.590 ;
        RECT 96.825 213.885 99.065 214.265 ;
        RECT 96.820 213.125 99.060 213.505 ;
        RECT 94.970 212.565 95.350 212.945 ;
        RECT 96.820 211.285 99.060 211.665 ;
        RECT 94.970 210.725 95.350 211.105 ;
        RECT 96.820 209.445 99.060 209.825 ;
        RECT 94.970 208.885 95.350 209.265 ;
        RECT 100.195 206.735 101.945 210.545 ;
        RECT 104.035 206.735 105.785 212.385 ;
        RECT 107.875 206.735 109.625 215.030 ;
        RECT 111.715 206.735 113.465 216.870 ;
        RECT 115.555 206.735 117.305 218.710 ;
        RECT 119.395 206.735 121.145 221.355 ;
        RECT 123.235 206.735 124.985 223.195 ;
        RECT 129.270 222.095 131.510 222.475 ;
        RECT 127.420 221.535 127.800 221.915 ;
        RECT 129.275 220.210 131.515 220.590 ;
        RECT 129.270 219.450 131.510 219.830 ;
        RECT 127.420 218.890 127.800 219.270 ;
        RECT 129.270 217.610 131.510 217.990 ;
        RECT 127.420 217.050 127.800 217.430 ;
        RECT 129.270 215.770 131.510 216.150 ;
        RECT 127.420 215.210 127.800 215.590 ;
        RECT 129.275 213.885 131.515 214.265 ;
        RECT 129.270 213.125 131.510 213.505 ;
        RECT 127.420 212.565 127.800 212.945 ;
        RECT 129.270 211.285 131.510 211.665 ;
        RECT 127.420 210.725 127.800 211.105 ;
        RECT 129.270 209.445 131.510 209.825 ;
        RECT 127.420 208.885 127.800 209.265 ;
        RECT 132.645 206.735 134.395 210.545 ;
        RECT 136.485 206.735 138.235 212.385 ;
        RECT 140.325 206.735 142.075 215.030 ;
        RECT 144.165 206.735 145.915 216.870 ;
        RECT 148.005 206.735 149.755 218.710 ;
        RECT 151.845 206.735 153.595 221.355 ;
        RECT 155.685 206.735 157.435 223.195 ;
        RECT 159.870 221.535 160.250 221.915 ;
        RECT 162.315 220.225 162.695 220.605 ;
        RECT 164.355 220.225 164.735 220.605 ;
        RECT 166.140 220.225 166.520 220.605 ;
        RECT 159.870 218.890 160.250 219.270 ;
        RECT 159.870 217.050 160.250 217.430 ;
        RECT 162.315 217.225 162.695 217.605 ;
        RECT 164.355 217.225 164.735 217.605 ;
        RECT 166.140 217.225 166.520 217.605 ;
        RECT 159.870 215.210 160.250 215.590 ;
        RECT 162.315 214.225 162.695 214.605 ;
        RECT 164.355 214.225 164.735 214.605 ;
        RECT 166.140 214.225 166.520 214.605 ;
        RECT 159.870 212.565 160.250 212.945 ;
        RECT 162.315 211.225 162.695 211.605 ;
        RECT 164.355 211.225 164.735 211.605 ;
        RECT 166.140 211.225 166.520 211.605 ;
        RECT 159.870 210.725 160.250 211.105 ;
        RECT 159.870 208.885 160.250 209.265 ;
        RECT 162.315 208.225 162.695 208.605 ;
        RECT 164.355 208.225 164.735 208.605 ;
        RECT 166.140 208.225 166.520 208.605 ;
        RECT 34.060 206.350 34.440 206.540 ;
        RECT 37.900 206.350 38.280 206.540 ;
        RECT 41.740 206.350 42.120 206.540 ;
        RECT 45.580 206.350 45.960 206.540 ;
        RECT 49.420 206.350 49.800 206.540 ;
        RECT 53.260 206.350 53.640 206.540 ;
        RECT 57.100 206.350 57.480 206.540 ;
        RECT 60.940 206.350 61.320 206.540 ;
        RECT 66.510 206.350 66.890 206.540 ;
        RECT 70.350 206.350 70.730 206.540 ;
        RECT 74.190 206.350 74.570 206.540 ;
        RECT 78.030 206.350 78.410 206.540 ;
        RECT 81.870 206.350 82.250 206.540 ;
        RECT 85.710 206.350 86.090 206.540 ;
        RECT 89.550 206.350 89.930 206.540 ;
        RECT 93.390 206.350 93.770 206.540 ;
        RECT 98.960 206.350 99.340 206.540 ;
        RECT 102.800 206.350 103.180 206.540 ;
        RECT 106.640 206.350 107.020 206.540 ;
        RECT 110.480 206.350 110.860 206.540 ;
        RECT 114.320 206.350 114.700 206.540 ;
        RECT 118.160 206.350 118.540 206.540 ;
        RECT 122.000 206.350 122.380 206.540 ;
        RECT 125.840 206.350 126.220 206.540 ;
        RECT 131.410 206.350 131.790 206.540 ;
        RECT 135.250 206.350 135.630 206.540 ;
        RECT 139.090 206.350 139.470 206.540 ;
        RECT 142.930 206.350 143.310 206.540 ;
        RECT 146.770 206.350 147.150 206.540 ;
        RECT 150.610 206.350 150.990 206.540 ;
        RECT 154.450 206.350 154.830 206.540 ;
        RECT 158.290 206.350 158.670 206.540 ;
        RECT 28.390 205.540 166.790 206.350 ;
        RECT 25.200 203.725 25.580 204.105 ;
        RECT 28.390 204.090 29.200 205.540 ;
        RECT 161.300 205.350 161.680 205.540 ;
        RECT 163.340 205.350 163.720 205.540 ;
        RECT 165.380 205.350 165.760 205.540 ;
        RECT 161.300 204.090 161.680 204.280 ;
        RECT 163.340 204.090 163.720 204.280 ;
        RECT 165.380 204.090 165.760 204.280 ;
        RECT 28.390 203.280 166.790 204.090 ;
        RECT 32.140 203.090 32.520 203.280 ;
        RECT 35.980 203.090 36.360 203.280 ;
        RECT 39.820 203.090 40.200 203.280 ;
        RECT 43.660 203.090 44.040 203.280 ;
        RECT 47.500 203.090 47.880 203.280 ;
        RECT 51.340 203.090 51.720 203.280 ;
        RECT 55.180 203.090 55.560 203.280 ;
        RECT 59.020 203.090 59.400 203.280 ;
        RECT 64.590 203.090 64.970 203.280 ;
        RECT 68.430 203.090 68.810 203.280 ;
        RECT 72.270 203.090 72.650 203.280 ;
        RECT 76.110 203.090 76.490 203.280 ;
        RECT 79.950 203.090 80.330 203.280 ;
        RECT 83.790 203.090 84.170 203.280 ;
        RECT 87.630 203.090 88.010 203.280 ;
        RECT 91.470 203.090 91.850 203.280 ;
        RECT 97.040 203.090 97.420 203.280 ;
        RECT 100.880 203.090 101.260 203.280 ;
        RECT 104.720 203.090 105.100 203.280 ;
        RECT 108.560 203.090 108.940 203.280 ;
        RECT 112.400 203.090 112.780 203.280 ;
        RECT 116.240 203.090 116.620 203.280 ;
        RECT 120.080 203.090 120.460 203.280 ;
        RECT 123.920 203.090 124.300 203.280 ;
        RECT 129.490 203.090 129.870 203.280 ;
        RECT 133.330 203.090 133.710 203.280 ;
        RECT 137.170 203.090 137.550 203.280 ;
        RECT 141.010 203.090 141.390 203.280 ;
        RECT 144.850 203.090 145.230 203.280 ;
        RECT 148.690 203.090 149.070 203.280 ;
        RECT 152.530 203.090 152.910 203.280 ;
        RECT 156.370 203.090 156.750 203.280 ;
        RECT 25.200 200.725 25.580 201.105 ;
        RECT 27.480 198.390 27.830 202.580 ;
        RECT 25.200 197.725 25.580 198.105 ;
        RECT 28.110 197.035 28.460 200.950 ;
        RECT 29.120 200.725 29.500 201.105 ;
        RECT 31.920 199.760 34.160 200.140 ;
        RECT 37.215 199.040 38.965 202.895 ;
        RECT 29.120 197.725 29.500 198.105 ;
        RECT 31.920 197.920 34.160 198.300 ;
        RECT 41.055 197.195 42.805 202.895 ;
        RECT 27.705 196.710 28.460 197.035 ;
        RECT 28.110 196.705 28.460 196.710 ;
        RECT 31.920 196.075 34.160 196.455 ;
        RECT 31.925 195.315 34.165 195.695 ;
        RECT 25.200 194.725 25.580 195.105 ;
        RECT 29.120 194.725 29.500 195.105 ;
        RECT 44.895 194.555 46.645 202.895 ;
        RECT 31.920 193.435 34.160 193.815 ;
        RECT 48.735 192.715 50.485 202.895 ;
        RECT 25.200 191.725 25.580 192.105 ;
        RECT 29.120 191.725 29.500 192.105 ;
        RECT 31.920 191.595 34.160 191.975 ;
        RECT 52.575 190.870 54.325 202.895 ;
        RECT 31.920 189.750 34.160 190.130 ;
        RECT 25.200 188.725 25.580 189.105 ;
        RECT 29.120 188.725 29.500 189.105 ;
        RECT 31.925 188.990 34.165 189.370 ;
        RECT 56.415 188.230 58.165 202.895 ;
        RECT 31.920 187.110 34.160 187.490 ;
        RECT 60.255 186.390 62.005 202.895 ;
        RECT 62.520 200.320 62.900 200.700 ;
        RECT 64.370 199.760 66.610 200.140 ;
        RECT 69.665 199.040 71.415 202.895 ;
        RECT 62.520 198.480 62.900 198.860 ;
        RECT 64.370 197.920 66.610 198.300 ;
        RECT 73.505 197.195 75.255 202.895 ;
        RECT 62.520 196.635 62.900 197.015 ;
        RECT 64.370 196.075 66.610 196.455 ;
        RECT 64.375 195.315 66.615 195.695 ;
        RECT 77.345 194.555 79.095 202.895 ;
        RECT 62.520 193.995 62.900 194.375 ;
        RECT 64.370 193.435 66.610 193.815 ;
        RECT 81.185 192.715 82.935 202.895 ;
        RECT 62.520 192.155 62.900 192.535 ;
        RECT 64.370 191.595 66.610 191.975 ;
        RECT 85.025 190.870 86.775 202.895 ;
        RECT 62.520 190.310 62.900 190.690 ;
        RECT 64.370 189.750 66.610 190.130 ;
        RECT 64.375 188.990 66.615 189.370 ;
        RECT 88.865 188.230 90.615 202.895 ;
        RECT 62.520 187.670 62.900 188.050 ;
        RECT 64.370 187.110 66.610 187.490 ;
        RECT 92.705 186.390 94.455 202.895 ;
        RECT 94.970 200.320 95.350 200.700 ;
        RECT 96.820 199.760 99.060 200.140 ;
        RECT 102.115 199.040 103.865 202.895 ;
        RECT 94.970 198.480 95.350 198.860 ;
        RECT 96.820 197.920 99.060 198.300 ;
        RECT 105.955 197.195 107.705 202.895 ;
        RECT 94.970 196.635 95.350 197.015 ;
        RECT 96.820 196.075 99.060 196.455 ;
        RECT 96.825 195.315 99.065 195.695 ;
        RECT 109.795 194.555 111.545 202.895 ;
        RECT 94.970 193.995 95.350 194.375 ;
        RECT 96.820 193.435 99.060 193.815 ;
        RECT 113.635 192.715 115.385 202.895 ;
        RECT 94.970 192.155 95.350 192.535 ;
        RECT 96.820 191.595 99.060 191.975 ;
        RECT 117.475 190.870 119.225 202.895 ;
        RECT 94.970 190.310 95.350 190.690 ;
        RECT 96.820 189.750 99.060 190.130 ;
        RECT 96.825 188.990 99.065 189.370 ;
        RECT 121.315 188.230 123.065 202.895 ;
        RECT 94.970 187.670 95.350 188.050 ;
        RECT 96.820 187.110 99.060 187.490 ;
        RECT 125.155 186.390 126.905 202.895 ;
        RECT 127.420 200.320 127.800 200.700 ;
        RECT 129.270 199.760 131.510 200.140 ;
        RECT 134.565 199.040 136.315 202.895 ;
        RECT 127.420 198.480 127.800 198.860 ;
        RECT 129.270 197.920 131.510 198.300 ;
        RECT 138.405 197.195 140.155 202.895 ;
        RECT 127.420 196.635 127.800 197.015 ;
        RECT 129.270 196.075 131.510 196.455 ;
        RECT 129.275 195.315 131.515 195.695 ;
        RECT 142.245 194.555 143.995 202.895 ;
        RECT 127.420 193.995 127.800 194.375 ;
        RECT 129.270 193.435 131.510 193.815 ;
        RECT 146.085 192.715 147.835 202.895 ;
        RECT 127.420 192.155 127.800 192.535 ;
        RECT 129.270 191.595 131.510 191.975 ;
        RECT 149.925 190.870 151.675 202.895 ;
        RECT 127.420 190.310 127.800 190.690 ;
        RECT 129.270 189.750 131.510 190.130 ;
        RECT 129.275 188.990 131.515 189.370 ;
        RECT 153.765 188.230 155.515 202.895 ;
        RECT 127.420 187.670 127.800 188.050 ;
        RECT 129.270 187.110 131.510 187.490 ;
        RECT 157.605 186.390 159.355 202.895 ;
        RECT 162.315 202.225 162.695 202.605 ;
        RECT 164.355 202.225 164.735 202.605 ;
        RECT 166.140 202.225 166.520 202.605 ;
        RECT 159.870 200.320 160.250 200.700 ;
        RECT 162.315 199.225 162.695 199.605 ;
        RECT 164.355 199.225 164.735 199.605 ;
        RECT 166.140 199.225 166.520 199.605 ;
        RECT 159.870 198.480 160.250 198.860 ;
        RECT 159.870 196.635 160.250 197.015 ;
        RECT 162.315 196.225 162.695 196.605 ;
        RECT 164.355 196.225 164.735 196.605 ;
        RECT 166.140 196.225 166.520 196.605 ;
        RECT 159.870 193.995 160.250 194.375 ;
        RECT 162.315 193.225 162.695 193.605 ;
        RECT 164.355 193.225 164.735 193.605 ;
        RECT 166.140 193.225 166.520 193.605 ;
        RECT 159.870 192.155 160.250 192.535 ;
        RECT 159.870 190.310 160.250 190.690 ;
        RECT 162.315 190.225 162.695 190.605 ;
        RECT 164.355 190.225 164.735 190.605 ;
        RECT 166.140 190.225 166.520 190.605 ;
        RECT 159.870 187.670 160.250 188.050 ;
        RECT 162.315 187.225 162.695 187.605 ;
        RECT 164.355 187.225 164.735 187.605 ;
        RECT 166.140 187.225 166.520 187.605 ;
        RECT 25.200 185.725 25.580 186.105 ;
        RECT 29.120 185.725 29.500 186.105 ;
        RECT 62.520 185.830 62.900 186.210 ;
        RECT 94.970 185.830 95.350 186.210 ;
        RECT 127.420 185.830 127.800 186.210 ;
        RECT 159.870 185.830 160.250 186.210 ;
        RECT 31.920 185.270 34.160 185.650 ;
        RECT 64.370 185.270 66.610 185.650 ;
        RECT 96.820 185.270 99.060 185.650 ;
        RECT 129.270 185.270 131.510 185.650 ;
        RECT 31.920 184.550 34.160 184.930 ;
        RECT 64.370 184.550 66.610 184.930 ;
        RECT 96.820 184.550 99.060 184.930 ;
        RECT 129.270 184.550 131.510 184.930 ;
        RECT 62.520 183.990 62.900 184.370 ;
        RECT 94.970 183.990 95.350 184.370 ;
        RECT 127.420 183.990 127.800 184.370 ;
        RECT 159.870 183.990 160.250 184.370 ;
        RECT 25.200 182.340 25.580 182.720 ;
        RECT 29.120 182.340 29.500 182.720 ;
        RECT 31.920 182.710 34.160 183.090 ;
        RECT 31.925 180.825 34.165 181.205 ;
        RECT 31.920 180.065 34.160 180.445 ;
        RECT 25.200 179.340 25.580 179.720 ;
        RECT 29.120 179.340 29.500 179.720 ;
        RECT 31.920 178.225 34.160 178.605 ;
        RECT 25.200 176.340 25.580 176.720 ;
        RECT 29.120 176.340 29.500 176.720 ;
        RECT 31.920 176.385 34.160 176.765 ;
        RECT 31.925 174.500 34.165 174.880 ;
        RECT 31.920 173.740 34.160 174.120 ;
        RECT 25.200 173.340 25.580 173.720 ;
        RECT 29.120 173.340 29.500 173.720 ;
        RECT 31.920 171.900 34.160 172.280 ;
        RECT 25.200 170.340 25.580 170.720 ;
        RECT 29.120 170.340 29.500 170.720 ;
        RECT 31.920 170.060 34.160 170.440 ;
        RECT 25.200 167.340 25.580 167.720 ;
        RECT 29.120 167.340 29.500 167.720 ;
        RECT 35.295 167.350 37.045 171.160 ;
        RECT 39.135 167.350 40.885 173.000 ;
        RECT 42.975 167.350 44.725 175.645 ;
        RECT 46.815 167.350 48.565 177.485 ;
        RECT 50.655 167.350 52.405 179.325 ;
        RECT 54.495 167.350 56.245 181.970 ;
        RECT 58.335 167.350 60.085 183.810 ;
        RECT 64.370 182.710 66.610 183.090 ;
        RECT 62.520 182.150 62.900 182.530 ;
        RECT 64.375 180.825 66.615 181.205 ;
        RECT 64.370 180.065 66.610 180.445 ;
        RECT 62.520 179.505 62.900 179.885 ;
        RECT 64.370 178.225 66.610 178.605 ;
        RECT 62.520 177.665 62.900 178.045 ;
        RECT 64.370 176.385 66.610 176.765 ;
        RECT 62.520 175.825 62.900 176.205 ;
        RECT 64.375 174.500 66.615 174.880 ;
        RECT 64.370 173.740 66.610 174.120 ;
        RECT 62.520 173.180 62.900 173.560 ;
        RECT 64.370 171.900 66.610 172.280 ;
        RECT 62.520 171.340 62.900 171.720 ;
        RECT 64.370 170.060 66.610 170.440 ;
        RECT 62.520 169.500 62.900 169.880 ;
        RECT 67.745 167.350 69.495 171.160 ;
        RECT 71.585 167.350 73.335 173.000 ;
        RECT 75.425 167.350 77.175 175.645 ;
        RECT 79.265 167.350 81.015 177.485 ;
        RECT 83.105 167.350 84.855 179.325 ;
        RECT 86.945 167.350 88.695 181.970 ;
        RECT 90.785 167.350 92.535 183.810 ;
        RECT 96.820 182.710 99.060 183.090 ;
        RECT 94.970 182.150 95.350 182.530 ;
        RECT 96.825 180.825 99.065 181.205 ;
        RECT 96.820 180.065 99.060 180.445 ;
        RECT 94.970 179.505 95.350 179.885 ;
        RECT 96.820 178.225 99.060 178.605 ;
        RECT 94.970 177.665 95.350 178.045 ;
        RECT 96.820 176.385 99.060 176.765 ;
        RECT 94.970 175.825 95.350 176.205 ;
        RECT 96.825 174.500 99.065 174.880 ;
        RECT 96.820 173.740 99.060 174.120 ;
        RECT 94.970 173.180 95.350 173.560 ;
        RECT 96.820 171.900 99.060 172.280 ;
        RECT 94.970 171.340 95.350 171.720 ;
        RECT 96.820 170.060 99.060 170.440 ;
        RECT 94.970 169.500 95.350 169.880 ;
        RECT 100.195 167.350 101.945 171.160 ;
        RECT 104.035 167.350 105.785 173.000 ;
        RECT 107.875 167.350 109.625 175.645 ;
        RECT 111.715 167.350 113.465 177.485 ;
        RECT 115.555 167.350 117.305 179.325 ;
        RECT 119.395 167.350 121.145 181.970 ;
        RECT 123.235 167.350 124.985 183.810 ;
        RECT 129.270 182.710 131.510 183.090 ;
        RECT 127.420 182.150 127.800 182.530 ;
        RECT 129.275 180.825 131.515 181.205 ;
        RECT 129.270 180.065 131.510 180.445 ;
        RECT 127.420 179.505 127.800 179.885 ;
        RECT 129.270 178.225 131.510 178.605 ;
        RECT 127.420 177.665 127.800 178.045 ;
        RECT 129.270 176.385 131.510 176.765 ;
        RECT 127.420 175.825 127.800 176.205 ;
        RECT 129.275 174.500 131.515 174.880 ;
        RECT 129.270 173.740 131.510 174.120 ;
        RECT 127.420 173.180 127.800 173.560 ;
        RECT 129.270 171.900 131.510 172.280 ;
        RECT 127.420 171.340 127.800 171.720 ;
        RECT 129.270 170.060 131.510 170.440 ;
        RECT 127.420 169.500 127.800 169.880 ;
        RECT 132.645 167.350 134.395 171.160 ;
        RECT 136.485 167.350 138.235 173.000 ;
        RECT 140.325 167.350 142.075 175.645 ;
        RECT 144.165 167.350 145.915 177.485 ;
        RECT 148.005 167.350 149.755 179.325 ;
        RECT 151.845 167.350 153.595 181.970 ;
        RECT 155.685 167.350 157.435 183.810 ;
        RECT 159.870 182.150 160.250 182.530 ;
        RECT 162.315 180.840 162.695 181.220 ;
        RECT 164.355 180.840 164.735 181.220 ;
        RECT 166.140 180.840 166.520 181.220 ;
        RECT 159.870 179.505 160.250 179.885 ;
        RECT 159.870 177.665 160.250 178.045 ;
        RECT 162.315 177.840 162.695 178.220 ;
        RECT 164.355 177.840 164.735 178.220 ;
        RECT 166.140 177.840 166.520 178.220 ;
        RECT 159.870 175.825 160.250 176.205 ;
        RECT 162.315 174.840 162.695 175.220 ;
        RECT 164.355 174.840 164.735 175.220 ;
        RECT 166.140 174.840 166.520 175.220 ;
        RECT 159.870 173.180 160.250 173.560 ;
        RECT 162.315 171.840 162.695 172.220 ;
        RECT 164.355 171.840 164.735 172.220 ;
        RECT 166.140 171.840 166.520 172.220 ;
        RECT 159.870 171.340 160.250 171.720 ;
        RECT 159.870 169.500 160.250 169.880 ;
        RECT 162.315 168.840 162.695 169.220 ;
        RECT 164.355 168.840 164.735 169.220 ;
        RECT 166.140 168.840 166.520 169.220 ;
        RECT 34.060 166.965 34.440 167.155 ;
        RECT 37.900 166.965 38.280 167.155 ;
        RECT 41.740 166.965 42.120 167.155 ;
        RECT 45.580 166.965 45.960 167.155 ;
        RECT 49.420 166.965 49.800 167.155 ;
        RECT 53.260 166.965 53.640 167.155 ;
        RECT 57.100 166.965 57.480 167.155 ;
        RECT 60.940 166.965 61.320 167.155 ;
        RECT 66.510 166.965 66.890 167.155 ;
        RECT 70.350 166.965 70.730 167.155 ;
        RECT 74.190 166.965 74.570 167.155 ;
        RECT 78.030 166.965 78.410 167.155 ;
        RECT 81.870 166.965 82.250 167.155 ;
        RECT 85.710 166.965 86.090 167.155 ;
        RECT 89.550 166.965 89.930 167.155 ;
        RECT 93.390 166.965 93.770 167.155 ;
        RECT 98.960 166.965 99.340 167.155 ;
        RECT 102.800 166.965 103.180 167.155 ;
        RECT 106.640 166.965 107.020 167.155 ;
        RECT 110.480 166.965 110.860 167.155 ;
        RECT 114.320 166.965 114.700 167.155 ;
        RECT 118.160 166.965 118.540 167.155 ;
        RECT 122.000 166.965 122.380 167.155 ;
        RECT 125.840 166.965 126.220 167.155 ;
        RECT 131.410 166.965 131.790 167.155 ;
        RECT 135.250 166.965 135.630 167.155 ;
        RECT 139.090 166.965 139.470 167.155 ;
        RECT 142.930 166.965 143.310 167.155 ;
        RECT 146.770 166.965 147.150 167.155 ;
        RECT 150.610 166.965 150.990 167.155 ;
        RECT 154.450 166.965 154.830 167.155 ;
        RECT 158.290 166.965 158.670 167.155 ;
        RECT 28.390 166.155 166.790 166.965 ;
        RECT 25.200 164.340 25.580 164.720 ;
        RECT 28.390 164.705 29.200 166.155 ;
        RECT 161.300 165.965 161.680 166.155 ;
        RECT 163.340 165.965 163.720 166.155 ;
        RECT 165.380 165.965 165.760 166.155 ;
        RECT 161.300 164.705 161.680 164.895 ;
        RECT 163.340 164.705 163.720 164.895 ;
        RECT 165.380 164.705 165.760 164.895 ;
        RECT 28.390 163.895 166.790 164.705 ;
        RECT 32.140 163.705 32.520 163.895 ;
        RECT 35.980 163.705 36.360 163.895 ;
        RECT 39.820 163.705 40.200 163.895 ;
        RECT 43.660 163.705 44.040 163.895 ;
        RECT 47.500 163.705 47.880 163.895 ;
        RECT 51.340 163.705 51.720 163.895 ;
        RECT 55.180 163.705 55.560 163.895 ;
        RECT 59.020 163.705 59.400 163.895 ;
        RECT 64.590 163.705 64.970 163.895 ;
        RECT 68.430 163.705 68.810 163.895 ;
        RECT 72.270 163.705 72.650 163.895 ;
        RECT 76.110 163.705 76.490 163.895 ;
        RECT 79.950 163.705 80.330 163.895 ;
        RECT 83.790 163.705 84.170 163.895 ;
        RECT 87.630 163.705 88.010 163.895 ;
        RECT 91.470 163.705 91.850 163.895 ;
        RECT 97.040 163.705 97.420 163.895 ;
        RECT 100.880 163.705 101.260 163.895 ;
        RECT 104.720 163.705 105.100 163.895 ;
        RECT 108.560 163.705 108.940 163.895 ;
        RECT 112.400 163.705 112.780 163.895 ;
        RECT 116.240 163.705 116.620 163.895 ;
        RECT 120.080 163.705 120.460 163.895 ;
        RECT 123.920 163.705 124.300 163.895 ;
        RECT 129.490 163.705 129.870 163.895 ;
        RECT 133.330 163.705 133.710 163.895 ;
        RECT 137.170 163.705 137.550 163.895 ;
        RECT 141.010 163.705 141.390 163.895 ;
        RECT 144.850 163.705 145.230 163.895 ;
        RECT 148.690 163.705 149.070 163.895 ;
        RECT 152.530 163.705 152.910 163.895 ;
        RECT 156.370 163.705 156.750 163.895 ;
        RECT 25.200 161.340 25.580 161.720 ;
        RECT 27.480 159.005 27.830 163.195 ;
        RECT 25.200 158.340 25.580 158.720 ;
        RECT 28.110 157.650 28.460 161.565 ;
        RECT 29.120 161.340 29.500 161.720 ;
        RECT 31.920 160.375 34.160 160.755 ;
        RECT 37.215 159.655 38.965 163.510 ;
        RECT 29.120 158.340 29.500 158.720 ;
        RECT 31.920 158.535 34.160 158.915 ;
        RECT 41.055 157.810 42.805 163.510 ;
        RECT 27.705 157.325 28.460 157.650 ;
        RECT 28.110 157.320 28.460 157.325 ;
        RECT 31.920 156.690 34.160 157.070 ;
        RECT 31.925 155.930 34.165 156.310 ;
        RECT 25.200 155.340 25.580 155.720 ;
        RECT 29.120 155.340 29.500 155.720 ;
        RECT 44.895 155.170 46.645 163.510 ;
        RECT 31.920 154.050 34.160 154.430 ;
        RECT 48.735 153.330 50.485 163.510 ;
        RECT 25.200 152.340 25.580 152.720 ;
        RECT 29.120 152.340 29.500 152.720 ;
        RECT 31.920 152.210 34.160 152.590 ;
        RECT 52.575 151.485 54.325 163.510 ;
        RECT 31.920 150.365 34.160 150.745 ;
        RECT 25.200 149.340 25.580 149.720 ;
        RECT 29.120 149.340 29.500 149.720 ;
        RECT 31.925 149.605 34.165 149.985 ;
        RECT 56.415 148.845 58.165 163.510 ;
        RECT 31.920 147.725 34.160 148.105 ;
        RECT 60.255 147.005 62.005 163.510 ;
        RECT 62.520 160.935 62.900 161.315 ;
        RECT 64.370 160.375 66.610 160.755 ;
        RECT 69.665 159.655 71.415 163.510 ;
        RECT 62.520 159.095 62.900 159.475 ;
        RECT 64.370 158.535 66.610 158.915 ;
        RECT 73.505 157.810 75.255 163.510 ;
        RECT 62.520 157.250 62.900 157.630 ;
        RECT 64.370 156.690 66.610 157.070 ;
        RECT 64.375 155.930 66.615 156.310 ;
        RECT 77.345 155.170 79.095 163.510 ;
        RECT 62.520 154.610 62.900 154.990 ;
        RECT 64.370 154.050 66.610 154.430 ;
        RECT 81.185 153.330 82.935 163.510 ;
        RECT 62.520 152.770 62.900 153.150 ;
        RECT 64.370 152.210 66.610 152.590 ;
        RECT 85.025 151.485 86.775 163.510 ;
        RECT 62.520 150.925 62.900 151.305 ;
        RECT 64.370 150.365 66.610 150.745 ;
        RECT 64.375 149.605 66.615 149.985 ;
        RECT 88.865 148.845 90.615 163.510 ;
        RECT 62.520 148.285 62.900 148.665 ;
        RECT 64.370 147.725 66.610 148.105 ;
        RECT 92.705 147.005 94.455 163.510 ;
        RECT 94.970 160.935 95.350 161.315 ;
        RECT 96.820 160.375 99.060 160.755 ;
        RECT 102.115 159.655 103.865 163.510 ;
        RECT 94.970 159.095 95.350 159.475 ;
        RECT 96.820 158.535 99.060 158.915 ;
        RECT 105.955 157.810 107.705 163.510 ;
        RECT 94.970 157.250 95.350 157.630 ;
        RECT 96.820 156.690 99.060 157.070 ;
        RECT 96.825 155.930 99.065 156.310 ;
        RECT 109.795 155.170 111.545 163.510 ;
        RECT 94.970 154.610 95.350 154.990 ;
        RECT 96.820 154.050 99.060 154.430 ;
        RECT 113.635 153.330 115.385 163.510 ;
        RECT 94.970 152.770 95.350 153.150 ;
        RECT 96.820 152.210 99.060 152.590 ;
        RECT 117.475 151.485 119.225 163.510 ;
        RECT 94.970 150.925 95.350 151.305 ;
        RECT 96.820 150.365 99.060 150.745 ;
        RECT 96.825 149.605 99.065 149.985 ;
        RECT 121.315 148.845 123.065 163.510 ;
        RECT 94.970 148.285 95.350 148.665 ;
        RECT 96.820 147.725 99.060 148.105 ;
        RECT 125.155 147.005 126.905 163.510 ;
        RECT 127.420 160.935 127.800 161.315 ;
        RECT 129.270 160.375 131.510 160.755 ;
        RECT 134.565 159.655 136.315 163.510 ;
        RECT 127.420 159.095 127.800 159.475 ;
        RECT 129.270 158.535 131.510 158.915 ;
        RECT 138.405 157.810 140.155 163.510 ;
        RECT 127.420 157.250 127.800 157.630 ;
        RECT 129.270 156.690 131.510 157.070 ;
        RECT 129.275 155.930 131.515 156.310 ;
        RECT 142.245 155.170 143.995 163.510 ;
        RECT 127.420 154.610 127.800 154.990 ;
        RECT 129.270 154.050 131.510 154.430 ;
        RECT 146.085 153.330 147.835 163.510 ;
        RECT 127.420 152.770 127.800 153.150 ;
        RECT 129.270 152.210 131.510 152.590 ;
        RECT 149.925 151.485 151.675 163.510 ;
        RECT 127.420 150.925 127.800 151.305 ;
        RECT 129.270 150.365 131.510 150.745 ;
        RECT 129.275 149.605 131.515 149.985 ;
        RECT 153.765 148.845 155.515 163.510 ;
        RECT 127.420 148.285 127.800 148.665 ;
        RECT 129.270 147.725 131.510 148.105 ;
        RECT 157.605 147.005 159.355 163.510 ;
        RECT 162.315 162.840 162.695 163.220 ;
        RECT 164.355 162.840 164.735 163.220 ;
        RECT 166.140 162.840 166.520 163.220 ;
        RECT 159.870 160.935 160.250 161.315 ;
        RECT 162.315 159.840 162.695 160.220 ;
        RECT 164.355 159.840 164.735 160.220 ;
        RECT 166.140 159.840 166.520 160.220 ;
        RECT 159.870 159.095 160.250 159.475 ;
        RECT 159.870 157.250 160.250 157.630 ;
        RECT 162.315 156.840 162.695 157.220 ;
        RECT 164.355 156.840 164.735 157.220 ;
        RECT 166.140 156.840 166.520 157.220 ;
        RECT 159.870 154.610 160.250 154.990 ;
        RECT 162.315 153.840 162.695 154.220 ;
        RECT 164.355 153.840 164.735 154.220 ;
        RECT 166.140 153.840 166.520 154.220 ;
        RECT 159.870 152.770 160.250 153.150 ;
        RECT 159.870 150.925 160.250 151.305 ;
        RECT 162.315 150.840 162.695 151.220 ;
        RECT 164.355 150.840 164.735 151.220 ;
        RECT 166.140 150.840 166.520 151.220 ;
        RECT 159.870 148.285 160.250 148.665 ;
        RECT 162.315 147.840 162.695 148.220 ;
        RECT 164.355 147.840 164.735 148.220 ;
        RECT 166.140 147.840 166.520 148.220 ;
        RECT 25.200 146.340 25.580 146.720 ;
        RECT 29.120 146.340 29.500 146.720 ;
        RECT 62.520 146.445 62.900 146.825 ;
        RECT 94.970 146.445 95.350 146.825 ;
        RECT 127.420 146.445 127.800 146.825 ;
        RECT 159.870 146.445 160.250 146.825 ;
        RECT 31.920 145.885 34.160 146.265 ;
        RECT 64.370 145.885 66.610 146.265 ;
        RECT 96.820 145.885 99.060 146.265 ;
        RECT 129.270 145.885 131.510 146.265 ;
        RECT 31.920 145.165 34.160 145.545 ;
        RECT 64.370 145.165 66.610 145.545 ;
        RECT 96.820 145.165 99.060 145.545 ;
        RECT 129.270 145.165 131.510 145.545 ;
        RECT 62.520 144.605 62.900 144.985 ;
        RECT 94.970 144.605 95.350 144.985 ;
        RECT 127.420 144.605 127.800 144.985 ;
        RECT 159.870 144.605 160.250 144.985 ;
        RECT 25.200 142.955 25.580 143.335 ;
        RECT 29.120 142.955 29.500 143.335 ;
        RECT 31.920 143.325 34.160 143.705 ;
        RECT 31.925 141.440 34.165 141.820 ;
        RECT 31.920 140.680 34.160 141.060 ;
        RECT 25.200 139.955 25.580 140.335 ;
        RECT 29.120 139.955 29.500 140.335 ;
        RECT 31.920 138.840 34.160 139.220 ;
        RECT 25.200 136.955 25.580 137.335 ;
        RECT 29.120 136.955 29.500 137.335 ;
        RECT 31.920 137.000 34.160 137.380 ;
        RECT 31.925 135.115 34.165 135.495 ;
        RECT 31.920 134.355 34.160 134.735 ;
        RECT 25.200 133.955 25.580 134.335 ;
        RECT 29.120 133.955 29.500 134.335 ;
        RECT 31.920 132.515 34.160 132.895 ;
        RECT 25.200 130.955 25.580 131.335 ;
        RECT 29.120 130.955 29.500 131.335 ;
        RECT 31.920 130.675 34.160 131.055 ;
        RECT 25.200 127.955 25.580 128.335 ;
        RECT 29.120 127.955 29.500 128.335 ;
        RECT 35.295 127.965 37.045 131.775 ;
        RECT 39.135 127.965 40.885 133.615 ;
        RECT 42.975 127.965 44.725 136.260 ;
        RECT 46.815 127.965 48.565 138.100 ;
        RECT 50.655 127.965 52.405 139.940 ;
        RECT 54.495 127.965 56.245 142.585 ;
        RECT 58.335 127.965 60.085 144.425 ;
        RECT 64.370 143.325 66.610 143.705 ;
        RECT 62.520 142.765 62.900 143.145 ;
        RECT 64.375 141.440 66.615 141.820 ;
        RECT 64.370 140.680 66.610 141.060 ;
        RECT 62.520 140.120 62.900 140.500 ;
        RECT 64.370 138.840 66.610 139.220 ;
        RECT 62.520 138.280 62.900 138.660 ;
        RECT 64.370 137.000 66.610 137.380 ;
        RECT 62.520 136.440 62.900 136.820 ;
        RECT 64.375 135.115 66.615 135.495 ;
        RECT 64.370 134.355 66.610 134.735 ;
        RECT 62.520 133.795 62.900 134.175 ;
        RECT 64.370 132.515 66.610 132.895 ;
        RECT 62.520 131.955 62.900 132.335 ;
        RECT 64.370 130.675 66.610 131.055 ;
        RECT 62.520 130.115 62.900 130.495 ;
        RECT 67.745 127.965 69.495 131.775 ;
        RECT 71.585 127.965 73.335 133.615 ;
        RECT 75.425 127.965 77.175 136.260 ;
        RECT 79.265 127.965 81.015 138.100 ;
        RECT 83.105 127.965 84.855 139.940 ;
        RECT 86.945 127.965 88.695 142.585 ;
        RECT 90.785 127.965 92.535 144.425 ;
        RECT 96.820 143.325 99.060 143.705 ;
        RECT 94.970 142.765 95.350 143.145 ;
        RECT 96.825 141.440 99.065 141.820 ;
        RECT 96.820 140.680 99.060 141.060 ;
        RECT 94.970 140.120 95.350 140.500 ;
        RECT 96.820 138.840 99.060 139.220 ;
        RECT 94.970 138.280 95.350 138.660 ;
        RECT 96.820 137.000 99.060 137.380 ;
        RECT 94.970 136.440 95.350 136.820 ;
        RECT 96.825 135.115 99.065 135.495 ;
        RECT 96.820 134.355 99.060 134.735 ;
        RECT 94.970 133.795 95.350 134.175 ;
        RECT 96.820 132.515 99.060 132.895 ;
        RECT 94.970 131.955 95.350 132.335 ;
        RECT 96.820 130.675 99.060 131.055 ;
        RECT 94.970 130.115 95.350 130.495 ;
        RECT 100.195 127.965 101.945 131.775 ;
        RECT 104.035 127.965 105.785 133.615 ;
        RECT 107.875 127.965 109.625 136.260 ;
        RECT 111.715 127.965 113.465 138.100 ;
        RECT 115.555 127.965 117.305 139.940 ;
        RECT 119.395 127.965 121.145 142.585 ;
        RECT 123.235 127.965 124.985 144.425 ;
        RECT 129.270 143.325 131.510 143.705 ;
        RECT 127.420 142.765 127.800 143.145 ;
        RECT 129.275 141.440 131.515 141.820 ;
        RECT 129.270 140.680 131.510 141.060 ;
        RECT 127.420 140.120 127.800 140.500 ;
        RECT 129.270 138.840 131.510 139.220 ;
        RECT 127.420 138.280 127.800 138.660 ;
        RECT 129.270 137.000 131.510 137.380 ;
        RECT 127.420 136.440 127.800 136.820 ;
        RECT 129.275 135.115 131.515 135.495 ;
        RECT 129.270 134.355 131.510 134.735 ;
        RECT 127.420 133.795 127.800 134.175 ;
        RECT 129.270 132.515 131.510 132.895 ;
        RECT 127.420 131.955 127.800 132.335 ;
        RECT 129.270 130.675 131.510 131.055 ;
        RECT 127.420 130.115 127.800 130.495 ;
        RECT 132.645 127.965 134.395 131.775 ;
        RECT 136.485 127.965 138.235 133.615 ;
        RECT 140.325 127.965 142.075 136.260 ;
        RECT 144.165 127.965 145.915 138.100 ;
        RECT 148.005 127.965 149.755 139.940 ;
        RECT 151.845 127.965 153.595 142.585 ;
        RECT 155.685 127.965 157.435 144.425 ;
        RECT 159.870 142.765 160.250 143.145 ;
        RECT 162.315 141.455 162.695 141.835 ;
        RECT 164.355 141.455 164.735 141.835 ;
        RECT 166.140 141.455 166.520 141.835 ;
        RECT 159.870 140.120 160.250 140.500 ;
        RECT 159.870 138.280 160.250 138.660 ;
        RECT 162.315 138.455 162.695 138.835 ;
        RECT 164.355 138.455 164.735 138.835 ;
        RECT 166.140 138.455 166.520 138.835 ;
        RECT 159.870 136.440 160.250 136.820 ;
        RECT 162.315 135.455 162.695 135.835 ;
        RECT 164.355 135.455 164.735 135.835 ;
        RECT 166.140 135.455 166.520 135.835 ;
        RECT 159.870 133.795 160.250 134.175 ;
        RECT 162.315 132.455 162.695 132.835 ;
        RECT 164.355 132.455 164.735 132.835 ;
        RECT 166.140 132.455 166.520 132.835 ;
        RECT 159.870 131.955 160.250 132.335 ;
        RECT 159.870 130.115 160.250 130.495 ;
        RECT 162.315 129.455 162.695 129.835 ;
        RECT 164.355 129.455 164.735 129.835 ;
        RECT 166.140 129.455 166.520 129.835 ;
        RECT 34.060 127.580 34.440 127.770 ;
        RECT 37.900 127.580 38.280 127.770 ;
        RECT 41.740 127.580 42.120 127.770 ;
        RECT 45.580 127.580 45.960 127.770 ;
        RECT 49.420 127.580 49.800 127.770 ;
        RECT 53.260 127.580 53.640 127.770 ;
        RECT 57.100 127.580 57.480 127.770 ;
        RECT 60.940 127.580 61.320 127.770 ;
        RECT 66.510 127.580 66.890 127.770 ;
        RECT 70.350 127.580 70.730 127.770 ;
        RECT 74.190 127.580 74.570 127.770 ;
        RECT 78.030 127.580 78.410 127.770 ;
        RECT 81.870 127.580 82.250 127.770 ;
        RECT 85.710 127.580 86.090 127.770 ;
        RECT 89.550 127.580 89.930 127.770 ;
        RECT 93.390 127.580 93.770 127.770 ;
        RECT 98.960 127.580 99.340 127.770 ;
        RECT 102.800 127.580 103.180 127.770 ;
        RECT 106.640 127.580 107.020 127.770 ;
        RECT 110.480 127.580 110.860 127.770 ;
        RECT 114.320 127.580 114.700 127.770 ;
        RECT 118.160 127.580 118.540 127.770 ;
        RECT 122.000 127.580 122.380 127.770 ;
        RECT 125.840 127.580 126.220 127.770 ;
        RECT 131.410 127.580 131.790 127.770 ;
        RECT 135.250 127.580 135.630 127.770 ;
        RECT 139.090 127.580 139.470 127.770 ;
        RECT 142.930 127.580 143.310 127.770 ;
        RECT 146.770 127.580 147.150 127.770 ;
        RECT 150.610 127.580 150.990 127.770 ;
        RECT 154.450 127.580 154.830 127.770 ;
        RECT 158.290 127.580 158.670 127.770 ;
        RECT 28.390 126.770 166.790 127.580 ;
        RECT 25.200 124.955 25.580 125.335 ;
        RECT 28.390 125.320 29.200 126.770 ;
        RECT 161.300 126.580 161.680 126.770 ;
        RECT 163.340 126.580 163.720 126.770 ;
        RECT 165.380 126.580 165.760 126.770 ;
        RECT 161.300 125.320 161.680 125.510 ;
        RECT 163.340 125.320 163.720 125.510 ;
        RECT 165.380 125.320 165.760 125.510 ;
        RECT 28.390 124.510 166.790 125.320 ;
        RECT 32.140 124.320 32.520 124.510 ;
        RECT 35.980 124.320 36.360 124.510 ;
        RECT 39.820 124.320 40.200 124.510 ;
        RECT 43.660 124.320 44.040 124.510 ;
        RECT 47.500 124.320 47.880 124.510 ;
        RECT 51.340 124.320 51.720 124.510 ;
        RECT 55.180 124.320 55.560 124.510 ;
        RECT 59.020 124.320 59.400 124.510 ;
        RECT 64.590 124.320 64.970 124.510 ;
        RECT 68.430 124.320 68.810 124.510 ;
        RECT 72.270 124.320 72.650 124.510 ;
        RECT 76.110 124.320 76.490 124.510 ;
        RECT 79.950 124.320 80.330 124.510 ;
        RECT 83.790 124.320 84.170 124.510 ;
        RECT 87.630 124.320 88.010 124.510 ;
        RECT 91.470 124.320 91.850 124.510 ;
        RECT 97.040 124.320 97.420 124.510 ;
        RECT 100.880 124.320 101.260 124.510 ;
        RECT 104.720 124.320 105.100 124.510 ;
        RECT 108.560 124.320 108.940 124.510 ;
        RECT 112.400 124.320 112.780 124.510 ;
        RECT 116.240 124.320 116.620 124.510 ;
        RECT 120.080 124.320 120.460 124.510 ;
        RECT 123.920 124.320 124.300 124.510 ;
        RECT 129.490 124.320 129.870 124.510 ;
        RECT 133.330 124.320 133.710 124.510 ;
        RECT 137.170 124.320 137.550 124.510 ;
        RECT 141.010 124.320 141.390 124.510 ;
        RECT 144.850 124.320 145.230 124.510 ;
        RECT 148.690 124.320 149.070 124.510 ;
        RECT 152.530 124.320 152.910 124.510 ;
        RECT 156.370 124.320 156.750 124.510 ;
        RECT 25.200 121.955 25.580 122.335 ;
        RECT 27.480 119.620 27.830 123.810 ;
        RECT 25.200 118.955 25.580 119.335 ;
        RECT 28.110 118.265 28.460 122.180 ;
        RECT 29.120 121.955 29.500 122.335 ;
        RECT 31.920 120.990 34.160 121.370 ;
        RECT 37.215 120.270 38.965 124.125 ;
        RECT 29.120 118.955 29.500 119.335 ;
        RECT 31.920 119.150 34.160 119.530 ;
        RECT 41.055 118.425 42.805 124.125 ;
        RECT 27.705 117.940 28.460 118.265 ;
        RECT 28.110 117.935 28.460 117.940 ;
        RECT 31.920 117.305 34.160 117.685 ;
        RECT 31.925 116.545 34.165 116.925 ;
        RECT 25.200 115.955 25.580 116.335 ;
        RECT 29.120 115.955 29.500 116.335 ;
        RECT 44.895 115.785 46.645 124.125 ;
        RECT 31.920 114.665 34.160 115.045 ;
        RECT 48.735 113.945 50.485 124.125 ;
        RECT 25.200 112.955 25.580 113.335 ;
        RECT 29.120 112.955 29.500 113.335 ;
        RECT 31.920 112.825 34.160 113.205 ;
        RECT 52.575 112.100 54.325 124.125 ;
        RECT 31.920 110.980 34.160 111.360 ;
        RECT 25.200 109.955 25.580 110.335 ;
        RECT 29.120 109.955 29.500 110.335 ;
        RECT 31.925 110.220 34.165 110.600 ;
        RECT 56.415 109.460 58.165 124.125 ;
        RECT 31.920 108.340 34.160 108.720 ;
        RECT 60.255 107.620 62.005 124.125 ;
        RECT 62.520 121.550 62.900 121.930 ;
        RECT 64.370 120.990 66.610 121.370 ;
        RECT 69.665 120.270 71.415 124.125 ;
        RECT 62.520 119.710 62.900 120.090 ;
        RECT 64.370 119.150 66.610 119.530 ;
        RECT 73.505 118.425 75.255 124.125 ;
        RECT 62.520 117.865 62.900 118.245 ;
        RECT 64.370 117.305 66.610 117.685 ;
        RECT 64.375 116.545 66.615 116.925 ;
        RECT 77.345 115.785 79.095 124.125 ;
        RECT 62.520 115.225 62.900 115.605 ;
        RECT 64.370 114.665 66.610 115.045 ;
        RECT 81.185 113.945 82.935 124.125 ;
        RECT 62.520 113.385 62.900 113.765 ;
        RECT 64.370 112.825 66.610 113.205 ;
        RECT 85.025 112.100 86.775 124.125 ;
        RECT 62.520 111.540 62.900 111.920 ;
        RECT 64.370 110.980 66.610 111.360 ;
        RECT 64.375 110.220 66.615 110.600 ;
        RECT 88.865 109.460 90.615 124.125 ;
        RECT 62.520 108.900 62.900 109.280 ;
        RECT 64.370 108.340 66.610 108.720 ;
        RECT 92.705 107.620 94.455 124.125 ;
        RECT 94.970 121.550 95.350 121.930 ;
        RECT 96.820 120.990 99.060 121.370 ;
        RECT 102.115 120.270 103.865 124.125 ;
        RECT 94.970 119.710 95.350 120.090 ;
        RECT 96.820 119.150 99.060 119.530 ;
        RECT 105.955 118.425 107.705 124.125 ;
        RECT 94.970 117.865 95.350 118.245 ;
        RECT 96.820 117.305 99.060 117.685 ;
        RECT 96.825 116.545 99.065 116.925 ;
        RECT 109.795 115.785 111.545 124.125 ;
        RECT 94.970 115.225 95.350 115.605 ;
        RECT 96.820 114.665 99.060 115.045 ;
        RECT 113.635 113.945 115.385 124.125 ;
        RECT 94.970 113.385 95.350 113.765 ;
        RECT 96.820 112.825 99.060 113.205 ;
        RECT 117.475 112.100 119.225 124.125 ;
        RECT 94.970 111.540 95.350 111.920 ;
        RECT 96.820 110.980 99.060 111.360 ;
        RECT 96.825 110.220 99.065 110.600 ;
        RECT 121.315 109.460 123.065 124.125 ;
        RECT 94.970 108.900 95.350 109.280 ;
        RECT 96.820 108.340 99.060 108.720 ;
        RECT 125.155 107.620 126.905 124.125 ;
        RECT 127.420 121.550 127.800 121.930 ;
        RECT 129.270 120.990 131.510 121.370 ;
        RECT 134.565 120.270 136.315 124.125 ;
        RECT 127.420 119.710 127.800 120.090 ;
        RECT 129.270 119.150 131.510 119.530 ;
        RECT 138.405 118.425 140.155 124.125 ;
        RECT 127.420 117.865 127.800 118.245 ;
        RECT 129.270 117.305 131.510 117.685 ;
        RECT 129.275 116.545 131.515 116.925 ;
        RECT 142.245 115.785 143.995 124.125 ;
        RECT 127.420 115.225 127.800 115.605 ;
        RECT 129.270 114.665 131.510 115.045 ;
        RECT 146.085 113.945 147.835 124.125 ;
        RECT 127.420 113.385 127.800 113.765 ;
        RECT 129.270 112.825 131.510 113.205 ;
        RECT 149.925 112.100 151.675 124.125 ;
        RECT 127.420 111.540 127.800 111.920 ;
        RECT 129.270 110.980 131.510 111.360 ;
        RECT 129.275 110.220 131.515 110.600 ;
        RECT 153.765 109.460 155.515 124.125 ;
        RECT 127.420 108.900 127.800 109.280 ;
        RECT 129.270 108.340 131.510 108.720 ;
        RECT 157.605 107.620 159.355 124.125 ;
        RECT 162.315 123.455 162.695 123.835 ;
        RECT 164.355 123.455 164.735 123.835 ;
        RECT 166.140 123.455 166.520 123.835 ;
        RECT 159.870 121.550 160.250 121.930 ;
        RECT 162.315 120.455 162.695 120.835 ;
        RECT 164.355 120.455 164.735 120.835 ;
        RECT 166.140 120.455 166.520 120.835 ;
        RECT 159.870 119.710 160.250 120.090 ;
        RECT 159.870 117.865 160.250 118.245 ;
        RECT 162.315 117.455 162.695 117.835 ;
        RECT 164.355 117.455 164.735 117.835 ;
        RECT 166.140 117.455 166.520 117.835 ;
        RECT 159.870 115.225 160.250 115.605 ;
        RECT 162.315 114.455 162.695 114.835 ;
        RECT 164.355 114.455 164.735 114.835 ;
        RECT 166.140 114.455 166.520 114.835 ;
        RECT 159.870 113.385 160.250 113.765 ;
        RECT 159.870 111.540 160.250 111.920 ;
        RECT 162.315 111.455 162.695 111.835 ;
        RECT 164.355 111.455 164.735 111.835 ;
        RECT 166.140 111.455 166.520 111.835 ;
        RECT 159.870 108.900 160.250 109.280 ;
        RECT 162.315 108.455 162.695 108.835 ;
        RECT 164.355 108.455 164.735 108.835 ;
        RECT 166.140 108.455 166.520 108.835 ;
        RECT 25.200 106.955 25.580 107.335 ;
        RECT 29.120 106.955 29.500 107.335 ;
        RECT 62.520 107.060 62.900 107.440 ;
        RECT 94.970 107.060 95.350 107.440 ;
        RECT 127.420 107.060 127.800 107.440 ;
        RECT 159.870 107.060 160.250 107.440 ;
        RECT 31.920 106.500 34.160 106.880 ;
        RECT 64.370 106.500 66.610 106.880 ;
        RECT 96.820 106.500 99.060 106.880 ;
        RECT 129.270 106.500 131.510 106.880 ;
        RECT 31.920 105.780 34.160 106.160 ;
        RECT 64.370 105.780 66.610 106.160 ;
        RECT 96.820 105.780 99.060 106.160 ;
        RECT 129.270 105.780 131.510 106.160 ;
        RECT 62.520 105.220 62.900 105.600 ;
        RECT 94.970 105.220 95.350 105.600 ;
        RECT 127.420 105.220 127.800 105.600 ;
        RECT 159.870 105.220 160.250 105.600 ;
        RECT 25.200 103.570 25.580 103.950 ;
        RECT 29.120 103.570 29.500 103.950 ;
        RECT 31.920 103.940 34.160 104.320 ;
        RECT 31.925 102.055 34.165 102.435 ;
        RECT 31.920 101.295 34.160 101.675 ;
        RECT 25.200 100.570 25.580 100.950 ;
        RECT 29.120 100.570 29.500 100.950 ;
        RECT 31.920 99.455 34.160 99.835 ;
        RECT 25.200 97.570 25.580 97.950 ;
        RECT 29.120 97.570 29.500 97.950 ;
        RECT 31.920 97.615 34.160 97.995 ;
        RECT 31.925 95.730 34.165 96.110 ;
        RECT 31.920 94.970 34.160 95.350 ;
        RECT 25.200 94.570 25.580 94.950 ;
        RECT 29.120 94.570 29.500 94.950 ;
        RECT 31.920 93.130 34.160 93.510 ;
        RECT 25.200 91.570 25.580 91.950 ;
        RECT 29.120 91.570 29.500 91.950 ;
        RECT 31.920 91.290 34.160 91.670 ;
        RECT 25.200 88.570 25.580 88.950 ;
        RECT 29.120 88.570 29.500 88.950 ;
        RECT 35.295 88.580 37.045 92.390 ;
        RECT 39.135 88.580 40.885 94.230 ;
        RECT 42.975 88.580 44.725 96.875 ;
        RECT 46.815 88.580 48.565 98.715 ;
        RECT 50.655 88.580 52.405 100.555 ;
        RECT 54.495 88.580 56.245 103.200 ;
        RECT 58.335 88.580 60.085 105.040 ;
        RECT 64.370 103.940 66.610 104.320 ;
        RECT 62.520 103.380 62.900 103.760 ;
        RECT 64.375 102.055 66.615 102.435 ;
        RECT 64.370 101.295 66.610 101.675 ;
        RECT 62.520 100.735 62.900 101.115 ;
        RECT 64.370 99.455 66.610 99.835 ;
        RECT 62.520 98.895 62.900 99.275 ;
        RECT 64.370 97.615 66.610 97.995 ;
        RECT 62.520 97.055 62.900 97.435 ;
        RECT 64.375 95.730 66.615 96.110 ;
        RECT 64.370 94.970 66.610 95.350 ;
        RECT 62.520 94.410 62.900 94.790 ;
        RECT 64.370 93.130 66.610 93.510 ;
        RECT 62.520 92.570 62.900 92.950 ;
        RECT 64.370 91.290 66.610 91.670 ;
        RECT 62.520 90.730 62.900 91.110 ;
        RECT 67.745 88.580 69.495 92.390 ;
        RECT 71.585 88.580 73.335 94.230 ;
        RECT 75.425 88.580 77.175 96.875 ;
        RECT 79.265 88.580 81.015 98.715 ;
        RECT 83.105 88.580 84.855 100.555 ;
        RECT 86.945 88.580 88.695 103.200 ;
        RECT 90.785 88.580 92.535 105.040 ;
        RECT 96.820 103.940 99.060 104.320 ;
        RECT 94.970 103.380 95.350 103.760 ;
        RECT 96.825 102.055 99.065 102.435 ;
        RECT 96.820 101.295 99.060 101.675 ;
        RECT 94.970 100.735 95.350 101.115 ;
        RECT 96.820 99.455 99.060 99.835 ;
        RECT 94.970 98.895 95.350 99.275 ;
        RECT 96.820 97.615 99.060 97.995 ;
        RECT 94.970 97.055 95.350 97.435 ;
        RECT 96.825 95.730 99.065 96.110 ;
        RECT 96.820 94.970 99.060 95.350 ;
        RECT 94.970 94.410 95.350 94.790 ;
        RECT 96.820 93.130 99.060 93.510 ;
        RECT 94.970 92.570 95.350 92.950 ;
        RECT 96.820 91.290 99.060 91.670 ;
        RECT 94.970 90.730 95.350 91.110 ;
        RECT 100.195 88.580 101.945 92.390 ;
        RECT 104.035 88.580 105.785 94.230 ;
        RECT 107.875 88.580 109.625 96.875 ;
        RECT 111.715 88.580 113.465 98.715 ;
        RECT 115.555 88.580 117.305 100.555 ;
        RECT 119.395 88.580 121.145 103.200 ;
        RECT 123.235 88.580 124.985 105.040 ;
        RECT 129.270 103.940 131.510 104.320 ;
        RECT 127.420 103.380 127.800 103.760 ;
        RECT 129.275 102.055 131.515 102.435 ;
        RECT 129.270 101.295 131.510 101.675 ;
        RECT 127.420 100.735 127.800 101.115 ;
        RECT 129.270 99.455 131.510 99.835 ;
        RECT 127.420 98.895 127.800 99.275 ;
        RECT 129.270 97.615 131.510 97.995 ;
        RECT 127.420 97.055 127.800 97.435 ;
        RECT 129.275 95.730 131.515 96.110 ;
        RECT 129.270 94.970 131.510 95.350 ;
        RECT 127.420 94.410 127.800 94.790 ;
        RECT 129.270 93.130 131.510 93.510 ;
        RECT 127.420 92.570 127.800 92.950 ;
        RECT 129.270 91.290 131.510 91.670 ;
        RECT 127.420 90.730 127.800 91.110 ;
        RECT 132.645 88.580 134.395 92.390 ;
        RECT 136.485 88.580 138.235 94.230 ;
        RECT 140.325 88.580 142.075 96.875 ;
        RECT 144.165 88.580 145.915 98.715 ;
        RECT 148.005 88.580 149.755 100.555 ;
        RECT 151.845 88.580 153.595 103.200 ;
        RECT 155.685 88.580 157.435 105.040 ;
        RECT 159.870 103.380 160.250 103.760 ;
        RECT 162.315 102.070 162.695 102.450 ;
        RECT 164.355 102.070 164.735 102.450 ;
        RECT 166.140 102.070 166.520 102.450 ;
        RECT 159.870 100.735 160.250 101.115 ;
        RECT 159.870 98.895 160.250 99.275 ;
        RECT 162.315 99.070 162.695 99.450 ;
        RECT 164.355 99.070 164.735 99.450 ;
        RECT 166.140 99.070 166.520 99.450 ;
        RECT 159.870 97.055 160.250 97.435 ;
        RECT 162.315 96.070 162.695 96.450 ;
        RECT 164.355 96.070 164.735 96.450 ;
        RECT 166.140 96.070 166.520 96.450 ;
        RECT 159.870 94.410 160.250 94.790 ;
        RECT 162.315 93.070 162.695 93.450 ;
        RECT 164.355 93.070 164.735 93.450 ;
        RECT 166.140 93.070 166.520 93.450 ;
        RECT 159.870 92.570 160.250 92.950 ;
        RECT 159.870 90.730 160.250 91.110 ;
        RECT 162.315 90.070 162.695 90.450 ;
        RECT 164.355 90.070 164.735 90.450 ;
        RECT 166.140 90.070 166.520 90.450 ;
        RECT 34.060 88.195 34.440 88.385 ;
        RECT 37.900 88.195 38.280 88.385 ;
        RECT 41.740 88.195 42.120 88.385 ;
        RECT 45.580 88.195 45.960 88.385 ;
        RECT 49.420 88.195 49.800 88.385 ;
        RECT 53.260 88.195 53.640 88.385 ;
        RECT 57.100 88.195 57.480 88.385 ;
        RECT 60.940 88.195 61.320 88.385 ;
        RECT 66.510 88.195 66.890 88.385 ;
        RECT 70.350 88.195 70.730 88.385 ;
        RECT 74.190 88.195 74.570 88.385 ;
        RECT 78.030 88.195 78.410 88.385 ;
        RECT 81.870 88.195 82.250 88.385 ;
        RECT 85.710 88.195 86.090 88.385 ;
        RECT 89.550 88.195 89.930 88.385 ;
        RECT 93.390 88.195 93.770 88.385 ;
        RECT 98.960 88.195 99.340 88.385 ;
        RECT 102.800 88.195 103.180 88.385 ;
        RECT 106.640 88.195 107.020 88.385 ;
        RECT 110.480 88.195 110.860 88.385 ;
        RECT 114.320 88.195 114.700 88.385 ;
        RECT 118.160 88.195 118.540 88.385 ;
        RECT 122.000 88.195 122.380 88.385 ;
        RECT 125.840 88.195 126.220 88.385 ;
        RECT 131.410 88.195 131.790 88.385 ;
        RECT 135.250 88.195 135.630 88.385 ;
        RECT 139.090 88.195 139.470 88.385 ;
        RECT 142.930 88.195 143.310 88.385 ;
        RECT 146.770 88.195 147.150 88.385 ;
        RECT 150.610 88.195 150.990 88.385 ;
        RECT 154.450 88.195 154.830 88.385 ;
        RECT 158.290 88.195 158.670 88.385 ;
        RECT 28.390 87.385 166.790 88.195 ;
        RECT 25.200 85.570 25.580 85.950 ;
        RECT 28.390 85.935 29.200 87.385 ;
        RECT 161.300 87.195 161.680 87.385 ;
        RECT 163.340 87.195 163.720 87.385 ;
        RECT 165.380 87.195 165.760 87.385 ;
        RECT 161.300 85.935 161.680 86.125 ;
        RECT 163.340 85.935 163.720 86.125 ;
        RECT 165.380 85.935 165.760 86.125 ;
        RECT 28.390 85.125 166.790 85.935 ;
        RECT 32.140 84.935 32.520 85.125 ;
        RECT 35.980 84.935 36.360 85.125 ;
        RECT 39.820 84.935 40.200 85.125 ;
        RECT 43.660 84.935 44.040 85.125 ;
        RECT 47.500 84.935 47.880 85.125 ;
        RECT 51.340 84.935 51.720 85.125 ;
        RECT 55.180 84.935 55.560 85.125 ;
        RECT 59.020 84.935 59.400 85.125 ;
        RECT 64.590 84.935 64.970 85.125 ;
        RECT 68.430 84.935 68.810 85.125 ;
        RECT 72.270 84.935 72.650 85.125 ;
        RECT 76.110 84.935 76.490 85.125 ;
        RECT 79.950 84.935 80.330 85.125 ;
        RECT 83.790 84.935 84.170 85.125 ;
        RECT 87.630 84.935 88.010 85.125 ;
        RECT 91.470 84.935 91.850 85.125 ;
        RECT 97.040 84.935 97.420 85.125 ;
        RECT 100.880 84.935 101.260 85.125 ;
        RECT 104.720 84.935 105.100 85.125 ;
        RECT 108.560 84.935 108.940 85.125 ;
        RECT 112.400 84.935 112.780 85.125 ;
        RECT 116.240 84.935 116.620 85.125 ;
        RECT 120.080 84.935 120.460 85.125 ;
        RECT 123.920 84.935 124.300 85.125 ;
        RECT 129.490 84.935 129.870 85.125 ;
        RECT 133.330 84.935 133.710 85.125 ;
        RECT 137.170 84.935 137.550 85.125 ;
        RECT 141.010 84.935 141.390 85.125 ;
        RECT 144.850 84.935 145.230 85.125 ;
        RECT 148.690 84.935 149.070 85.125 ;
        RECT 152.530 84.935 152.910 85.125 ;
        RECT 156.370 84.935 156.750 85.125 ;
        RECT 25.200 82.570 25.580 82.950 ;
        RECT 27.480 80.235 27.830 84.425 ;
        RECT 25.200 79.570 25.580 79.950 ;
        RECT 28.110 78.880 28.460 82.795 ;
        RECT 29.120 82.570 29.500 82.950 ;
        RECT 31.920 81.605 34.160 81.985 ;
        RECT 37.215 80.885 38.965 84.740 ;
        RECT 29.120 79.570 29.500 79.950 ;
        RECT 31.920 79.765 34.160 80.145 ;
        RECT 41.055 79.040 42.805 84.740 ;
        RECT 27.705 78.555 28.460 78.880 ;
        RECT 28.110 78.550 28.460 78.555 ;
        RECT 31.920 77.920 34.160 78.300 ;
        RECT 31.925 77.160 34.165 77.540 ;
        RECT 25.200 76.570 25.580 76.950 ;
        RECT 29.120 76.570 29.500 76.950 ;
        RECT 44.895 76.400 46.645 84.740 ;
        RECT 31.920 75.280 34.160 75.660 ;
        RECT 48.735 74.560 50.485 84.740 ;
        RECT 25.200 73.570 25.580 73.950 ;
        RECT 29.120 73.570 29.500 73.950 ;
        RECT 31.920 73.440 34.160 73.820 ;
        RECT 52.575 72.715 54.325 84.740 ;
        RECT 31.920 71.595 34.160 71.975 ;
        RECT 25.200 70.570 25.580 70.950 ;
        RECT 29.120 70.570 29.500 70.950 ;
        RECT 31.925 70.835 34.165 71.215 ;
        RECT 56.415 70.075 58.165 84.740 ;
        RECT 31.920 68.955 34.160 69.335 ;
        RECT 60.255 68.235 62.005 84.740 ;
        RECT 62.520 82.165 62.900 82.545 ;
        RECT 64.370 81.605 66.610 81.985 ;
        RECT 69.665 80.885 71.415 84.740 ;
        RECT 62.520 80.325 62.900 80.705 ;
        RECT 64.370 79.765 66.610 80.145 ;
        RECT 73.505 79.040 75.255 84.740 ;
        RECT 62.520 78.480 62.900 78.860 ;
        RECT 64.370 77.920 66.610 78.300 ;
        RECT 64.375 77.160 66.615 77.540 ;
        RECT 77.345 76.400 79.095 84.740 ;
        RECT 62.520 75.840 62.900 76.220 ;
        RECT 64.370 75.280 66.610 75.660 ;
        RECT 81.185 74.560 82.935 84.740 ;
        RECT 62.520 74.000 62.900 74.380 ;
        RECT 64.370 73.440 66.610 73.820 ;
        RECT 85.025 72.715 86.775 84.740 ;
        RECT 62.520 72.155 62.900 72.535 ;
        RECT 64.370 71.595 66.610 71.975 ;
        RECT 64.375 70.835 66.615 71.215 ;
        RECT 88.865 70.075 90.615 84.740 ;
        RECT 62.520 69.515 62.900 69.895 ;
        RECT 64.370 68.955 66.610 69.335 ;
        RECT 92.705 68.235 94.455 84.740 ;
        RECT 94.970 82.165 95.350 82.545 ;
        RECT 96.820 81.605 99.060 81.985 ;
        RECT 102.115 80.885 103.865 84.740 ;
        RECT 94.970 80.325 95.350 80.705 ;
        RECT 96.820 79.765 99.060 80.145 ;
        RECT 105.955 79.040 107.705 84.740 ;
        RECT 94.970 78.480 95.350 78.860 ;
        RECT 96.820 77.920 99.060 78.300 ;
        RECT 96.825 77.160 99.065 77.540 ;
        RECT 109.795 76.400 111.545 84.740 ;
        RECT 94.970 75.840 95.350 76.220 ;
        RECT 96.820 75.280 99.060 75.660 ;
        RECT 113.635 74.560 115.385 84.740 ;
        RECT 94.970 74.000 95.350 74.380 ;
        RECT 96.820 73.440 99.060 73.820 ;
        RECT 117.475 72.715 119.225 84.740 ;
        RECT 94.970 72.155 95.350 72.535 ;
        RECT 96.820 71.595 99.060 71.975 ;
        RECT 96.825 70.835 99.065 71.215 ;
        RECT 121.315 70.075 123.065 84.740 ;
        RECT 94.970 69.515 95.350 69.895 ;
        RECT 96.820 68.955 99.060 69.335 ;
        RECT 125.155 68.235 126.905 84.740 ;
        RECT 127.420 82.165 127.800 82.545 ;
        RECT 129.270 81.605 131.510 81.985 ;
        RECT 134.565 80.885 136.315 84.740 ;
        RECT 127.420 80.325 127.800 80.705 ;
        RECT 129.270 79.765 131.510 80.145 ;
        RECT 138.405 79.040 140.155 84.740 ;
        RECT 127.420 78.480 127.800 78.860 ;
        RECT 129.270 77.920 131.510 78.300 ;
        RECT 129.275 77.160 131.515 77.540 ;
        RECT 142.245 76.400 143.995 84.740 ;
        RECT 127.420 75.840 127.800 76.220 ;
        RECT 129.270 75.280 131.510 75.660 ;
        RECT 146.085 74.560 147.835 84.740 ;
        RECT 127.420 74.000 127.800 74.380 ;
        RECT 129.270 73.440 131.510 73.820 ;
        RECT 149.925 72.715 151.675 84.740 ;
        RECT 127.420 72.155 127.800 72.535 ;
        RECT 129.270 71.595 131.510 71.975 ;
        RECT 129.275 70.835 131.515 71.215 ;
        RECT 153.765 70.075 155.515 84.740 ;
        RECT 127.420 69.515 127.800 69.895 ;
        RECT 129.270 68.955 131.510 69.335 ;
        RECT 157.605 68.235 159.355 84.740 ;
        RECT 162.315 84.070 162.695 84.450 ;
        RECT 164.355 84.070 164.735 84.450 ;
        RECT 166.140 84.070 166.520 84.450 ;
        RECT 159.870 82.165 160.250 82.545 ;
        RECT 162.315 81.070 162.695 81.450 ;
        RECT 164.355 81.070 164.735 81.450 ;
        RECT 166.140 81.070 166.520 81.450 ;
        RECT 159.870 80.325 160.250 80.705 ;
        RECT 159.870 78.480 160.250 78.860 ;
        RECT 162.315 78.070 162.695 78.450 ;
        RECT 164.355 78.070 164.735 78.450 ;
        RECT 166.140 78.070 166.520 78.450 ;
        RECT 159.870 75.840 160.250 76.220 ;
        RECT 162.315 75.070 162.695 75.450 ;
        RECT 164.355 75.070 164.735 75.450 ;
        RECT 166.140 75.070 166.520 75.450 ;
        RECT 159.870 74.000 160.250 74.380 ;
        RECT 159.870 72.155 160.250 72.535 ;
        RECT 162.315 72.070 162.695 72.450 ;
        RECT 164.355 72.070 164.735 72.450 ;
        RECT 166.140 72.070 166.520 72.450 ;
        RECT 159.870 69.515 160.250 69.895 ;
        RECT 162.315 69.070 162.695 69.450 ;
        RECT 164.355 69.070 164.735 69.450 ;
        RECT 166.140 69.070 166.520 69.450 ;
        RECT 25.200 67.570 25.580 67.950 ;
        RECT 29.120 67.570 29.500 67.950 ;
        RECT 62.520 67.675 62.900 68.055 ;
        RECT 94.970 67.675 95.350 68.055 ;
        RECT 127.420 67.675 127.800 68.055 ;
        RECT 159.870 67.675 160.250 68.055 ;
        RECT 31.920 67.115 34.160 67.495 ;
        RECT 64.370 67.115 66.610 67.495 ;
        RECT 96.820 67.115 99.060 67.495 ;
        RECT 129.270 67.115 131.510 67.495 ;
      LAYER Metal3 ;
        RECT 31.920 381.475 34.160 381.855 ;
        RECT 64.370 381.475 66.610 381.855 ;
        RECT 96.820 381.475 99.060 381.855 ;
        RECT 129.270 381.475 131.510 381.855 ;
        RECT 53.700 381.245 54.080 381.295 ;
        RECT 62.520 381.245 62.900 381.295 ;
        RECT 53.700 380.965 62.900 381.245 ;
        RECT 53.700 380.915 54.080 380.965 ;
        RECT 62.520 380.915 62.900 380.965 ;
        RECT 86.150 381.245 86.530 381.295 ;
        RECT 94.970 381.245 95.350 381.295 ;
        RECT 86.150 380.965 95.350 381.245 ;
        RECT 86.150 380.915 86.530 380.965 ;
        RECT 94.970 380.915 95.350 380.965 ;
        RECT 118.600 381.245 118.980 381.295 ;
        RECT 127.420 381.245 127.800 381.295 ;
        RECT 118.600 380.965 127.800 381.245 ;
        RECT 118.600 380.915 118.980 380.965 ;
        RECT 127.420 380.915 127.800 380.965 ;
        RECT 151.050 381.245 151.430 381.295 ;
        RECT 159.870 381.245 160.250 381.295 ;
        RECT 151.050 380.965 160.250 381.245 ;
        RECT 151.050 380.915 151.430 380.965 ;
        RECT 159.870 380.915 160.250 380.965 ;
        RECT 25.200 379.265 25.580 379.645 ;
        RECT 29.120 379.265 29.500 379.645 ;
        RECT 31.920 379.635 34.160 380.015 ;
        RECT 64.370 379.635 66.610 380.015 ;
        RECT 96.820 379.635 99.060 380.015 ;
        RECT 129.270 379.635 131.510 380.015 ;
        RECT 54.980 379.405 55.360 379.455 ;
        RECT 62.520 379.405 62.900 379.455 ;
        RECT 54.980 379.125 62.900 379.405 ;
        RECT 54.980 379.075 55.360 379.125 ;
        RECT 62.520 379.075 62.900 379.125 ;
        RECT 87.430 379.405 87.810 379.455 ;
        RECT 94.970 379.405 95.350 379.455 ;
        RECT 87.430 379.125 95.350 379.405 ;
        RECT 87.430 379.075 87.810 379.125 ;
        RECT 94.970 379.075 95.350 379.125 ;
        RECT 119.880 379.405 120.260 379.455 ;
        RECT 127.420 379.405 127.800 379.455 ;
        RECT 119.880 379.125 127.800 379.405 ;
        RECT 119.880 379.075 120.260 379.125 ;
        RECT 127.420 379.075 127.800 379.125 ;
        RECT 152.330 379.405 152.710 379.455 ;
        RECT 159.870 379.405 160.250 379.455 ;
        RECT 152.330 379.125 160.250 379.405 ;
        RECT 152.330 379.075 152.710 379.125 ;
        RECT 159.870 379.075 160.250 379.125 ;
        RECT 31.925 377.750 34.165 378.130 ;
        RECT 64.375 377.750 66.615 378.130 ;
        RECT 96.825 377.750 99.065 378.130 ;
        RECT 129.275 377.750 131.515 378.130 ;
        RECT 162.315 377.765 162.695 378.145 ;
        RECT 164.355 377.765 164.735 378.145 ;
        RECT 166.140 377.765 166.520 378.145 ;
        RECT 31.920 376.990 34.160 377.370 ;
        RECT 64.370 376.990 66.610 377.370 ;
        RECT 96.820 376.990 99.060 377.370 ;
        RECT 129.270 376.990 131.510 377.370 ;
        RECT 56.260 376.760 56.640 376.810 ;
        RECT 62.520 376.760 62.900 376.810 ;
        RECT 25.200 376.265 25.580 376.645 ;
        RECT 29.120 376.265 29.500 376.645 ;
        RECT 56.260 376.480 62.900 376.760 ;
        RECT 56.260 376.430 56.640 376.480 ;
        RECT 62.520 376.430 62.900 376.480 ;
        RECT 88.710 376.760 89.090 376.810 ;
        RECT 94.970 376.760 95.350 376.810 ;
        RECT 88.710 376.480 95.350 376.760 ;
        RECT 88.710 376.430 89.090 376.480 ;
        RECT 94.970 376.430 95.350 376.480 ;
        RECT 121.160 376.760 121.540 376.810 ;
        RECT 127.420 376.760 127.800 376.810 ;
        RECT 121.160 376.480 127.800 376.760 ;
        RECT 121.160 376.430 121.540 376.480 ;
        RECT 127.420 376.430 127.800 376.480 ;
        RECT 153.610 376.760 153.990 376.810 ;
        RECT 159.870 376.760 160.250 376.810 ;
        RECT 153.610 376.480 160.250 376.760 ;
        RECT 153.610 376.430 153.990 376.480 ;
        RECT 159.870 376.430 160.250 376.480 ;
        RECT 31.920 375.150 34.160 375.530 ;
        RECT 64.370 375.150 66.610 375.530 ;
        RECT 96.820 375.150 99.060 375.530 ;
        RECT 129.270 375.150 131.510 375.530 ;
        RECT 57.540 374.920 57.920 374.970 ;
        RECT 62.520 374.920 62.900 374.970 ;
        RECT 57.540 374.640 62.900 374.920 ;
        RECT 57.540 374.590 57.920 374.640 ;
        RECT 62.520 374.590 62.900 374.640 ;
        RECT 89.990 374.920 90.370 374.970 ;
        RECT 94.970 374.920 95.350 374.970 ;
        RECT 89.990 374.640 95.350 374.920 ;
        RECT 89.990 374.590 90.370 374.640 ;
        RECT 94.970 374.590 95.350 374.640 ;
        RECT 122.440 374.920 122.820 374.970 ;
        RECT 127.420 374.920 127.800 374.970 ;
        RECT 122.440 374.640 127.800 374.920 ;
        RECT 122.440 374.590 122.820 374.640 ;
        RECT 127.420 374.590 127.800 374.640 ;
        RECT 154.890 374.920 155.270 374.970 ;
        RECT 159.870 374.920 160.250 374.970 ;
        RECT 154.890 374.640 160.250 374.920 ;
        RECT 162.315 374.765 162.695 375.145 ;
        RECT 164.355 374.765 164.735 375.145 ;
        RECT 166.140 374.765 166.520 375.145 ;
        RECT 154.890 374.590 155.270 374.640 ;
        RECT 159.870 374.590 160.250 374.640 ;
        RECT 25.200 373.265 25.580 373.645 ;
        RECT 29.120 373.265 29.500 373.645 ;
        RECT 31.920 373.310 34.160 373.690 ;
        RECT 64.370 373.310 66.610 373.690 ;
        RECT 96.820 373.310 99.060 373.690 ;
        RECT 129.270 373.310 131.510 373.690 ;
        RECT 58.820 373.080 59.200 373.130 ;
        RECT 62.520 373.080 62.900 373.130 ;
        RECT 58.820 372.800 62.900 373.080 ;
        RECT 58.820 372.750 59.200 372.800 ;
        RECT 62.520 372.750 62.900 372.800 ;
        RECT 91.270 373.080 91.650 373.130 ;
        RECT 94.970 373.080 95.350 373.130 ;
        RECT 91.270 372.800 95.350 373.080 ;
        RECT 91.270 372.750 91.650 372.800 ;
        RECT 94.970 372.750 95.350 372.800 ;
        RECT 123.720 373.080 124.100 373.130 ;
        RECT 127.420 373.080 127.800 373.130 ;
        RECT 123.720 372.800 127.800 373.080 ;
        RECT 123.720 372.750 124.100 372.800 ;
        RECT 127.420 372.750 127.800 372.800 ;
        RECT 156.170 373.080 156.550 373.130 ;
        RECT 159.870 373.080 160.250 373.130 ;
        RECT 156.170 372.800 160.250 373.080 ;
        RECT 156.170 372.750 156.550 372.800 ;
        RECT 159.870 372.750 160.250 372.800 ;
        RECT 31.925 371.425 34.165 371.805 ;
        RECT 64.375 371.425 66.615 371.805 ;
        RECT 96.825 371.425 99.065 371.805 ;
        RECT 129.275 371.425 131.515 371.805 ;
        RECT 162.315 371.765 162.695 372.145 ;
        RECT 164.355 371.765 164.735 372.145 ;
        RECT 166.140 371.765 166.520 372.145 ;
        RECT 31.920 370.665 34.160 371.045 ;
        RECT 64.370 370.665 66.610 371.045 ;
        RECT 96.820 370.665 99.060 371.045 ;
        RECT 129.270 370.665 131.510 371.045 ;
        RECT 25.200 370.265 25.580 370.645 ;
        RECT 29.120 370.265 29.500 370.645 ;
        RECT 60.100 370.435 60.480 370.485 ;
        RECT 62.520 370.435 62.900 370.485 ;
        RECT 60.100 370.155 62.900 370.435 ;
        RECT 60.100 370.105 60.480 370.155 ;
        RECT 62.520 370.105 62.900 370.155 ;
        RECT 92.550 370.435 92.930 370.485 ;
        RECT 94.970 370.435 95.350 370.485 ;
        RECT 92.550 370.155 95.350 370.435 ;
        RECT 92.550 370.105 92.930 370.155 ;
        RECT 94.970 370.105 95.350 370.155 ;
        RECT 125.000 370.435 125.380 370.485 ;
        RECT 127.420 370.435 127.800 370.485 ;
        RECT 125.000 370.155 127.800 370.435 ;
        RECT 125.000 370.105 125.380 370.155 ;
        RECT 127.420 370.105 127.800 370.155 ;
        RECT 157.450 370.435 157.830 370.485 ;
        RECT 159.870 370.435 160.250 370.485 ;
        RECT 157.450 370.155 160.250 370.435 ;
        RECT 157.450 370.105 157.830 370.155 ;
        RECT 159.870 370.105 160.250 370.155 ;
        RECT 31.920 368.825 34.160 369.205 ;
        RECT 64.370 368.825 66.610 369.205 ;
        RECT 96.820 368.825 99.060 369.205 ;
        RECT 129.270 368.825 131.510 369.205 ;
        RECT 162.315 368.765 162.695 369.145 ;
        RECT 164.355 368.765 164.735 369.145 ;
        RECT 166.140 368.765 166.520 369.145 ;
        RECT 61.380 368.595 61.760 368.645 ;
        RECT 62.520 368.595 62.900 368.645 ;
        RECT 61.380 368.315 62.900 368.595 ;
        RECT 61.380 368.265 61.760 368.315 ;
        RECT 62.520 368.265 62.900 368.315 ;
        RECT 93.830 368.595 94.210 368.645 ;
        RECT 94.970 368.595 95.350 368.645 ;
        RECT 93.830 368.315 95.350 368.595 ;
        RECT 93.830 368.265 94.210 368.315 ;
        RECT 94.970 368.265 95.350 368.315 ;
        RECT 126.280 368.595 126.660 368.645 ;
        RECT 127.420 368.595 127.800 368.645 ;
        RECT 126.280 368.315 127.800 368.595 ;
        RECT 126.280 368.265 126.660 368.315 ;
        RECT 127.420 368.265 127.800 368.315 ;
        RECT 158.730 368.595 159.110 368.645 ;
        RECT 159.870 368.595 160.250 368.645 ;
        RECT 158.730 368.315 160.250 368.595 ;
        RECT 158.730 368.265 159.110 368.315 ;
        RECT 159.870 368.265 160.250 368.315 ;
        RECT 25.200 367.265 25.580 367.645 ;
        RECT 29.120 367.265 29.500 367.645 ;
        RECT 31.920 366.985 34.160 367.365 ;
        RECT 64.370 366.985 66.610 367.365 ;
        RECT 96.820 366.985 99.060 367.365 ;
        RECT 129.270 366.985 131.510 367.365 ;
        RECT 62.520 366.425 63.040 366.805 ;
        RECT 94.970 366.425 95.490 366.805 ;
        RECT 127.420 366.425 127.940 366.805 ;
        RECT 159.870 366.425 160.390 366.805 ;
        RECT 162.315 365.765 162.695 366.145 ;
        RECT 164.355 365.765 164.735 366.145 ;
        RECT 166.140 365.765 166.520 366.145 ;
        RECT 25.200 364.265 25.580 364.645 ;
        RECT 29.120 364.265 29.500 364.645 ;
        RECT 25.200 361.265 25.580 361.645 ;
        RECT 162.315 359.765 162.695 360.145 ;
        RECT 164.355 359.765 164.735 360.145 ;
        RECT 166.140 359.765 166.520 360.145 ;
        RECT 25.200 358.265 25.580 358.645 ;
        RECT 29.120 358.265 29.500 358.645 ;
        RECT 62.020 357.860 62.900 358.240 ;
        RECT 94.470 357.860 95.350 358.240 ;
        RECT 126.920 357.860 127.800 358.240 ;
        RECT 159.370 357.860 160.250 358.240 ;
        RECT 31.920 357.300 34.160 357.680 ;
        RECT 64.370 357.300 66.610 357.680 ;
        RECT 96.820 357.300 99.060 357.680 ;
        RECT 129.270 357.300 131.510 357.680 ;
        RECT 162.315 356.765 162.695 357.145 ;
        RECT 164.355 356.765 164.735 357.145 ;
        RECT 166.140 356.765 166.520 357.145 ;
        RECT 60.740 356.350 61.120 356.400 ;
        RECT 62.520 356.350 62.900 356.400 ;
        RECT 60.740 356.070 62.900 356.350 ;
        RECT 60.740 356.020 61.120 356.070 ;
        RECT 62.520 356.020 62.900 356.070 ;
        RECT 93.190 356.350 93.570 356.400 ;
        RECT 94.970 356.350 95.350 356.400 ;
        RECT 93.190 356.070 95.350 356.350 ;
        RECT 93.190 356.020 93.570 356.070 ;
        RECT 94.970 356.020 95.350 356.070 ;
        RECT 125.640 356.350 126.020 356.400 ;
        RECT 127.420 356.350 127.800 356.400 ;
        RECT 125.640 356.070 127.800 356.350 ;
        RECT 125.640 356.020 126.020 356.070 ;
        RECT 127.420 356.020 127.800 356.070 ;
        RECT 158.090 356.350 158.470 356.400 ;
        RECT 159.870 356.350 160.250 356.400 ;
        RECT 158.090 356.070 160.250 356.350 ;
        RECT 158.090 356.020 158.470 356.070 ;
        RECT 159.870 356.020 160.250 356.070 ;
        RECT 25.200 355.265 25.580 355.645 ;
        RECT 29.120 355.265 29.500 355.645 ;
        RECT 31.920 355.460 34.160 355.840 ;
        RECT 64.370 355.460 66.610 355.840 ;
        RECT 96.820 355.460 99.060 355.840 ;
        RECT 129.270 355.460 131.510 355.840 ;
        RECT 59.460 354.505 59.840 354.555 ;
        RECT 62.520 354.505 62.900 354.555 ;
        RECT 59.460 354.225 62.900 354.505 ;
        RECT 59.460 354.175 59.840 354.225 ;
        RECT 62.520 354.175 62.900 354.225 ;
        RECT 91.910 354.505 92.290 354.555 ;
        RECT 94.970 354.505 95.350 354.555 ;
        RECT 91.910 354.225 95.350 354.505 ;
        RECT 91.910 354.175 92.290 354.225 ;
        RECT 94.970 354.175 95.350 354.225 ;
        RECT 124.360 354.505 124.740 354.555 ;
        RECT 127.420 354.505 127.800 354.555 ;
        RECT 124.360 354.225 127.800 354.505 ;
        RECT 124.360 354.175 124.740 354.225 ;
        RECT 127.420 354.175 127.800 354.225 ;
        RECT 156.810 354.505 157.190 354.555 ;
        RECT 159.870 354.505 160.250 354.555 ;
        RECT 156.810 354.225 160.250 354.505 ;
        RECT 156.810 354.175 157.190 354.225 ;
        RECT 159.870 354.175 160.250 354.225 ;
        RECT 31.920 353.615 34.160 353.995 ;
        RECT 64.370 353.615 66.610 353.995 ;
        RECT 96.820 353.615 99.060 353.995 ;
        RECT 129.270 353.615 131.510 353.995 ;
        RECT 162.315 353.765 162.695 354.145 ;
        RECT 164.355 353.765 164.735 354.145 ;
        RECT 166.140 353.765 166.520 354.145 ;
        RECT 31.925 352.855 34.165 353.235 ;
        RECT 64.375 352.855 66.615 353.235 ;
        RECT 96.825 352.855 99.065 353.235 ;
        RECT 129.275 352.855 131.515 353.235 ;
        RECT 25.200 352.265 25.580 352.645 ;
        RECT 29.120 352.265 29.500 352.645 ;
        RECT 58.180 351.865 58.560 351.915 ;
        RECT 62.520 351.865 62.900 351.915 ;
        RECT 58.180 351.585 62.900 351.865 ;
        RECT 58.180 351.535 58.560 351.585 ;
        RECT 62.520 351.535 62.900 351.585 ;
        RECT 90.630 351.865 91.010 351.915 ;
        RECT 94.970 351.865 95.350 351.915 ;
        RECT 90.630 351.585 95.350 351.865 ;
        RECT 90.630 351.535 91.010 351.585 ;
        RECT 94.970 351.535 95.350 351.585 ;
        RECT 123.080 351.865 123.460 351.915 ;
        RECT 127.420 351.865 127.800 351.915 ;
        RECT 123.080 351.585 127.800 351.865 ;
        RECT 123.080 351.535 123.460 351.585 ;
        RECT 127.420 351.535 127.800 351.585 ;
        RECT 155.530 351.865 155.910 351.915 ;
        RECT 159.870 351.865 160.250 351.915 ;
        RECT 155.530 351.585 160.250 351.865 ;
        RECT 155.530 351.535 155.910 351.585 ;
        RECT 159.870 351.535 160.250 351.585 ;
        RECT 31.920 350.975 34.160 351.355 ;
        RECT 64.370 350.975 66.610 351.355 ;
        RECT 96.820 350.975 99.060 351.355 ;
        RECT 129.270 350.975 131.510 351.355 ;
        RECT 162.315 350.765 162.695 351.145 ;
        RECT 164.355 350.765 164.735 351.145 ;
        RECT 166.140 350.765 166.520 351.145 ;
        RECT 56.900 350.025 57.280 350.075 ;
        RECT 62.520 350.025 62.900 350.075 ;
        RECT 56.900 349.745 62.900 350.025 ;
        RECT 56.900 349.695 57.280 349.745 ;
        RECT 62.520 349.695 62.900 349.745 ;
        RECT 89.350 350.025 89.730 350.075 ;
        RECT 94.970 350.025 95.350 350.075 ;
        RECT 89.350 349.745 95.350 350.025 ;
        RECT 89.350 349.695 89.730 349.745 ;
        RECT 94.970 349.695 95.350 349.745 ;
        RECT 121.800 350.025 122.180 350.075 ;
        RECT 127.420 350.025 127.800 350.075 ;
        RECT 121.800 349.745 127.800 350.025 ;
        RECT 121.800 349.695 122.180 349.745 ;
        RECT 127.420 349.695 127.800 349.745 ;
        RECT 154.250 350.025 154.630 350.075 ;
        RECT 159.870 350.025 160.250 350.075 ;
        RECT 154.250 349.745 160.250 350.025 ;
        RECT 154.250 349.695 154.630 349.745 ;
        RECT 159.870 349.695 160.250 349.745 ;
        RECT 25.200 349.265 25.580 349.645 ;
        RECT 29.120 349.265 29.500 349.645 ;
        RECT 31.920 349.135 34.160 349.515 ;
        RECT 64.370 349.135 66.610 349.515 ;
        RECT 96.820 349.135 99.060 349.515 ;
        RECT 129.270 349.135 131.510 349.515 ;
        RECT 55.620 348.180 56.000 348.230 ;
        RECT 62.520 348.180 62.900 348.230 ;
        RECT 55.620 347.900 62.900 348.180 ;
        RECT 55.620 347.850 56.000 347.900 ;
        RECT 62.520 347.850 62.900 347.900 ;
        RECT 88.070 348.180 88.450 348.230 ;
        RECT 94.970 348.180 95.350 348.230 ;
        RECT 88.070 347.900 95.350 348.180 ;
        RECT 88.070 347.850 88.450 347.900 ;
        RECT 94.970 347.850 95.350 347.900 ;
        RECT 120.520 348.180 120.900 348.230 ;
        RECT 127.420 348.180 127.800 348.230 ;
        RECT 120.520 347.900 127.800 348.180 ;
        RECT 120.520 347.850 120.900 347.900 ;
        RECT 127.420 347.850 127.800 347.900 ;
        RECT 152.970 348.180 153.350 348.230 ;
        RECT 159.870 348.180 160.250 348.230 ;
        RECT 152.970 347.900 160.250 348.180 ;
        RECT 152.970 347.850 153.350 347.900 ;
        RECT 159.870 347.850 160.250 347.900 ;
        RECT 162.315 347.765 162.695 348.145 ;
        RECT 164.355 347.765 164.735 348.145 ;
        RECT 166.140 347.765 166.520 348.145 ;
        RECT 31.920 347.290 34.160 347.670 ;
        RECT 64.370 347.290 66.610 347.670 ;
        RECT 96.820 347.290 99.060 347.670 ;
        RECT 129.270 347.290 131.510 347.670 ;
        RECT 25.200 346.265 25.580 346.645 ;
        RECT 29.120 346.265 29.500 346.645 ;
        RECT 31.925 346.530 34.165 346.910 ;
        RECT 64.375 346.530 66.615 346.910 ;
        RECT 96.825 346.530 99.065 346.910 ;
        RECT 129.275 346.530 131.515 346.910 ;
        RECT 54.340 345.540 54.720 345.590 ;
        RECT 62.520 345.540 62.900 345.590 ;
        RECT 54.340 345.260 62.900 345.540 ;
        RECT 54.340 345.210 54.720 345.260 ;
        RECT 62.520 345.210 62.900 345.260 ;
        RECT 86.790 345.540 87.170 345.590 ;
        RECT 94.970 345.540 95.350 345.590 ;
        RECT 86.790 345.260 95.350 345.540 ;
        RECT 86.790 345.210 87.170 345.260 ;
        RECT 94.970 345.210 95.350 345.260 ;
        RECT 119.240 345.540 119.620 345.590 ;
        RECT 127.420 345.540 127.800 345.590 ;
        RECT 119.240 345.260 127.800 345.540 ;
        RECT 119.240 345.210 119.620 345.260 ;
        RECT 127.420 345.210 127.800 345.260 ;
        RECT 151.690 345.540 152.070 345.590 ;
        RECT 159.870 345.540 160.250 345.590 ;
        RECT 151.690 345.260 160.250 345.540 ;
        RECT 151.690 345.210 152.070 345.260 ;
        RECT 159.870 345.210 160.250 345.260 ;
        RECT 31.920 344.650 34.160 345.030 ;
        RECT 64.370 344.650 66.610 345.030 ;
        RECT 96.820 344.650 99.060 345.030 ;
        RECT 129.270 344.650 131.510 345.030 ;
        RECT 162.315 344.765 162.695 345.145 ;
        RECT 164.355 344.765 164.735 345.145 ;
        RECT 166.140 344.765 166.520 345.145 ;
        RECT 53.060 343.700 53.440 343.750 ;
        RECT 62.520 343.700 62.900 343.750 ;
        RECT 25.200 343.265 25.580 343.645 ;
        RECT 29.120 343.265 29.500 343.645 ;
        RECT 53.060 343.420 62.900 343.700 ;
        RECT 53.060 343.370 53.440 343.420 ;
        RECT 62.520 343.370 62.900 343.420 ;
        RECT 85.510 343.700 85.890 343.750 ;
        RECT 94.970 343.700 95.350 343.750 ;
        RECT 85.510 343.420 95.350 343.700 ;
        RECT 85.510 343.370 85.890 343.420 ;
        RECT 94.970 343.370 95.350 343.420 ;
        RECT 117.960 343.700 118.340 343.750 ;
        RECT 127.420 343.700 127.800 343.750 ;
        RECT 117.960 343.420 127.800 343.700 ;
        RECT 117.960 343.370 118.340 343.420 ;
        RECT 127.420 343.370 127.800 343.420 ;
        RECT 150.410 343.700 150.790 343.750 ;
        RECT 159.870 343.700 160.250 343.750 ;
        RECT 150.410 343.420 160.250 343.700 ;
        RECT 150.410 343.370 150.790 343.420 ;
        RECT 159.870 343.370 160.250 343.420 ;
        RECT 31.920 342.810 34.160 343.190 ;
        RECT 64.370 342.810 66.610 343.190 ;
        RECT 96.820 342.810 99.060 343.190 ;
        RECT 129.270 342.810 131.510 343.190 ;
        RECT 31.920 342.090 34.160 342.470 ;
        RECT 64.370 342.090 66.610 342.470 ;
        RECT 96.820 342.090 99.060 342.470 ;
        RECT 129.270 342.090 131.510 342.470 ;
        RECT 53.700 341.860 54.080 341.910 ;
        RECT 62.520 341.860 62.900 341.910 ;
        RECT 53.700 341.580 62.900 341.860 ;
        RECT 53.700 341.530 54.080 341.580 ;
        RECT 62.520 341.530 62.900 341.580 ;
        RECT 86.150 341.860 86.530 341.910 ;
        RECT 94.970 341.860 95.350 341.910 ;
        RECT 86.150 341.580 95.350 341.860 ;
        RECT 86.150 341.530 86.530 341.580 ;
        RECT 94.970 341.530 95.350 341.580 ;
        RECT 118.600 341.860 118.980 341.910 ;
        RECT 127.420 341.860 127.800 341.910 ;
        RECT 118.600 341.580 127.800 341.860 ;
        RECT 118.600 341.530 118.980 341.580 ;
        RECT 127.420 341.530 127.800 341.580 ;
        RECT 151.050 341.860 151.430 341.910 ;
        RECT 159.870 341.860 160.250 341.910 ;
        RECT 151.050 341.580 160.250 341.860 ;
        RECT 151.050 341.530 151.430 341.580 ;
        RECT 159.870 341.530 160.250 341.580 ;
        RECT 25.200 339.880 25.580 340.260 ;
        RECT 29.120 339.880 29.500 340.260 ;
        RECT 31.920 340.250 34.160 340.630 ;
        RECT 64.370 340.250 66.610 340.630 ;
        RECT 96.820 340.250 99.060 340.630 ;
        RECT 129.270 340.250 131.510 340.630 ;
        RECT 54.980 340.020 55.360 340.070 ;
        RECT 62.520 340.020 62.900 340.070 ;
        RECT 54.980 339.740 62.900 340.020 ;
        RECT 54.980 339.690 55.360 339.740 ;
        RECT 62.520 339.690 62.900 339.740 ;
        RECT 87.430 340.020 87.810 340.070 ;
        RECT 94.970 340.020 95.350 340.070 ;
        RECT 87.430 339.740 95.350 340.020 ;
        RECT 87.430 339.690 87.810 339.740 ;
        RECT 94.970 339.690 95.350 339.740 ;
        RECT 119.880 340.020 120.260 340.070 ;
        RECT 127.420 340.020 127.800 340.070 ;
        RECT 119.880 339.740 127.800 340.020 ;
        RECT 119.880 339.690 120.260 339.740 ;
        RECT 127.420 339.690 127.800 339.740 ;
        RECT 152.330 340.020 152.710 340.070 ;
        RECT 159.870 340.020 160.250 340.070 ;
        RECT 152.330 339.740 160.250 340.020 ;
        RECT 152.330 339.690 152.710 339.740 ;
        RECT 159.870 339.690 160.250 339.740 ;
        RECT 31.925 338.365 34.165 338.745 ;
        RECT 64.375 338.365 66.615 338.745 ;
        RECT 96.825 338.365 99.065 338.745 ;
        RECT 129.275 338.365 131.515 338.745 ;
        RECT 162.315 338.380 162.695 338.760 ;
        RECT 164.355 338.380 164.735 338.760 ;
        RECT 166.140 338.380 166.520 338.760 ;
        RECT 31.920 337.605 34.160 337.985 ;
        RECT 64.370 337.605 66.610 337.985 ;
        RECT 96.820 337.605 99.060 337.985 ;
        RECT 129.270 337.605 131.510 337.985 ;
        RECT 56.260 337.375 56.640 337.425 ;
        RECT 62.520 337.375 62.900 337.425 ;
        RECT 25.200 336.880 25.580 337.260 ;
        RECT 29.120 336.880 29.500 337.260 ;
        RECT 56.260 337.095 62.900 337.375 ;
        RECT 56.260 337.045 56.640 337.095 ;
        RECT 62.520 337.045 62.900 337.095 ;
        RECT 88.710 337.375 89.090 337.425 ;
        RECT 94.970 337.375 95.350 337.425 ;
        RECT 88.710 337.095 95.350 337.375 ;
        RECT 88.710 337.045 89.090 337.095 ;
        RECT 94.970 337.045 95.350 337.095 ;
        RECT 121.160 337.375 121.540 337.425 ;
        RECT 127.420 337.375 127.800 337.425 ;
        RECT 121.160 337.095 127.800 337.375 ;
        RECT 121.160 337.045 121.540 337.095 ;
        RECT 127.420 337.045 127.800 337.095 ;
        RECT 153.610 337.375 153.990 337.425 ;
        RECT 159.870 337.375 160.250 337.425 ;
        RECT 153.610 337.095 160.250 337.375 ;
        RECT 153.610 337.045 153.990 337.095 ;
        RECT 159.870 337.045 160.250 337.095 ;
        RECT 31.920 335.765 34.160 336.145 ;
        RECT 64.370 335.765 66.610 336.145 ;
        RECT 96.820 335.765 99.060 336.145 ;
        RECT 129.270 335.765 131.510 336.145 ;
        RECT 57.540 335.535 57.920 335.585 ;
        RECT 62.520 335.535 62.900 335.585 ;
        RECT 57.540 335.255 62.900 335.535 ;
        RECT 57.540 335.205 57.920 335.255 ;
        RECT 62.520 335.205 62.900 335.255 ;
        RECT 89.990 335.535 90.370 335.585 ;
        RECT 94.970 335.535 95.350 335.585 ;
        RECT 89.990 335.255 95.350 335.535 ;
        RECT 89.990 335.205 90.370 335.255 ;
        RECT 94.970 335.205 95.350 335.255 ;
        RECT 122.440 335.535 122.820 335.585 ;
        RECT 127.420 335.535 127.800 335.585 ;
        RECT 122.440 335.255 127.800 335.535 ;
        RECT 122.440 335.205 122.820 335.255 ;
        RECT 127.420 335.205 127.800 335.255 ;
        RECT 154.890 335.535 155.270 335.585 ;
        RECT 159.870 335.535 160.250 335.585 ;
        RECT 154.890 335.255 160.250 335.535 ;
        RECT 162.315 335.380 162.695 335.760 ;
        RECT 164.355 335.380 164.735 335.760 ;
        RECT 166.140 335.380 166.520 335.760 ;
        RECT 154.890 335.205 155.270 335.255 ;
        RECT 159.870 335.205 160.250 335.255 ;
        RECT 25.200 333.880 25.580 334.260 ;
        RECT 29.120 333.880 29.500 334.260 ;
        RECT 31.920 333.925 34.160 334.305 ;
        RECT 64.370 333.925 66.610 334.305 ;
        RECT 96.820 333.925 99.060 334.305 ;
        RECT 129.270 333.925 131.510 334.305 ;
        RECT 58.820 333.695 59.200 333.745 ;
        RECT 62.520 333.695 62.900 333.745 ;
        RECT 58.820 333.415 62.900 333.695 ;
        RECT 58.820 333.365 59.200 333.415 ;
        RECT 62.520 333.365 62.900 333.415 ;
        RECT 91.270 333.695 91.650 333.745 ;
        RECT 94.970 333.695 95.350 333.745 ;
        RECT 91.270 333.415 95.350 333.695 ;
        RECT 91.270 333.365 91.650 333.415 ;
        RECT 94.970 333.365 95.350 333.415 ;
        RECT 123.720 333.695 124.100 333.745 ;
        RECT 127.420 333.695 127.800 333.745 ;
        RECT 123.720 333.415 127.800 333.695 ;
        RECT 123.720 333.365 124.100 333.415 ;
        RECT 127.420 333.365 127.800 333.415 ;
        RECT 156.170 333.695 156.550 333.745 ;
        RECT 159.870 333.695 160.250 333.745 ;
        RECT 156.170 333.415 160.250 333.695 ;
        RECT 156.170 333.365 156.550 333.415 ;
        RECT 159.870 333.365 160.250 333.415 ;
        RECT 31.925 332.040 34.165 332.420 ;
        RECT 64.375 332.040 66.615 332.420 ;
        RECT 96.825 332.040 99.065 332.420 ;
        RECT 129.275 332.040 131.515 332.420 ;
        RECT 162.315 332.380 162.695 332.760 ;
        RECT 164.355 332.380 164.735 332.760 ;
        RECT 166.140 332.380 166.520 332.760 ;
        RECT 31.920 331.280 34.160 331.660 ;
        RECT 64.370 331.280 66.610 331.660 ;
        RECT 96.820 331.280 99.060 331.660 ;
        RECT 129.270 331.280 131.510 331.660 ;
        RECT 25.200 330.880 25.580 331.260 ;
        RECT 29.120 330.880 29.500 331.260 ;
        RECT 60.100 331.050 60.480 331.100 ;
        RECT 62.520 331.050 62.900 331.100 ;
        RECT 60.100 330.770 62.900 331.050 ;
        RECT 60.100 330.720 60.480 330.770 ;
        RECT 62.520 330.720 62.900 330.770 ;
        RECT 92.550 331.050 92.930 331.100 ;
        RECT 94.970 331.050 95.350 331.100 ;
        RECT 92.550 330.770 95.350 331.050 ;
        RECT 92.550 330.720 92.930 330.770 ;
        RECT 94.970 330.720 95.350 330.770 ;
        RECT 125.000 331.050 125.380 331.100 ;
        RECT 127.420 331.050 127.800 331.100 ;
        RECT 125.000 330.770 127.800 331.050 ;
        RECT 125.000 330.720 125.380 330.770 ;
        RECT 127.420 330.720 127.800 330.770 ;
        RECT 157.450 331.050 157.830 331.100 ;
        RECT 159.870 331.050 160.250 331.100 ;
        RECT 157.450 330.770 160.250 331.050 ;
        RECT 157.450 330.720 157.830 330.770 ;
        RECT 159.870 330.720 160.250 330.770 ;
        RECT 31.920 329.440 34.160 329.820 ;
        RECT 64.370 329.440 66.610 329.820 ;
        RECT 96.820 329.440 99.060 329.820 ;
        RECT 129.270 329.440 131.510 329.820 ;
        RECT 162.315 329.380 162.695 329.760 ;
        RECT 164.355 329.380 164.735 329.760 ;
        RECT 166.140 329.380 166.520 329.760 ;
        RECT 61.380 329.210 61.760 329.260 ;
        RECT 62.520 329.210 62.900 329.260 ;
        RECT 61.380 328.930 62.900 329.210 ;
        RECT 61.380 328.880 61.760 328.930 ;
        RECT 62.520 328.880 62.900 328.930 ;
        RECT 93.830 329.210 94.210 329.260 ;
        RECT 94.970 329.210 95.350 329.260 ;
        RECT 93.830 328.930 95.350 329.210 ;
        RECT 93.830 328.880 94.210 328.930 ;
        RECT 94.970 328.880 95.350 328.930 ;
        RECT 126.280 329.210 126.660 329.260 ;
        RECT 127.420 329.210 127.800 329.260 ;
        RECT 126.280 328.930 127.800 329.210 ;
        RECT 126.280 328.880 126.660 328.930 ;
        RECT 127.420 328.880 127.800 328.930 ;
        RECT 158.730 329.210 159.110 329.260 ;
        RECT 159.870 329.210 160.250 329.260 ;
        RECT 158.730 328.930 160.250 329.210 ;
        RECT 158.730 328.880 159.110 328.930 ;
        RECT 159.870 328.880 160.250 328.930 ;
        RECT 25.200 327.880 25.580 328.260 ;
        RECT 29.120 327.880 29.500 328.260 ;
        RECT 31.920 327.600 34.160 327.980 ;
        RECT 64.370 327.600 66.610 327.980 ;
        RECT 96.820 327.600 99.060 327.980 ;
        RECT 129.270 327.600 131.510 327.980 ;
        RECT 62.520 327.040 63.040 327.420 ;
        RECT 94.970 327.040 95.490 327.420 ;
        RECT 127.420 327.040 127.940 327.420 ;
        RECT 159.870 327.040 160.390 327.420 ;
        RECT 162.315 326.380 162.695 326.760 ;
        RECT 164.355 326.380 164.735 326.760 ;
        RECT 166.140 326.380 166.520 326.760 ;
        RECT 25.200 324.880 25.580 325.260 ;
        RECT 29.120 324.880 29.500 325.260 ;
        RECT 25.200 321.880 25.580 322.260 ;
        RECT 162.315 320.380 162.695 320.760 ;
        RECT 164.355 320.380 164.735 320.760 ;
        RECT 166.140 320.380 166.520 320.760 ;
        RECT 25.200 318.880 25.580 319.260 ;
        RECT 29.120 318.880 29.500 319.260 ;
        RECT 62.020 318.475 62.900 318.855 ;
        RECT 94.470 318.475 95.350 318.855 ;
        RECT 126.920 318.475 127.800 318.855 ;
        RECT 159.370 318.475 160.250 318.855 ;
        RECT 31.920 317.915 34.160 318.295 ;
        RECT 64.370 317.915 66.610 318.295 ;
        RECT 96.820 317.915 99.060 318.295 ;
        RECT 129.270 317.915 131.510 318.295 ;
        RECT 162.315 317.380 162.695 317.760 ;
        RECT 164.355 317.380 164.735 317.760 ;
        RECT 166.140 317.380 166.520 317.760 ;
        RECT 60.740 316.965 61.120 317.015 ;
        RECT 62.520 316.965 62.900 317.015 ;
        RECT 60.740 316.685 62.900 316.965 ;
        RECT 60.740 316.635 61.120 316.685 ;
        RECT 62.520 316.635 62.900 316.685 ;
        RECT 93.190 316.965 93.570 317.015 ;
        RECT 94.970 316.965 95.350 317.015 ;
        RECT 93.190 316.685 95.350 316.965 ;
        RECT 93.190 316.635 93.570 316.685 ;
        RECT 94.970 316.635 95.350 316.685 ;
        RECT 125.640 316.965 126.020 317.015 ;
        RECT 127.420 316.965 127.800 317.015 ;
        RECT 125.640 316.685 127.800 316.965 ;
        RECT 125.640 316.635 126.020 316.685 ;
        RECT 127.420 316.635 127.800 316.685 ;
        RECT 158.090 316.965 158.470 317.015 ;
        RECT 159.870 316.965 160.250 317.015 ;
        RECT 158.090 316.685 160.250 316.965 ;
        RECT 158.090 316.635 158.470 316.685 ;
        RECT 159.870 316.635 160.250 316.685 ;
        RECT 25.200 315.880 25.580 316.260 ;
        RECT 29.120 315.880 29.500 316.260 ;
        RECT 31.920 316.075 34.160 316.455 ;
        RECT 64.370 316.075 66.610 316.455 ;
        RECT 96.820 316.075 99.060 316.455 ;
        RECT 129.270 316.075 131.510 316.455 ;
        RECT 59.460 315.120 59.840 315.170 ;
        RECT 62.520 315.120 62.900 315.170 ;
        RECT 59.460 314.840 62.900 315.120 ;
        RECT 59.460 314.790 59.840 314.840 ;
        RECT 62.520 314.790 62.900 314.840 ;
        RECT 91.910 315.120 92.290 315.170 ;
        RECT 94.970 315.120 95.350 315.170 ;
        RECT 91.910 314.840 95.350 315.120 ;
        RECT 91.910 314.790 92.290 314.840 ;
        RECT 94.970 314.790 95.350 314.840 ;
        RECT 124.360 315.120 124.740 315.170 ;
        RECT 127.420 315.120 127.800 315.170 ;
        RECT 124.360 314.840 127.800 315.120 ;
        RECT 124.360 314.790 124.740 314.840 ;
        RECT 127.420 314.790 127.800 314.840 ;
        RECT 156.810 315.120 157.190 315.170 ;
        RECT 159.870 315.120 160.250 315.170 ;
        RECT 156.810 314.840 160.250 315.120 ;
        RECT 156.810 314.790 157.190 314.840 ;
        RECT 159.870 314.790 160.250 314.840 ;
        RECT 31.920 314.230 34.160 314.610 ;
        RECT 64.370 314.230 66.610 314.610 ;
        RECT 96.820 314.230 99.060 314.610 ;
        RECT 129.270 314.230 131.510 314.610 ;
        RECT 162.315 314.380 162.695 314.760 ;
        RECT 164.355 314.380 164.735 314.760 ;
        RECT 166.140 314.380 166.520 314.760 ;
        RECT 31.925 313.470 34.165 313.850 ;
        RECT 64.375 313.470 66.615 313.850 ;
        RECT 96.825 313.470 99.065 313.850 ;
        RECT 129.275 313.470 131.515 313.850 ;
        RECT 25.200 312.880 25.580 313.260 ;
        RECT 29.120 312.880 29.500 313.260 ;
        RECT 58.180 312.480 58.560 312.530 ;
        RECT 62.520 312.480 62.900 312.530 ;
        RECT 58.180 312.200 62.900 312.480 ;
        RECT 58.180 312.150 58.560 312.200 ;
        RECT 62.520 312.150 62.900 312.200 ;
        RECT 90.630 312.480 91.010 312.530 ;
        RECT 94.970 312.480 95.350 312.530 ;
        RECT 90.630 312.200 95.350 312.480 ;
        RECT 90.630 312.150 91.010 312.200 ;
        RECT 94.970 312.150 95.350 312.200 ;
        RECT 123.080 312.480 123.460 312.530 ;
        RECT 127.420 312.480 127.800 312.530 ;
        RECT 123.080 312.200 127.800 312.480 ;
        RECT 123.080 312.150 123.460 312.200 ;
        RECT 127.420 312.150 127.800 312.200 ;
        RECT 155.530 312.480 155.910 312.530 ;
        RECT 159.870 312.480 160.250 312.530 ;
        RECT 155.530 312.200 160.250 312.480 ;
        RECT 155.530 312.150 155.910 312.200 ;
        RECT 159.870 312.150 160.250 312.200 ;
        RECT 31.920 311.590 34.160 311.970 ;
        RECT 64.370 311.590 66.610 311.970 ;
        RECT 96.820 311.590 99.060 311.970 ;
        RECT 129.270 311.590 131.510 311.970 ;
        RECT 162.315 311.380 162.695 311.760 ;
        RECT 164.355 311.380 164.735 311.760 ;
        RECT 166.140 311.380 166.520 311.760 ;
        RECT 56.900 310.640 57.280 310.690 ;
        RECT 62.520 310.640 62.900 310.690 ;
        RECT 56.900 310.360 62.900 310.640 ;
        RECT 56.900 310.310 57.280 310.360 ;
        RECT 62.520 310.310 62.900 310.360 ;
        RECT 89.350 310.640 89.730 310.690 ;
        RECT 94.970 310.640 95.350 310.690 ;
        RECT 89.350 310.360 95.350 310.640 ;
        RECT 89.350 310.310 89.730 310.360 ;
        RECT 94.970 310.310 95.350 310.360 ;
        RECT 121.800 310.640 122.180 310.690 ;
        RECT 127.420 310.640 127.800 310.690 ;
        RECT 121.800 310.360 127.800 310.640 ;
        RECT 121.800 310.310 122.180 310.360 ;
        RECT 127.420 310.310 127.800 310.360 ;
        RECT 154.250 310.640 154.630 310.690 ;
        RECT 159.870 310.640 160.250 310.690 ;
        RECT 154.250 310.360 160.250 310.640 ;
        RECT 154.250 310.310 154.630 310.360 ;
        RECT 159.870 310.310 160.250 310.360 ;
        RECT 25.200 309.880 25.580 310.260 ;
        RECT 29.120 309.880 29.500 310.260 ;
        RECT 31.920 309.750 34.160 310.130 ;
        RECT 64.370 309.750 66.610 310.130 ;
        RECT 96.820 309.750 99.060 310.130 ;
        RECT 129.270 309.750 131.510 310.130 ;
        RECT 55.620 308.795 56.000 308.845 ;
        RECT 62.520 308.795 62.900 308.845 ;
        RECT 55.620 308.515 62.900 308.795 ;
        RECT 55.620 308.465 56.000 308.515 ;
        RECT 62.520 308.465 62.900 308.515 ;
        RECT 88.070 308.795 88.450 308.845 ;
        RECT 94.970 308.795 95.350 308.845 ;
        RECT 88.070 308.515 95.350 308.795 ;
        RECT 88.070 308.465 88.450 308.515 ;
        RECT 94.970 308.465 95.350 308.515 ;
        RECT 120.520 308.795 120.900 308.845 ;
        RECT 127.420 308.795 127.800 308.845 ;
        RECT 120.520 308.515 127.800 308.795 ;
        RECT 120.520 308.465 120.900 308.515 ;
        RECT 127.420 308.465 127.800 308.515 ;
        RECT 152.970 308.795 153.350 308.845 ;
        RECT 159.870 308.795 160.250 308.845 ;
        RECT 152.970 308.515 160.250 308.795 ;
        RECT 152.970 308.465 153.350 308.515 ;
        RECT 159.870 308.465 160.250 308.515 ;
        RECT 162.315 308.380 162.695 308.760 ;
        RECT 164.355 308.380 164.735 308.760 ;
        RECT 166.140 308.380 166.520 308.760 ;
        RECT 31.920 307.905 34.160 308.285 ;
        RECT 64.370 307.905 66.610 308.285 ;
        RECT 96.820 307.905 99.060 308.285 ;
        RECT 129.270 307.905 131.510 308.285 ;
        RECT 25.200 306.880 25.580 307.260 ;
        RECT 29.120 306.880 29.500 307.260 ;
        RECT 31.925 307.145 34.165 307.525 ;
        RECT 64.375 307.145 66.615 307.525 ;
        RECT 96.825 307.145 99.065 307.525 ;
        RECT 129.275 307.145 131.515 307.525 ;
        RECT 54.340 306.155 54.720 306.205 ;
        RECT 62.520 306.155 62.900 306.205 ;
        RECT 54.340 305.875 62.900 306.155 ;
        RECT 54.340 305.825 54.720 305.875 ;
        RECT 62.520 305.825 62.900 305.875 ;
        RECT 86.790 306.155 87.170 306.205 ;
        RECT 94.970 306.155 95.350 306.205 ;
        RECT 86.790 305.875 95.350 306.155 ;
        RECT 86.790 305.825 87.170 305.875 ;
        RECT 94.970 305.825 95.350 305.875 ;
        RECT 119.240 306.155 119.620 306.205 ;
        RECT 127.420 306.155 127.800 306.205 ;
        RECT 119.240 305.875 127.800 306.155 ;
        RECT 119.240 305.825 119.620 305.875 ;
        RECT 127.420 305.825 127.800 305.875 ;
        RECT 151.690 306.155 152.070 306.205 ;
        RECT 159.870 306.155 160.250 306.205 ;
        RECT 151.690 305.875 160.250 306.155 ;
        RECT 151.690 305.825 152.070 305.875 ;
        RECT 159.870 305.825 160.250 305.875 ;
        RECT 31.920 305.265 34.160 305.645 ;
        RECT 64.370 305.265 66.610 305.645 ;
        RECT 96.820 305.265 99.060 305.645 ;
        RECT 129.270 305.265 131.510 305.645 ;
        RECT 162.315 305.380 162.695 305.760 ;
        RECT 164.355 305.380 164.735 305.760 ;
        RECT 166.140 305.380 166.520 305.760 ;
        RECT 53.060 304.315 53.440 304.365 ;
        RECT 62.520 304.315 62.900 304.365 ;
        RECT 25.200 303.880 25.580 304.260 ;
        RECT 29.120 303.880 29.500 304.260 ;
        RECT 53.060 304.035 62.900 304.315 ;
        RECT 53.060 303.985 53.440 304.035 ;
        RECT 62.520 303.985 62.900 304.035 ;
        RECT 85.510 304.315 85.890 304.365 ;
        RECT 94.970 304.315 95.350 304.365 ;
        RECT 85.510 304.035 95.350 304.315 ;
        RECT 85.510 303.985 85.890 304.035 ;
        RECT 94.970 303.985 95.350 304.035 ;
        RECT 117.960 304.315 118.340 304.365 ;
        RECT 127.420 304.315 127.800 304.365 ;
        RECT 117.960 304.035 127.800 304.315 ;
        RECT 117.960 303.985 118.340 304.035 ;
        RECT 127.420 303.985 127.800 304.035 ;
        RECT 150.410 304.315 150.790 304.365 ;
        RECT 159.870 304.315 160.250 304.365 ;
        RECT 150.410 304.035 160.250 304.315 ;
        RECT 150.410 303.985 150.790 304.035 ;
        RECT 159.870 303.985 160.250 304.035 ;
        RECT 31.920 303.425 34.160 303.805 ;
        RECT 64.370 303.425 66.610 303.805 ;
        RECT 96.820 303.425 99.060 303.805 ;
        RECT 129.270 303.425 131.510 303.805 ;
        RECT 31.920 302.705 34.160 303.085 ;
        RECT 64.370 302.705 66.610 303.085 ;
        RECT 96.820 302.705 99.060 303.085 ;
        RECT 129.270 302.705 131.510 303.085 ;
        RECT 53.700 302.475 54.080 302.525 ;
        RECT 62.520 302.475 62.900 302.525 ;
        RECT 53.700 302.195 62.900 302.475 ;
        RECT 53.700 302.145 54.080 302.195 ;
        RECT 62.520 302.145 62.900 302.195 ;
        RECT 86.150 302.475 86.530 302.525 ;
        RECT 94.970 302.475 95.350 302.525 ;
        RECT 86.150 302.195 95.350 302.475 ;
        RECT 86.150 302.145 86.530 302.195 ;
        RECT 94.970 302.145 95.350 302.195 ;
        RECT 118.600 302.475 118.980 302.525 ;
        RECT 127.420 302.475 127.800 302.525 ;
        RECT 118.600 302.195 127.800 302.475 ;
        RECT 118.600 302.145 118.980 302.195 ;
        RECT 127.420 302.145 127.800 302.195 ;
        RECT 151.050 302.475 151.430 302.525 ;
        RECT 159.870 302.475 160.250 302.525 ;
        RECT 151.050 302.195 160.250 302.475 ;
        RECT 151.050 302.145 151.430 302.195 ;
        RECT 159.870 302.145 160.250 302.195 ;
        RECT 25.200 300.495 25.580 300.875 ;
        RECT 29.120 300.495 29.500 300.875 ;
        RECT 31.920 300.865 34.160 301.245 ;
        RECT 64.370 300.865 66.610 301.245 ;
        RECT 96.820 300.865 99.060 301.245 ;
        RECT 129.270 300.865 131.510 301.245 ;
        RECT 54.980 300.635 55.360 300.685 ;
        RECT 62.520 300.635 62.900 300.685 ;
        RECT 54.980 300.355 62.900 300.635 ;
        RECT 54.980 300.305 55.360 300.355 ;
        RECT 62.520 300.305 62.900 300.355 ;
        RECT 87.430 300.635 87.810 300.685 ;
        RECT 94.970 300.635 95.350 300.685 ;
        RECT 87.430 300.355 95.350 300.635 ;
        RECT 87.430 300.305 87.810 300.355 ;
        RECT 94.970 300.305 95.350 300.355 ;
        RECT 119.880 300.635 120.260 300.685 ;
        RECT 127.420 300.635 127.800 300.685 ;
        RECT 119.880 300.355 127.800 300.635 ;
        RECT 119.880 300.305 120.260 300.355 ;
        RECT 127.420 300.305 127.800 300.355 ;
        RECT 152.330 300.635 152.710 300.685 ;
        RECT 159.870 300.635 160.250 300.685 ;
        RECT 152.330 300.355 160.250 300.635 ;
        RECT 152.330 300.305 152.710 300.355 ;
        RECT 159.870 300.305 160.250 300.355 ;
        RECT 31.925 298.980 34.165 299.360 ;
        RECT 64.375 298.980 66.615 299.360 ;
        RECT 96.825 298.980 99.065 299.360 ;
        RECT 129.275 298.980 131.515 299.360 ;
        RECT 162.315 298.995 162.695 299.375 ;
        RECT 164.355 298.995 164.735 299.375 ;
        RECT 166.140 298.995 166.520 299.375 ;
        RECT 31.920 298.220 34.160 298.600 ;
        RECT 64.370 298.220 66.610 298.600 ;
        RECT 96.820 298.220 99.060 298.600 ;
        RECT 129.270 298.220 131.510 298.600 ;
        RECT 56.260 297.990 56.640 298.040 ;
        RECT 62.520 297.990 62.900 298.040 ;
        RECT 25.200 297.495 25.580 297.875 ;
        RECT 29.120 297.495 29.500 297.875 ;
        RECT 56.260 297.710 62.900 297.990 ;
        RECT 56.260 297.660 56.640 297.710 ;
        RECT 62.520 297.660 62.900 297.710 ;
        RECT 88.710 297.990 89.090 298.040 ;
        RECT 94.970 297.990 95.350 298.040 ;
        RECT 88.710 297.710 95.350 297.990 ;
        RECT 88.710 297.660 89.090 297.710 ;
        RECT 94.970 297.660 95.350 297.710 ;
        RECT 121.160 297.990 121.540 298.040 ;
        RECT 127.420 297.990 127.800 298.040 ;
        RECT 121.160 297.710 127.800 297.990 ;
        RECT 121.160 297.660 121.540 297.710 ;
        RECT 127.420 297.660 127.800 297.710 ;
        RECT 153.610 297.990 153.990 298.040 ;
        RECT 159.870 297.990 160.250 298.040 ;
        RECT 153.610 297.710 160.250 297.990 ;
        RECT 153.610 297.660 153.990 297.710 ;
        RECT 159.870 297.660 160.250 297.710 ;
        RECT 31.920 296.380 34.160 296.760 ;
        RECT 64.370 296.380 66.610 296.760 ;
        RECT 96.820 296.380 99.060 296.760 ;
        RECT 129.270 296.380 131.510 296.760 ;
        RECT 57.540 296.150 57.920 296.200 ;
        RECT 62.520 296.150 62.900 296.200 ;
        RECT 57.540 295.870 62.900 296.150 ;
        RECT 57.540 295.820 57.920 295.870 ;
        RECT 62.520 295.820 62.900 295.870 ;
        RECT 89.990 296.150 90.370 296.200 ;
        RECT 94.970 296.150 95.350 296.200 ;
        RECT 89.990 295.870 95.350 296.150 ;
        RECT 89.990 295.820 90.370 295.870 ;
        RECT 94.970 295.820 95.350 295.870 ;
        RECT 122.440 296.150 122.820 296.200 ;
        RECT 127.420 296.150 127.800 296.200 ;
        RECT 122.440 295.870 127.800 296.150 ;
        RECT 122.440 295.820 122.820 295.870 ;
        RECT 127.420 295.820 127.800 295.870 ;
        RECT 154.890 296.150 155.270 296.200 ;
        RECT 159.870 296.150 160.250 296.200 ;
        RECT 154.890 295.870 160.250 296.150 ;
        RECT 162.315 295.995 162.695 296.375 ;
        RECT 164.355 295.995 164.735 296.375 ;
        RECT 166.140 295.995 166.520 296.375 ;
        RECT 154.890 295.820 155.270 295.870 ;
        RECT 159.870 295.820 160.250 295.870 ;
        RECT 25.200 294.495 25.580 294.875 ;
        RECT 29.120 294.495 29.500 294.875 ;
        RECT 31.920 294.540 34.160 294.920 ;
        RECT 64.370 294.540 66.610 294.920 ;
        RECT 96.820 294.540 99.060 294.920 ;
        RECT 129.270 294.540 131.510 294.920 ;
        RECT 58.820 294.310 59.200 294.360 ;
        RECT 62.520 294.310 62.900 294.360 ;
        RECT 58.820 294.030 62.900 294.310 ;
        RECT 58.820 293.980 59.200 294.030 ;
        RECT 62.520 293.980 62.900 294.030 ;
        RECT 91.270 294.310 91.650 294.360 ;
        RECT 94.970 294.310 95.350 294.360 ;
        RECT 91.270 294.030 95.350 294.310 ;
        RECT 91.270 293.980 91.650 294.030 ;
        RECT 94.970 293.980 95.350 294.030 ;
        RECT 123.720 294.310 124.100 294.360 ;
        RECT 127.420 294.310 127.800 294.360 ;
        RECT 123.720 294.030 127.800 294.310 ;
        RECT 123.720 293.980 124.100 294.030 ;
        RECT 127.420 293.980 127.800 294.030 ;
        RECT 156.170 294.310 156.550 294.360 ;
        RECT 159.870 294.310 160.250 294.360 ;
        RECT 156.170 294.030 160.250 294.310 ;
        RECT 156.170 293.980 156.550 294.030 ;
        RECT 159.870 293.980 160.250 294.030 ;
        RECT 31.925 292.655 34.165 293.035 ;
        RECT 64.375 292.655 66.615 293.035 ;
        RECT 96.825 292.655 99.065 293.035 ;
        RECT 129.275 292.655 131.515 293.035 ;
        RECT 162.315 292.995 162.695 293.375 ;
        RECT 164.355 292.995 164.735 293.375 ;
        RECT 166.140 292.995 166.520 293.375 ;
        RECT 31.920 291.895 34.160 292.275 ;
        RECT 64.370 291.895 66.610 292.275 ;
        RECT 96.820 291.895 99.060 292.275 ;
        RECT 129.270 291.895 131.510 292.275 ;
        RECT 25.200 291.495 25.580 291.875 ;
        RECT 29.120 291.495 29.500 291.875 ;
        RECT 60.100 291.665 60.480 291.715 ;
        RECT 62.520 291.665 62.900 291.715 ;
        RECT 60.100 291.385 62.900 291.665 ;
        RECT 60.100 291.335 60.480 291.385 ;
        RECT 62.520 291.335 62.900 291.385 ;
        RECT 92.550 291.665 92.930 291.715 ;
        RECT 94.970 291.665 95.350 291.715 ;
        RECT 92.550 291.385 95.350 291.665 ;
        RECT 92.550 291.335 92.930 291.385 ;
        RECT 94.970 291.335 95.350 291.385 ;
        RECT 125.000 291.665 125.380 291.715 ;
        RECT 127.420 291.665 127.800 291.715 ;
        RECT 125.000 291.385 127.800 291.665 ;
        RECT 125.000 291.335 125.380 291.385 ;
        RECT 127.420 291.335 127.800 291.385 ;
        RECT 157.450 291.665 157.830 291.715 ;
        RECT 159.870 291.665 160.250 291.715 ;
        RECT 157.450 291.385 160.250 291.665 ;
        RECT 157.450 291.335 157.830 291.385 ;
        RECT 159.870 291.335 160.250 291.385 ;
        RECT 31.920 290.055 34.160 290.435 ;
        RECT 64.370 290.055 66.610 290.435 ;
        RECT 96.820 290.055 99.060 290.435 ;
        RECT 129.270 290.055 131.510 290.435 ;
        RECT 162.315 289.995 162.695 290.375 ;
        RECT 164.355 289.995 164.735 290.375 ;
        RECT 166.140 289.995 166.520 290.375 ;
        RECT 61.380 289.825 61.760 289.875 ;
        RECT 62.520 289.825 62.900 289.875 ;
        RECT 61.380 289.545 62.900 289.825 ;
        RECT 61.380 289.495 61.760 289.545 ;
        RECT 62.520 289.495 62.900 289.545 ;
        RECT 93.830 289.825 94.210 289.875 ;
        RECT 94.970 289.825 95.350 289.875 ;
        RECT 93.830 289.545 95.350 289.825 ;
        RECT 93.830 289.495 94.210 289.545 ;
        RECT 94.970 289.495 95.350 289.545 ;
        RECT 126.280 289.825 126.660 289.875 ;
        RECT 127.420 289.825 127.800 289.875 ;
        RECT 126.280 289.545 127.800 289.825 ;
        RECT 126.280 289.495 126.660 289.545 ;
        RECT 127.420 289.495 127.800 289.545 ;
        RECT 158.730 289.825 159.110 289.875 ;
        RECT 159.870 289.825 160.250 289.875 ;
        RECT 158.730 289.545 160.250 289.825 ;
        RECT 158.730 289.495 159.110 289.545 ;
        RECT 159.870 289.495 160.250 289.545 ;
        RECT 25.200 288.495 25.580 288.875 ;
        RECT 29.120 288.495 29.500 288.875 ;
        RECT 31.920 288.215 34.160 288.595 ;
        RECT 64.370 288.215 66.610 288.595 ;
        RECT 96.820 288.215 99.060 288.595 ;
        RECT 129.270 288.215 131.510 288.595 ;
        RECT 62.520 287.655 63.040 288.035 ;
        RECT 94.970 287.655 95.490 288.035 ;
        RECT 127.420 287.655 127.940 288.035 ;
        RECT 159.870 287.655 160.390 288.035 ;
        RECT 162.315 286.995 162.695 287.375 ;
        RECT 164.355 286.995 164.735 287.375 ;
        RECT 166.140 286.995 166.520 287.375 ;
        RECT 25.200 285.495 25.580 285.875 ;
        RECT 29.120 285.495 29.500 285.875 ;
        RECT 25.200 282.495 25.580 282.875 ;
        RECT 162.315 280.995 162.695 281.375 ;
        RECT 164.355 280.995 164.735 281.375 ;
        RECT 166.140 280.995 166.520 281.375 ;
        RECT 25.200 279.495 25.580 279.875 ;
        RECT 29.120 279.495 29.500 279.875 ;
        RECT 62.020 279.090 62.900 279.470 ;
        RECT 94.470 279.090 95.350 279.470 ;
        RECT 126.920 279.090 127.800 279.470 ;
        RECT 159.370 279.090 160.250 279.470 ;
        RECT 31.920 278.530 34.160 278.910 ;
        RECT 64.370 278.530 66.610 278.910 ;
        RECT 96.820 278.530 99.060 278.910 ;
        RECT 129.270 278.530 131.510 278.910 ;
        RECT 162.315 277.995 162.695 278.375 ;
        RECT 164.355 277.995 164.735 278.375 ;
        RECT 166.140 277.995 166.520 278.375 ;
        RECT 60.740 277.580 61.120 277.630 ;
        RECT 62.520 277.580 62.900 277.630 ;
        RECT 60.740 277.300 62.900 277.580 ;
        RECT 60.740 277.250 61.120 277.300 ;
        RECT 62.520 277.250 62.900 277.300 ;
        RECT 93.190 277.580 93.570 277.630 ;
        RECT 94.970 277.580 95.350 277.630 ;
        RECT 93.190 277.300 95.350 277.580 ;
        RECT 93.190 277.250 93.570 277.300 ;
        RECT 94.970 277.250 95.350 277.300 ;
        RECT 125.640 277.580 126.020 277.630 ;
        RECT 127.420 277.580 127.800 277.630 ;
        RECT 125.640 277.300 127.800 277.580 ;
        RECT 125.640 277.250 126.020 277.300 ;
        RECT 127.420 277.250 127.800 277.300 ;
        RECT 158.090 277.580 158.470 277.630 ;
        RECT 159.870 277.580 160.250 277.630 ;
        RECT 158.090 277.300 160.250 277.580 ;
        RECT 158.090 277.250 158.470 277.300 ;
        RECT 159.870 277.250 160.250 277.300 ;
        RECT 25.200 276.495 25.580 276.875 ;
        RECT 29.120 276.495 29.500 276.875 ;
        RECT 31.920 276.690 34.160 277.070 ;
        RECT 64.370 276.690 66.610 277.070 ;
        RECT 96.820 276.690 99.060 277.070 ;
        RECT 129.270 276.690 131.510 277.070 ;
        RECT 59.460 275.735 59.840 275.785 ;
        RECT 62.520 275.735 62.900 275.785 ;
        RECT 59.460 275.455 62.900 275.735 ;
        RECT 59.460 275.405 59.840 275.455 ;
        RECT 62.520 275.405 62.900 275.455 ;
        RECT 91.910 275.735 92.290 275.785 ;
        RECT 94.970 275.735 95.350 275.785 ;
        RECT 91.910 275.455 95.350 275.735 ;
        RECT 91.910 275.405 92.290 275.455 ;
        RECT 94.970 275.405 95.350 275.455 ;
        RECT 124.360 275.735 124.740 275.785 ;
        RECT 127.420 275.735 127.800 275.785 ;
        RECT 124.360 275.455 127.800 275.735 ;
        RECT 124.360 275.405 124.740 275.455 ;
        RECT 127.420 275.405 127.800 275.455 ;
        RECT 156.810 275.735 157.190 275.785 ;
        RECT 159.870 275.735 160.250 275.785 ;
        RECT 156.810 275.455 160.250 275.735 ;
        RECT 156.810 275.405 157.190 275.455 ;
        RECT 159.870 275.405 160.250 275.455 ;
        RECT 31.920 274.845 34.160 275.225 ;
        RECT 64.370 274.845 66.610 275.225 ;
        RECT 96.820 274.845 99.060 275.225 ;
        RECT 129.270 274.845 131.510 275.225 ;
        RECT 162.315 274.995 162.695 275.375 ;
        RECT 164.355 274.995 164.735 275.375 ;
        RECT 166.140 274.995 166.520 275.375 ;
        RECT 31.925 274.085 34.165 274.465 ;
        RECT 64.375 274.085 66.615 274.465 ;
        RECT 96.825 274.085 99.065 274.465 ;
        RECT 129.275 274.085 131.515 274.465 ;
        RECT 25.200 273.495 25.580 273.875 ;
        RECT 29.120 273.495 29.500 273.875 ;
        RECT 58.180 273.095 58.560 273.145 ;
        RECT 62.520 273.095 62.900 273.145 ;
        RECT 58.180 272.815 62.900 273.095 ;
        RECT 58.180 272.765 58.560 272.815 ;
        RECT 62.520 272.765 62.900 272.815 ;
        RECT 90.630 273.095 91.010 273.145 ;
        RECT 94.970 273.095 95.350 273.145 ;
        RECT 90.630 272.815 95.350 273.095 ;
        RECT 90.630 272.765 91.010 272.815 ;
        RECT 94.970 272.765 95.350 272.815 ;
        RECT 123.080 273.095 123.460 273.145 ;
        RECT 127.420 273.095 127.800 273.145 ;
        RECT 123.080 272.815 127.800 273.095 ;
        RECT 123.080 272.765 123.460 272.815 ;
        RECT 127.420 272.765 127.800 272.815 ;
        RECT 155.530 273.095 155.910 273.145 ;
        RECT 159.870 273.095 160.250 273.145 ;
        RECT 155.530 272.815 160.250 273.095 ;
        RECT 155.530 272.765 155.910 272.815 ;
        RECT 159.870 272.765 160.250 272.815 ;
        RECT 31.920 272.205 34.160 272.585 ;
        RECT 64.370 272.205 66.610 272.585 ;
        RECT 96.820 272.205 99.060 272.585 ;
        RECT 129.270 272.205 131.510 272.585 ;
        RECT 162.315 271.995 162.695 272.375 ;
        RECT 164.355 271.995 164.735 272.375 ;
        RECT 166.140 271.995 166.520 272.375 ;
        RECT 56.900 271.255 57.280 271.305 ;
        RECT 62.520 271.255 62.900 271.305 ;
        RECT 56.900 270.975 62.900 271.255 ;
        RECT 56.900 270.925 57.280 270.975 ;
        RECT 62.520 270.925 62.900 270.975 ;
        RECT 89.350 271.255 89.730 271.305 ;
        RECT 94.970 271.255 95.350 271.305 ;
        RECT 89.350 270.975 95.350 271.255 ;
        RECT 89.350 270.925 89.730 270.975 ;
        RECT 94.970 270.925 95.350 270.975 ;
        RECT 121.800 271.255 122.180 271.305 ;
        RECT 127.420 271.255 127.800 271.305 ;
        RECT 121.800 270.975 127.800 271.255 ;
        RECT 121.800 270.925 122.180 270.975 ;
        RECT 127.420 270.925 127.800 270.975 ;
        RECT 154.250 271.255 154.630 271.305 ;
        RECT 159.870 271.255 160.250 271.305 ;
        RECT 154.250 270.975 160.250 271.255 ;
        RECT 154.250 270.925 154.630 270.975 ;
        RECT 159.870 270.925 160.250 270.975 ;
        RECT 25.200 270.495 25.580 270.875 ;
        RECT 29.120 270.495 29.500 270.875 ;
        RECT 31.920 270.365 34.160 270.745 ;
        RECT 64.370 270.365 66.610 270.745 ;
        RECT 96.820 270.365 99.060 270.745 ;
        RECT 129.270 270.365 131.510 270.745 ;
        RECT 55.620 269.410 56.000 269.460 ;
        RECT 62.520 269.410 62.900 269.460 ;
        RECT 55.620 269.130 62.900 269.410 ;
        RECT 55.620 269.080 56.000 269.130 ;
        RECT 62.520 269.080 62.900 269.130 ;
        RECT 88.070 269.410 88.450 269.460 ;
        RECT 94.970 269.410 95.350 269.460 ;
        RECT 88.070 269.130 95.350 269.410 ;
        RECT 88.070 269.080 88.450 269.130 ;
        RECT 94.970 269.080 95.350 269.130 ;
        RECT 120.520 269.410 120.900 269.460 ;
        RECT 127.420 269.410 127.800 269.460 ;
        RECT 120.520 269.130 127.800 269.410 ;
        RECT 120.520 269.080 120.900 269.130 ;
        RECT 127.420 269.080 127.800 269.130 ;
        RECT 152.970 269.410 153.350 269.460 ;
        RECT 159.870 269.410 160.250 269.460 ;
        RECT 152.970 269.130 160.250 269.410 ;
        RECT 152.970 269.080 153.350 269.130 ;
        RECT 159.870 269.080 160.250 269.130 ;
        RECT 162.315 268.995 162.695 269.375 ;
        RECT 164.355 268.995 164.735 269.375 ;
        RECT 166.140 268.995 166.520 269.375 ;
        RECT 31.920 268.520 34.160 268.900 ;
        RECT 64.370 268.520 66.610 268.900 ;
        RECT 96.820 268.520 99.060 268.900 ;
        RECT 129.270 268.520 131.510 268.900 ;
        RECT 25.200 267.495 25.580 267.875 ;
        RECT 29.120 267.495 29.500 267.875 ;
        RECT 31.925 267.760 34.165 268.140 ;
        RECT 64.375 267.760 66.615 268.140 ;
        RECT 96.825 267.760 99.065 268.140 ;
        RECT 129.275 267.760 131.515 268.140 ;
        RECT 54.340 266.770 54.720 266.820 ;
        RECT 62.520 266.770 62.900 266.820 ;
        RECT 54.340 266.490 62.900 266.770 ;
        RECT 54.340 266.440 54.720 266.490 ;
        RECT 62.520 266.440 62.900 266.490 ;
        RECT 86.790 266.770 87.170 266.820 ;
        RECT 94.970 266.770 95.350 266.820 ;
        RECT 86.790 266.490 95.350 266.770 ;
        RECT 86.790 266.440 87.170 266.490 ;
        RECT 94.970 266.440 95.350 266.490 ;
        RECT 119.240 266.770 119.620 266.820 ;
        RECT 127.420 266.770 127.800 266.820 ;
        RECT 119.240 266.490 127.800 266.770 ;
        RECT 119.240 266.440 119.620 266.490 ;
        RECT 127.420 266.440 127.800 266.490 ;
        RECT 151.690 266.770 152.070 266.820 ;
        RECT 159.870 266.770 160.250 266.820 ;
        RECT 151.690 266.490 160.250 266.770 ;
        RECT 151.690 266.440 152.070 266.490 ;
        RECT 159.870 266.440 160.250 266.490 ;
        RECT 31.920 265.880 34.160 266.260 ;
        RECT 64.370 265.880 66.610 266.260 ;
        RECT 96.820 265.880 99.060 266.260 ;
        RECT 129.270 265.880 131.510 266.260 ;
        RECT 162.315 265.995 162.695 266.375 ;
        RECT 164.355 265.995 164.735 266.375 ;
        RECT 166.140 265.995 166.520 266.375 ;
        RECT 53.060 264.930 53.440 264.980 ;
        RECT 62.520 264.930 62.900 264.980 ;
        RECT 25.200 264.495 25.580 264.875 ;
        RECT 29.120 264.495 29.500 264.875 ;
        RECT 53.060 264.650 62.900 264.930 ;
        RECT 53.060 264.600 53.440 264.650 ;
        RECT 62.520 264.600 62.900 264.650 ;
        RECT 85.510 264.930 85.890 264.980 ;
        RECT 94.970 264.930 95.350 264.980 ;
        RECT 85.510 264.650 95.350 264.930 ;
        RECT 85.510 264.600 85.890 264.650 ;
        RECT 94.970 264.600 95.350 264.650 ;
        RECT 117.960 264.930 118.340 264.980 ;
        RECT 127.420 264.930 127.800 264.980 ;
        RECT 117.960 264.650 127.800 264.930 ;
        RECT 117.960 264.600 118.340 264.650 ;
        RECT 127.420 264.600 127.800 264.650 ;
        RECT 150.410 264.930 150.790 264.980 ;
        RECT 159.870 264.930 160.250 264.980 ;
        RECT 150.410 264.650 160.250 264.930 ;
        RECT 150.410 264.600 150.790 264.650 ;
        RECT 159.870 264.600 160.250 264.650 ;
        RECT 31.920 264.040 34.160 264.420 ;
        RECT 64.370 264.040 66.610 264.420 ;
        RECT 96.820 264.040 99.060 264.420 ;
        RECT 129.270 264.040 131.510 264.420 ;
        RECT 31.920 263.320 34.160 263.700 ;
        RECT 64.370 263.320 66.610 263.700 ;
        RECT 96.820 263.320 99.060 263.700 ;
        RECT 129.270 263.320 131.510 263.700 ;
        RECT 53.700 263.090 54.080 263.140 ;
        RECT 62.520 263.090 62.900 263.140 ;
        RECT 53.700 262.810 62.900 263.090 ;
        RECT 53.700 262.760 54.080 262.810 ;
        RECT 62.520 262.760 62.900 262.810 ;
        RECT 86.150 263.090 86.530 263.140 ;
        RECT 94.970 263.090 95.350 263.140 ;
        RECT 86.150 262.810 95.350 263.090 ;
        RECT 86.150 262.760 86.530 262.810 ;
        RECT 94.970 262.760 95.350 262.810 ;
        RECT 118.600 263.090 118.980 263.140 ;
        RECT 127.420 263.090 127.800 263.140 ;
        RECT 118.600 262.810 127.800 263.090 ;
        RECT 118.600 262.760 118.980 262.810 ;
        RECT 127.420 262.760 127.800 262.810 ;
        RECT 151.050 263.090 151.430 263.140 ;
        RECT 159.870 263.090 160.250 263.140 ;
        RECT 151.050 262.810 160.250 263.090 ;
        RECT 151.050 262.760 151.430 262.810 ;
        RECT 159.870 262.760 160.250 262.810 ;
        RECT 25.200 261.110 25.580 261.490 ;
        RECT 29.120 261.110 29.500 261.490 ;
        RECT 31.920 261.480 34.160 261.860 ;
        RECT 64.370 261.480 66.610 261.860 ;
        RECT 96.820 261.480 99.060 261.860 ;
        RECT 129.270 261.480 131.510 261.860 ;
        RECT 54.980 261.250 55.360 261.300 ;
        RECT 62.520 261.250 62.900 261.300 ;
        RECT 54.980 260.970 62.900 261.250 ;
        RECT 54.980 260.920 55.360 260.970 ;
        RECT 62.520 260.920 62.900 260.970 ;
        RECT 87.430 261.250 87.810 261.300 ;
        RECT 94.970 261.250 95.350 261.300 ;
        RECT 87.430 260.970 95.350 261.250 ;
        RECT 87.430 260.920 87.810 260.970 ;
        RECT 94.970 260.920 95.350 260.970 ;
        RECT 119.880 261.250 120.260 261.300 ;
        RECT 127.420 261.250 127.800 261.300 ;
        RECT 119.880 260.970 127.800 261.250 ;
        RECT 119.880 260.920 120.260 260.970 ;
        RECT 127.420 260.920 127.800 260.970 ;
        RECT 152.330 261.250 152.710 261.300 ;
        RECT 159.870 261.250 160.250 261.300 ;
        RECT 152.330 260.970 160.250 261.250 ;
        RECT 152.330 260.920 152.710 260.970 ;
        RECT 159.870 260.920 160.250 260.970 ;
        RECT 31.925 259.595 34.165 259.975 ;
        RECT 64.375 259.595 66.615 259.975 ;
        RECT 96.825 259.595 99.065 259.975 ;
        RECT 129.275 259.595 131.515 259.975 ;
        RECT 162.315 259.610 162.695 259.990 ;
        RECT 164.355 259.610 164.735 259.990 ;
        RECT 166.140 259.610 166.520 259.990 ;
        RECT 31.920 258.835 34.160 259.215 ;
        RECT 64.370 258.835 66.610 259.215 ;
        RECT 96.820 258.835 99.060 259.215 ;
        RECT 129.270 258.835 131.510 259.215 ;
        RECT 56.260 258.605 56.640 258.655 ;
        RECT 62.520 258.605 62.900 258.655 ;
        RECT 25.200 258.110 25.580 258.490 ;
        RECT 29.120 258.110 29.500 258.490 ;
        RECT 56.260 258.325 62.900 258.605 ;
        RECT 56.260 258.275 56.640 258.325 ;
        RECT 62.520 258.275 62.900 258.325 ;
        RECT 88.710 258.605 89.090 258.655 ;
        RECT 94.970 258.605 95.350 258.655 ;
        RECT 88.710 258.325 95.350 258.605 ;
        RECT 88.710 258.275 89.090 258.325 ;
        RECT 94.970 258.275 95.350 258.325 ;
        RECT 121.160 258.605 121.540 258.655 ;
        RECT 127.420 258.605 127.800 258.655 ;
        RECT 121.160 258.325 127.800 258.605 ;
        RECT 121.160 258.275 121.540 258.325 ;
        RECT 127.420 258.275 127.800 258.325 ;
        RECT 153.610 258.605 153.990 258.655 ;
        RECT 159.870 258.605 160.250 258.655 ;
        RECT 153.610 258.325 160.250 258.605 ;
        RECT 153.610 258.275 153.990 258.325 ;
        RECT 159.870 258.275 160.250 258.325 ;
        RECT 31.920 256.995 34.160 257.375 ;
        RECT 64.370 256.995 66.610 257.375 ;
        RECT 96.820 256.995 99.060 257.375 ;
        RECT 129.270 256.995 131.510 257.375 ;
        RECT 57.540 256.765 57.920 256.815 ;
        RECT 62.520 256.765 62.900 256.815 ;
        RECT 57.540 256.485 62.900 256.765 ;
        RECT 57.540 256.435 57.920 256.485 ;
        RECT 62.520 256.435 62.900 256.485 ;
        RECT 89.990 256.765 90.370 256.815 ;
        RECT 94.970 256.765 95.350 256.815 ;
        RECT 89.990 256.485 95.350 256.765 ;
        RECT 89.990 256.435 90.370 256.485 ;
        RECT 94.970 256.435 95.350 256.485 ;
        RECT 122.440 256.765 122.820 256.815 ;
        RECT 127.420 256.765 127.800 256.815 ;
        RECT 122.440 256.485 127.800 256.765 ;
        RECT 122.440 256.435 122.820 256.485 ;
        RECT 127.420 256.435 127.800 256.485 ;
        RECT 154.890 256.765 155.270 256.815 ;
        RECT 159.870 256.765 160.250 256.815 ;
        RECT 154.890 256.485 160.250 256.765 ;
        RECT 162.315 256.610 162.695 256.990 ;
        RECT 164.355 256.610 164.735 256.990 ;
        RECT 166.140 256.610 166.520 256.990 ;
        RECT 154.890 256.435 155.270 256.485 ;
        RECT 159.870 256.435 160.250 256.485 ;
        RECT 25.200 255.110 25.580 255.490 ;
        RECT 29.120 255.110 29.500 255.490 ;
        RECT 31.920 255.155 34.160 255.535 ;
        RECT 64.370 255.155 66.610 255.535 ;
        RECT 96.820 255.155 99.060 255.535 ;
        RECT 129.270 255.155 131.510 255.535 ;
        RECT 58.820 254.925 59.200 254.975 ;
        RECT 62.520 254.925 62.900 254.975 ;
        RECT 58.820 254.645 62.900 254.925 ;
        RECT 58.820 254.595 59.200 254.645 ;
        RECT 62.520 254.595 62.900 254.645 ;
        RECT 91.270 254.925 91.650 254.975 ;
        RECT 94.970 254.925 95.350 254.975 ;
        RECT 91.270 254.645 95.350 254.925 ;
        RECT 91.270 254.595 91.650 254.645 ;
        RECT 94.970 254.595 95.350 254.645 ;
        RECT 123.720 254.925 124.100 254.975 ;
        RECT 127.420 254.925 127.800 254.975 ;
        RECT 123.720 254.645 127.800 254.925 ;
        RECT 123.720 254.595 124.100 254.645 ;
        RECT 127.420 254.595 127.800 254.645 ;
        RECT 156.170 254.925 156.550 254.975 ;
        RECT 159.870 254.925 160.250 254.975 ;
        RECT 156.170 254.645 160.250 254.925 ;
        RECT 156.170 254.595 156.550 254.645 ;
        RECT 159.870 254.595 160.250 254.645 ;
        RECT 31.925 253.270 34.165 253.650 ;
        RECT 64.375 253.270 66.615 253.650 ;
        RECT 96.825 253.270 99.065 253.650 ;
        RECT 129.275 253.270 131.515 253.650 ;
        RECT 162.315 253.610 162.695 253.990 ;
        RECT 164.355 253.610 164.735 253.990 ;
        RECT 166.140 253.610 166.520 253.990 ;
        RECT 31.920 252.510 34.160 252.890 ;
        RECT 64.370 252.510 66.610 252.890 ;
        RECT 96.820 252.510 99.060 252.890 ;
        RECT 129.270 252.510 131.510 252.890 ;
        RECT 25.200 252.110 25.580 252.490 ;
        RECT 29.120 252.110 29.500 252.490 ;
        RECT 60.100 252.280 60.480 252.330 ;
        RECT 62.520 252.280 62.900 252.330 ;
        RECT 60.100 252.000 62.900 252.280 ;
        RECT 60.100 251.950 60.480 252.000 ;
        RECT 62.520 251.950 62.900 252.000 ;
        RECT 92.550 252.280 92.930 252.330 ;
        RECT 94.970 252.280 95.350 252.330 ;
        RECT 92.550 252.000 95.350 252.280 ;
        RECT 92.550 251.950 92.930 252.000 ;
        RECT 94.970 251.950 95.350 252.000 ;
        RECT 125.000 252.280 125.380 252.330 ;
        RECT 127.420 252.280 127.800 252.330 ;
        RECT 125.000 252.000 127.800 252.280 ;
        RECT 125.000 251.950 125.380 252.000 ;
        RECT 127.420 251.950 127.800 252.000 ;
        RECT 157.450 252.280 157.830 252.330 ;
        RECT 159.870 252.280 160.250 252.330 ;
        RECT 157.450 252.000 160.250 252.280 ;
        RECT 157.450 251.950 157.830 252.000 ;
        RECT 159.870 251.950 160.250 252.000 ;
        RECT 31.920 250.670 34.160 251.050 ;
        RECT 64.370 250.670 66.610 251.050 ;
        RECT 96.820 250.670 99.060 251.050 ;
        RECT 129.270 250.670 131.510 251.050 ;
        RECT 162.315 250.610 162.695 250.990 ;
        RECT 164.355 250.610 164.735 250.990 ;
        RECT 166.140 250.610 166.520 250.990 ;
        RECT 61.380 250.440 61.760 250.490 ;
        RECT 62.520 250.440 62.900 250.490 ;
        RECT 61.380 250.160 62.900 250.440 ;
        RECT 61.380 250.110 61.760 250.160 ;
        RECT 62.520 250.110 62.900 250.160 ;
        RECT 93.830 250.440 94.210 250.490 ;
        RECT 94.970 250.440 95.350 250.490 ;
        RECT 93.830 250.160 95.350 250.440 ;
        RECT 93.830 250.110 94.210 250.160 ;
        RECT 94.970 250.110 95.350 250.160 ;
        RECT 126.280 250.440 126.660 250.490 ;
        RECT 127.420 250.440 127.800 250.490 ;
        RECT 126.280 250.160 127.800 250.440 ;
        RECT 126.280 250.110 126.660 250.160 ;
        RECT 127.420 250.110 127.800 250.160 ;
        RECT 158.730 250.440 159.110 250.490 ;
        RECT 159.870 250.440 160.250 250.490 ;
        RECT 158.730 250.160 160.250 250.440 ;
        RECT 158.730 250.110 159.110 250.160 ;
        RECT 159.870 250.110 160.250 250.160 ;
        RECT 25.200 249.110 25.580 249.490 ;
        RECT 29.120 249.110 29.500 249.490 ;
        RECT 31.920 248.830 34.160 249.210 ;
        RECT 64.370 248.830 66.610 249.210 ;
        RECT 96.820 248.830 99.060 249.210 ;
        RECT 129.270 248.830 131.510 249.210 ;
        RECT 62.520 248.270 63.040 248.650 ;
        RECT 94.970 248.270 95.490 248.650 ;
        RECT 127.420 248.270 127.940 248.650 ;
        RECT 159.870 248.270 160.390 248.650 ;
        RECT 162.315 247.610 162.695 247.990 ;
        RECT 164.355 247.610 164.735 247.990 ;
        RECT 166.140 247.610 166.520 247.990 ;
        RECT 25.200 246.110 25.580 246.490 ;
        RECT 29.120 246.110 29.500 246.490 ;
        RECT 25.200 243.110 25.580 243.490 ;
        RECT 162.315 241.610 162.695 241.990 ;
        RECT 164.355 241.610 164.735 241.990 ;
        RECT 166.140 241.610 166.520 241.990 ;
        RECT 25.200 240.110 25.580 240.490 ;
        RECT 29.120 240.110 29.500 240.490 ;
        RECT 62.020 239.705 62.900 240.085 ;
        RECT 94.470 239.705 95.350 240.085 ;
        RECT 126.920 239.705 127.800 240.085 ;
        RECT 159.370 239.705 160.250 240.085 ;
        RECT 31.920 239.145 34.160 239.525 ;
        RECT 64.370 239.145 66.610 239.525 ;
        RECT 96.820 239.145 99.060 239.525 ;
        RECT 129.270 239.145 131.510 239.525 ;
        RECT 162.315 238.610 162.695 238.990 ;
        RECT 164.355 238.610 164.735 238.990 ;
        RECT 166.140 238.610 166.520 238.990 ;
        RECT 60.740 238.195 61.120 238.245 ;
        RECT 62.520 238.195 62.900 238.245 ;
        RECT 60.740 237.915 62.900 238.195 ;
        RECT 60.740 237.865 61.120 237.915 ;
        RECT 62.520 237.865 62.900 237.915 ;
        RECT 93.190 238.195 93.570 238.245 ;
        RECT 94.970 238.195 95.350 238.245 ;
        RECT 93.190 237.915 95.350 238.195 ;
        RECT 93.190 237.865 93.570 237.915 ;
        RECT 94.970 237.865 95.350 237.915 ;
        RECT 125.640 238.195 126.020 238.245 ;
        RECT 127.420 238.195 127.800 238.245 ;
        RECT 125.640 237.915 127.800 238.195 ;
        RECT 125.640 237.865 126.020 237.915 ;
        RECT 127.420 237.865 127.800 237.915 ;
        RECT 158.090 238.195 158.470 238.245 ;
        RECT 159.870 238.195 160.250 238.245 ;
        RECT 158.090 237.915 160.250 238.195 ;
        RECT 158.090 237.865 158.470 237.915 ;
        RECT 159.870 237.865 160.250 237.915 ;
        RECT 25.200 237.110 25.580 237.490 ;
        RECT 29.120 237.110 29.500 237.490 ;
        RECT 31.920 237.305 34.160 237.685 ;
        RECT 64.370 237.305 66.610 237.685 ;
        RECT 96.820 237.305 99.060 237.685 ;
        RECT 129.270 237.305 131.510 237.685 ;
        RECT 59.460 236.350 59.840 236.400 ;
        RECT 62.520 236.350 62.900 236.400 ;
        RECT 59.460 236.070 62.900 236.350 ;
        RECT 59.460 236.020 59.840 236.070 ;
        RECT 62.520 236.020 62.900 236.070 ;
        RECT 91.910 236.350 92.290 236.400 ;
        RECT 94.970 236.350 95.350 236.400 ;
        RECT 91.910 236.070 95.350 236.350 ;
        RECT 91.910 236.020 92.290 236.070 ;
        RECT 94.970 236.020 95.350 236.070 ;
        RECT 124.360 236.350 124.740 236.400 ;
        RECT 127.420 236.350 127.800 236.400 ;
        RECT 124.360 236.070 127.800 236.350 ;
        RECT 124.360 236.020 124.740 236.070 ;
        RECT 127.420 236.020 127.800 236.070 ;
        RECT 156.810 236.350 157.190 236.400 ;
        RECT 159.870 236.350 160.250 236.400 ;
        RECT 156.810 236.070 160.250 236.350 ;
        RECT 156.810 236.020 157.190 236.070 ;
        RECT 159.870 236.020 160.250 236.070 ;
        RECT 31.920 235.460 34.160 235.840 ;
        RECT 64.370 235.460 66.610 235.840 ;
        RECT 96.820 235.460 99.060 235.840 ;
        RECT 129.270 235.460 131.510 235.840 ;
        RECT 162.315 235.610 162.695 235.990 ;
        RECT 164.355 235.610 164.735 235.990 ;
        RECT 166.140 235.610 166.520 235.990 ;
        RECT 31.925 234.700 34.165 235.080 ;
        RECT 64.375 234.700 66.615 235.080 ;
        RECT 96.825 234.700 99.065 235.080 ;
        RECT 129.275 234.700 131.515 235.080 ;
        RECT 25.200 234.110 25.580 234.490 ;
        RECT 29.120 234.110 29.500 234.490 ;
        RECT 58.180 233.710 58.560 233.760 ;
        RECT 62.520 233.710 62.900 233.760 ;
        RECT 58.180 233.430 62.900 233.710 ;
        RECT 58.180 233.380 58.560 233.430 ;
        RECT 62.520 233.380 62.900 233.430 ;
        RECT 90.630 233.710 91.010 233.760 ;
        RECT 94.970 233.710 95.350 233.760 ;
        RECT 90.630 233.430 95.350 233.710 ;
        RECT 90.630 233.380 91.010 233.430 ;
        RECT 94.970 233.380 95.350 233.430 ;
        RECT 123.080 233.710 123.460 233.760 ;
        RECT 127.420 233.710 127.800 233.760 ;
        RECT 123.080 233.430 127.800 233.710 ;
        RECT 123.080 233.380 123.460 233.430 ;
        RECT 127.420 233.380 127.800 233.430 ;
        RECT 155.530 233.710 155.910 233.760 ;
        RECT 159.870 233.710 160.250 233.760 ;
        RECT 155.530 233.430 160.250 233.710 ;
        RECT 155.530 233.380 155.910 233.430 ;
        RECT 159.870 233.380 160.250 233.430 ;
        RECT 31.920 232.820 34.160 233.200 ;
        RECT 64.370 232.820 66.610 233.200 ;
        RECT 96.820 232.820 99.060 233.200 ;
        RECT 129.270 232.820 131.510 233.200 ;
        RECT 162.315 232.610 162.695 232.990 ;
        RECT 164.355 232.610 164.735 232.990 ;
        RECT 166.140 232.610 166.520 232.990 ;
        RECT 56.900 231.870 57.280 231.920 ;
        RECT 62.520 231.870 62.900 231.920 ;
        RECT 56.900 231.590 62.900 231.870 ;
        RECT 56.900 231.540 57.280 231.590 ;
        RECT 62.520 231.540 62.900 231.590 ;
        RECT 89.350 231.870 89.730 231.920 ;
        RECT 94.970 231.870 95.350 231.920 ;
        RECT 89.350 231.590 95.350 231.870 ;
        RECT 89.350 231.540 89.730 231.590 ;
        RECT 94.970 231.540 95.350 231.590 ;
        RECT 121.800 231.870 122.180 231.920 ;
        RECT 127.420 231.870 127.800 231.920 ;
        RECT 121.800 231.590 127.800 231.870 ;
        RECT 121.800 231.540 122.180 231.590 ;
        RECT 127.420 231.540 127.800 231.590 ;
        RECT 154.250 231.870 154.630 231.920 ;
        RECT 159.870 231.870 160.250 231.920 ;
        RECT 154.250 231.590 160.250 231.870 ;
        RECT 154.250 231.540 154.630 231.590 ;
        RECT 159.870 231.540 160.250 231.590 ;
        RECT 25.200 231.110 25.580 231.490 ;
        RECT 29.120 231.110 29.500 231.490 ;
        RECT 31.920 230.980 34.160 231.360 ;
        RECT 64.370 230.980 66.610 231.360 ;
        RECT 96.820 230.980 99.060 231.360 ;
        RECT 129.270 230.980 131.510 231.360 ;
        RECT 55.620 230.025 56.000 230.075 ;
        RECT 62.520 230.025 62.900 230.075 ;
        RECT 55.620 229.745 62.900 230.025 ;
        RECT 55.620 229.695 56.000 229.745 ;
        RECT 62.520 229.695 62.900 229.745 ;
        RECT 88.070 230.025 88.450 230.075 ;
        RECT 94.970 230.025 95.350 230.075 ;
        RECT 88.070 229.745 95.350 230.025 ;
        RECT 88.070 229.695 88.450 229.745 ;
        RECT 94.970 229.695 95.350 229.745 ;
        RECT 120.520 230.025 120.900 230.075 ;
        RECT 127.420 230.025 127.800 230.075 ;
        RECT 120.520 229.745 127.800 230.025 ;
        RECT 120.520 229.695 120.900 229.745 ;
        RECT 127.420 229.695 127.800 229.745 ;
        RECT 152.970 230.025 153.350 230.075 ;
        RECT 159.870 230.025 160.250 230.075 ;
        RECT 152.970 229.745 160.250 230.025 ;
        RECT 152.970 229.695 153.350 229.745 ;
        RECT 159.870 229.695 160.250 229.745 ;
        RECT 162.315 229.610 162.695 229.990 ;
        RECT 164.355 229.610 164.735 229.990 ;
        RECT 166.140 229.610 166.520 229.990 ;
        RECT 31.920 229.135 34.160 229.515 ;
        RECT 64.370 229.135 66.610 229.515 ;
        RECT 96.820 229.135 99.060 229.515 ;
        RECT 129.270 229.135 131.510 229.515 ;
        RECT 25.200 228.110 25.580 228.490 ;
        RECT 29.120 228.110 29.500 228.490 ;
        RECT 31.925 228.375 34.165 228.755 ;
        RECT 64.375 228.375 66.615 228.755 ;
        RECT 96.825 228.375 99.065 228.755 ;
        RECT 129.275 228.375 131.515 228.755 ;
        RECT 54.340 227.385 54.720 227.435 ;
        RECT 62.520 227.385 62.900 227.435 ;
        RECT 54.340 227.105 62.900 227.385 ;
        RECT 54.340 227.055 54.720 227.105 ;
        RECT 62.520 227.055 62.900 227.105 ;
        RECT 86.790 227.385 87.170 227.435 ;
        RECT 94.970 227.385 95.350 227.435 ;
        RECT 86.790 227.105 95.350 227.385 ;
        RECT 86.790 227.055 87.170 227.105 ;
        RECT 94.970 227.055 95.350 227.105 ;
        RECT 119.240 227.385 119.620 227.435 ;
        RECT 127.420 227.385 127.800 227.435 ;
        RECT 119.240 227.105 127.800 227.385 ;
        RECT 119.240 227.055 119.620 227.105 ;
        RECT 127.420 227.055 127.800 227.105 ;
        RECT 151.690 227.385 152.070 227.435 ;
        RECT 159.870 227.385 160.250 227.435 ;
        RECT 151.690 227.105 160.250 227.385 ;
        RECT 151.690 227.055 152.070 227.105 ;
        RECT 159.870 227.055 160.250 227.105 ;
        RECT 31.920 226.495 34.160 226.875 ;
        RECT 64.370 226.495 66.610 226.875 ;
        RECT 96.820 226.495 99.060 226.875 ;
        RECT 129.270 226.495 131.510 226.875 ;
        RECT 162.315 226.610 162.695 226.990 ;
        RECT 164.355 226.610 164.735 226.990 ;
        RECT 166.140 226.610 166.520 226.990 ;
        RECT 53.060 225.545 53.440 225.595 ;
        RECT 62.520 225.545 62.900 225.595 ;
        RECT 25.200 225.110 25.580 225.490 ;
        RECT 29.120 225.110 29.500 225.490 ;
        RECT 53.060 225.265 62.900 225.545 ;
        RECT 53.060 225.215 53.440 225.265 ;
        RECT 62.520 225.215 62.900 225.265 ;
        RECT 85.510 225.545 85.890 225.595 ;
        RECT 94.970 225.545 95.350 225.595 ;
        RECT 85.510 225.265 95.350 225.545 ;
        RECT 85.510 225.215 85.890 225.265 ;
        RECT 94.970 225.215 95.350 225.265 ;
        RECT 117.960 225.545 118.340 225.595 ;
        RECT 127.420 225.545 127.800 225.595 ;
        RECT 117.960 225.265 127.800 225.545 ;
        RECT 117.960 225.215 118.340 225.265 ;
        RECT 127.420 225.215 127.800 225.265 ;
        RECT 150.410 225.545 150.790 225.595 ;
        RECT 159.870 225.545 160.250 225.595 ;
        RECT 150.410 225.265 160.250 225.545 ;
        RECT 150.410 225.215 150.790 225.265 ;
        RECT 159.870 225.215 160.250 225.265 ;
        RECT 31.920 224.655 34.160 225.035 ;
        RECT 64.370 224.655 66.610 225.035 ;
        RECT 96.820 224.655 99.060 225.035 ;
        RECT 129.270 224.655 131.510 225.035 ;
        RECT 31.920 223.935 34.160 224.315 ;
        RECT 64.370 223.935 66.610 224.315 ;
        RECT 96.820 223.935 99.060 224.315 ;
        RECT 129.270 223.935 131.510 224.315 ;
        RECT 53.700 223.705 54.080 223.755 ;
        RECT 62.520 223.705 62.900 223.755 ;
        RECT 53.700 223.425 62.900 223.705 ;
        RECT 53.700 223.375 54.080 223.425 ;
        RECT 62.520 223.375 62.900 223.425 ;
        RECT 86.150 223.705 86.530 223.755 ;
        RECT 94.970 223.705 95.350 223.755 ;
        RECT 86.150 223.425 95.350 223.705 ;
        RECT 86.150 223.375 86.530 223.425 ;
        RECT 94.970 223.375 95.350 223.425 ;
        RECT 118.600 223.705 118.980 223.755 ;
        RECT 127.420 223.705 127.800 223.755 ;
        RECT 118.600 223.425 127.800 223.705 ;
        RECT 118.600 223.375 118.980 223.425 ;
        RECT 127.420 223.375 127.800 223.425 ;
        RECT 151.050 223.705 151.430 223.755 ;
        RECT 159.870 223.705 160.250 223.755 ;
        RECT 151.050 223.425 160.250 223.705 ;
        RECT 151.050 223.375 151.430 223.425 ;
        RECT 159.870 223.375 160.250 223.425 ;
        RECT 25.200 221.725 25.580 222.105 ;
        RECT 29.120 221.725 29.500 222.105 ;
        RECT 31.920 222.095 34.160 222.475 ;
        RECT 64.370 222.095 66.610 222.475 ;
        RECT 96.820 222.095 99.060 222.475 ;
        RECT 129.270 222.095 131.510 222.475 ;
        RECT 54.980 221.865 55.360 221.915 ;
        RECT 62.520 221.865 62.900 221.915 ;
        RECT 54.980 221.585 62.900 221.865 ;
        RECT 54.980 221.535 55.360 221.585 ;
        RECT 62.520 221.535 62.900 221.585 ;
        RECT 87.430 221.865 87.810 221.915 ;
        RECT 94.970 221.865 95.350 221.915 ;
        RECT 87.430 221.585 95.350 221.865 ;
        RECT 87.430 221.535 87.810 221.585 ;
        RECT 94.970 221.535 95.350 221.585 ;
        RECT 119.880 221.865 120.260 221.915 ;
        RECT 127.420 221.865 127.800 221.915 ;
        RECT 119.880 221.585 127.800 221.865 ;
        RECT 119.880 221.535 120.260 221.585 ;
        RECT 127.420 221.535 127.800 221.585 ;
        RECT 152.330 221.865 152.710 221.915 ;
        RECT 159.870 221.865 160.250 221.915 ;
        RECT 152.330 221.585 160.250 221.865 ;
        RECT 152.330 221.535 152.710 221.585 ;
        RECT 159.870 221.535 160.250 221.585 ;
        RECT 31.925 220.210 34.165 220.590 ;
        RECT 64.375 220.210 66.615 220.590 ;
        RECT 96.825 220.210 99.065 220.590 ;
        RECT 129.275 220.210 131.515 220.590 ;
        RECT 162.315 220.225 162.695 220.605 ;
        RECT 164.355 220.225 164.735 220.605 ;
        RECT 166.140 220.225 166.520 220.605 ;
        RECT 31.920 219.450 34.160 219.830 ;
        RECT 64.370 219.450 66.610 219.830 ;
        RECT 96.820 219.450 99.060 219.830 ;
        RECT 129.270 219.450 131.510 219.830 ;
        RECT 56.260 219.220 56.640 219.270 ;
        RECT 62.520 219.220 62.900 219.270 ;
        RECT 25.200 218.725 25.580 219.105 ;
        RECT 29.120 218.725 29.500 219.105 ;
        RECT 56.260 218.940 62.900 219.220 ;
        RECT 56.260 218.890 56.640 218.940 ;
        RECT 62.520 218.890 62.900 218.940 ;
        RECT 88.710 219.220 89.090 219.270 ;
        RECT 94.970 219.220 95.350 219.270 ;
        RECT 88.710 218.940 95.350 219.220 ;
        RECT 88.710 218.890 89.090 218.940 ;
        RECT 94.970 218.890 95.350 218.940 ;
        RECT 121.160 219.220 121.540 219.270 ;
        RECT 127.420 219.220 127.800 219.270 ;
        RECT 121.160 218.940 127.800 219.220 ;
        RECT 121.160 218.890 121.540 218.940 ;
        RECT 127.420 218.890 127.800 218.940 ;
        RECT 153.610 219.220 153.990 219.270 ;
        RECT 159.870 219.220 160.250 219.270 ;
        RECT 153.610 218.940 160.250 219.220 ;
        RECT 153.610 218.890 153.990 218.940 ;
        RECT 159.870 218.890 160.250 218.940 ;
        RECT 31.920 217.610 34.160 217.990 ;
        RECT 64.370 217.610 66.610 217.990 ;
        RECT 96.820 217.610 99.060 217.990 ;
        RECT 129.270 217.610 131.510 217.990 ;
        RECT 57.540 217.380 57.920 217.430 ;
        RECT 62.520 217.380 62.900 217.430 ;
        RECT 57.540 217.100 62.900 217.380 ;
        RECT 57.540 217.050 57.920 217.100 ;
        RECT 62.520 217.050 62.900 217.100 ;
        RECT 89.990 217.380 90.370 217.430 ;
        RECT 94.970 217.380 95.350 217.430 ;
        RECT 89.990 217.100 95.350 217.380 ;
        RECT 89.990 217.050 90.370 217.100 ;
        RECT 94.970 217.050 95.350 217.100 ;
        RECT 122.440 217.380 122.820 217.430 ;
        RECT 127.420 217.380 127.800 217.430 ;
        RECT 122.440 217.100 127.800 217.380 ;
        RECT 122.440 217.050 122.820 217.100 ;
        RECT 127.420 217.050 127.800 217.100 ;
        RECT 154.890 217.380 155.270 217.430 ;
        RECT 159.870 217.380 160.250 217.430 ;
        RECT 154.890 217.100 160.250 217.380 ;
        RECT 162.315 217.225 162.695 217.605 ;
        RECT 164.355 217.225 164.735 217.605 ;
        RECT 166.140 217.225 166.520 217.605 ;
        RECT 154.890 217.050 155.270 217.100 ;
        RECT 159.870 217.050 160.250 217.100 ;
        RECT 25.200 215.725 25.580 216.105 ;
        RECT 29.120 215.725 29.500 216.105 ;
        RECT 31.920 215.770 34.160 216.150 ;
        RECT 64.370 215.770 66.610 216.150 ;
        RECT 96.820 215.770 99.060 216.150 ;
        RECT 129.270 215.770 131.510 216.150 ;
        RECT 58.820 215.540 59.200 215.590 ;
        RECT 62.520 215.540 62.900 215.590 ;
        RECT 58.820 215.260 62.900 215.540 ;
        RECT 58.820 215.210 59.200 215.260 ;
        RECT 62.520 215.210 62.900 215.260 ;
        RECT 91.270 215.540 91.650 215.590 ;
        RECT 94.970 215.540 95.350 215.590 ;
        RECT 91.270 215.260 95.350 215.540 ;
        RECT 91.270 215.210 91.650 215.260 ;
        RECT 94.970 215.210 95.350 215.260 ;
        RECT 123.720 215.540 124.100 215.590 ;
        RECT 127.420 215.540 127.800 215.590 ;
        RECT 123.720 215.260 127.800 215.540 ;
        RECT 123.720 215.210 124.100 215.260 ;
        RECT 127.420 215.210 127.800 215.260 ;
        RECT 156.170 215.540 156.550 215.590 ;
        RECT 159.870 215.540 160.250 215.590 ;
        RECT 156.170 215.260 160.250 215.540 ;
        RECT 156.170 215.210 156.550 215.260 ;
        RECT 159.870 215.210 160.250 215.260 ;
        RECT 31.925 213.885 34.165 214.265 ;
        RECT 64.375 213.885 66.615 214.265 ;
        RECT 96.825 213.885 99.065 214.265 ;
        RECT 129.275 213.885 131.515 214.265 ;
        RECT 162.315 214.225 162.695 214.605 ;
        RECT 164.355 214.225 164.735 214.605 ;
        RECT 166.140 214.225 166.520 214.605 ;
        RECT 31.920 213.125 34.160 213.505 ;
        RECT 64.370 213.125 66.610 213.505 ;
        RECT 96.820 213.125 99.060 213.505 ;
        RECT 129.270 213.125 131.510 213.505 ;
        RECT 25.200 212.725 25.580 213.105 ;
        RECT 29.120 212.725 29.500 213.105 ;
        RECT 60.100 212.895 60.480 212.945 ;
        RECT 62.520 212.895 62.900 212.945 ;
        RECT 60.100 212.615 62.900 212.895 ;
        RECT 60.100 212.565 60.480 212.615 ;
        RECT 62.520 212.565 62.900 212.615 ;
        RECT 92.550 212.895 92.930 212.945 ;
        RECT 94.970 212.895 95.350 212.945 ;
        RECT 92.550 212.615 95.350 212.895 ;
        RECT 92.550 212.565 92.930 212.615 ;
        RECT 94.970 212.565 95.350 212.615 ;
        RECT 125.000 212.895 125.380 212.945 ;
        RECT 127.420 212.895 127.800 212.945 ;
        RECT 125.000 212.615 127.800 212.895 ;
        RECT 125.000 212.565 125.380 212.615 ;
        RECT 127.420 212.565 127.800 212.615 ;
        RECT 157.450 212.895 157.830 212.945 ;
        RECT 159.870 212.895 160.250 212.945 ;
        RECT 157.450 212.615 160.250 212.895 ;
        RECT 157.450 212.565 157.830 212.615 ;
        RECT 159.870 212.565 160.250 212.615 ;
        RECT 31.920 211.285 34.160 211.665 ;
        RECT 64.370 211.285 66.610 211.665 ;
        RECT 96.820 211.285 99.060 211.665 ;
        RECT 129.270 211.285 131.510 211.665 ;
        RECT 162.315 211.225 162.695 211.605 ;
        RECT 164.355 211.225 164.735 211.605 ;
        RECT 166.140 211.225 166.520 211.605 ;
        RECT 61.380 211.055 61.760 211.105 ;
        RECT 62.520 211.055 62.900 211.105 ;
        RECT 61.380 210.775 62.900 211.055 ;
        RECT 61.380 210.725 61.760 210.775 ;
        RECT 62.520 210.725 62.900 210.775 ;
        RECT 93.830 211.055 94.210 211.105 ;
        RECT 94.970 211.055 95.350 211.105 ;
        RECT 93.830 210.775 95.350 211.055 ;
        RECT 93.830 210.725 94.210 210.775 ;
        RECT 94.970 210.725 95.350 210.775 ;
        RECT 126.280 211.055 126.660 211.105 ;
        RECT 127.420 211.055 127.800 211.105 ;
        RECT 126.280 210.775 127.800 211.055 ;
        RECT 126.280 210.725 126.660 210.775 ;
        RECT 127.420 210.725 127.800 210.775 ;
        RECT 158.730 211.055 159.110 211.105 ;
        RECT 159.870 211.055 160.250 211.105 ;
        RECT 158.730 210.775 160.250 211.055 ;
        RECT 158.730 210.725 159.110 210.775 ;
        RECT 159.870 210.725 160.250 210.775 ;
        RECT 25.200 209.725 25.580 210.105 ;
        RECT 29.120 209.725 29.500 210.105 ;
        RECT 31.920 209.445 34.160 209.825 ;
        RECT 64.370 209.445 66.610 209.825 ;
        RECT 96.820 209.445 99.060 209.825 ;
        RECT 129.270 209.445 131.510 209.825 ;
        RECT 62.520 208.885 63.040 209.265 ;
        RECT 94.970 208.885 95.490 209.265 ;
        RECT 127.420 208.885 127.940 209.265 ;
        RECT 159.870 208.885 160.390 209.265 ;
        RECT 162.315 208.225 162.695 208.605 ;
        RECT 164.355 208.225 164.735 208.605 ;
        RECT 166.140 208.225 166.520 208.605 ;
        RECT 25.200 206.725 25.580 207.105 ;
        RECT 29.120 206.725 29.500 207.105 ;
        RECT 25.200 203.725 25.580 204.105 ;
        RECT 162.315 202.225 162.695 202.605 ;
        RECT 164.355 202.225 164.735 202.605 ;
        RECT 166.140 202.225 166.520 202.605 ;
        RECT 25.200 200.725 25.580 201.105 ;
        RECT 29.120 200.725 29.500 201.105 ;
        RECT 62.020 200.320 62.900 200.700 ;
        RECT 94.470 200.320 95.350 200.700 ;
        RECT 126.920 200.320 127.800 200.700 ;
        RECT 159.370 200.320 160.250 200.700 ;
        RECT 31.920 199.760 34.160 200.140 ;
        RECT 64.370 199.760 66.610 200.140 ;
        RECT 96.820 199.760 99.060 200.140 ;
        RECT 129.270 199.760 131.510 200.140 ;
        RECT 162.315 199.225 162.695 199.605 ;
        RECT 164.355 199.225 164.735 199.605 ;
        RECT 166.140 199.225 166.520 199.605 ;
        RECT 60.740 198.810 61.120 198.860 ;
        RECT 62.520 198.810 62.900 198.860 ;
        RECT 60.740 198.530 62.900 198.810 ;
        RECT 60.740 198.480 61.120 198.530 ;
        RECT 62.520 198.480 62.900 198.530 ;
        RECT 93.190 198.810 93.570 198.860 ;
        RECT 94.970 198.810 95.350 198.860 ;
        RECT 93.190 198.530 95.350 198.810 ;
        RECT 93.190 198.480 93.570 198.530 ;
        RECT 94.970 198.480 95.350 198.530 ;
        RECT 125.640 198.810 126.020 198.860 ;
        RECT 127.420 198.810 127.800 198.860 ;
        RECT 125.640 198.530 127.800 198.810 ;
        RECT 125.640 198.480 126.020 198.530 ;
        RECT 127.420 198.480 127.800 198.530 ;
        RECT 158.090 198.810 158.470 198.860 ;
        RECT 159.870 198.810 160.250 198.860 ;
        RECT 158.090 198.530 160.250 198.810 ;
        RECT 158.090 198.480 158.470 198.530 ;
        RECT 159.870 198.480 160.250 198.530 ;
        RECT 25.200 197.725 25.580 198.105 ;
        RECT 29.120 197.725 29.500 198.105 ;
        RECT 31.920 197.920 34.160 198.300 ;
        RECT 64.370 197.920 66.610 198.300 ;
        RECT 96.820 197.920 99.060 198.300 ;
        RECT 129.270 197.920 131.510 198.300 ;
        RECT 59.460 196.965 59.840 197.015 ;
        RECT 62.520 196.965 62.900 197.015 ;
        RECT 59.460 196.685 62.900 196.965 ;
        RECT 59.460 196.635 59.840 196.685 ;
        RECT 62.520 196.635 62.900 196.685 ;
        RECT 91.910 196.965 92.290 197.015 ;
        RECT 94.970 196.965 95.350 197.015 ;
        RECT 91.910 196.685 95.350 196.965 ;
        RECT 91.910 196.635 92.290 196.685 ;
        RECT 94.970 196.635 95.350 196.685 ;
        RECT 124.360 196.965 124.740 197.015 ;
        RECT 127.420 196.965 127.800 197.015 ;
        RECT 124.360 196.685 127.800 196.965 ;
        RECT 124.360 196.635 124.740 196.685 ;
        RECT 127.420 196.635 127.800 196.685 ;
        RECT 156.810 196.965 157.190 197.015 ;
        RECT 159.870 196.965 160.250 197.015 ;
        RECT 156.810 196.685 160.250 196.965 ;
        RECT 156.810 196.635 157.190 196.685 ;
        RECT 159.870 196.635 160.250 196.685 ;
        RECT 31.920 196.075 34.160 196.455 ;
        RECT 64.370 196.075 66.610 196.455 ;
        RECT 96.820 196.075 99.060 196.455 ;
        RECT 129.270 196.075 131.510 196.455 ;
        RECT 162.315 196.225 162.695 196.605 ;
        RECT 164.355 196.225 164.735 196.605 ;
        RECT 166.140 196.225 166.520 196.605 ;
        RECT 31.925 195.315 34.165 195.695 ;
        RECT 64.375 195.315 66.615 195.695 ;
        RECT 96.825 195.315 99.065 195.695 ;
        RECT 129.275 195.315 131.515 195.695 ;
        RECT 25.200 194.725 25.580 195.105 ;
        RECT 29.120 194.725 29.500 195.105 ;
        RECT 58.180 194.325 58.560 194.375 ;
        RECT 62.520 194.325 62.900 194.375 ;
        RECT 58.180 194.045 62.900 194.325 ;
        RECT 58.180 193.995 58.560 194.045 ;
        RECT 62.520 193.995 62.900 194.045 ;
        RECT 90.630 194.325 91.010 194.375 ;
        RECT 94.970 194.325 95.350 194.375 ;
        RECT 90.630 194.045 95.350 194.325 ;
        RECT 90.630 193.995 91.010 194.045 ;
        RECT 94.970 193.995 95.350 194.045 ;
        RECT 123.080 194.325 123.460 194.375 ;
        RECT 127.420 194.325 127.800 194.375 ;
        RECT 123.080 194.045 127.800 194.325 ;
        RECT 123.080 193.995 123.460 194.045 ;
        RECT 127.420 193.995 127.800 194.045 ;
        RECT 155.530 194.325 155.910 194.375 ;
        RECT 159.870 194.325 160.250 194.375 ;
        RECT 155.530 194.045 160.250 194.325 ;
        RECT 155.530 193.995 155.910 194.045 ;
        RECT 159.870 193.995 160.250 194.045 ;
        RECT 31.920 193.435 34.160 193.815 ;
        RECT 64.370 193.435 66.610 193.815 ;
        RECT 96.820 193.435 99.060 193.815 ;
        RECT 129.270 193.435 131.510 193.815 ;
        RECT 162.315 193.225 162.695 193.605 ;
        RECT 164.355 193.225 164.735 193.605 ;
        RECT 166.140 193.225 166.520 193.605 ;
        RECT 56.900 192.485 57.280 192.535 ;
        RECT 62.520 192.485 62.900 192.535 ;
        RECT 56.900 192.205 62.900 192.485 ;
        RECT 56.900 192.155 57.280 192.205 ;
        RECT 62.520 192.155 62.900 192.205 ;
        RECT 89.350 192.485 89.730 192.535 ;
        RECT 94.970 192.485 95.350 192.535 ;
        RECT 89.350 192.205 95.350 192.485 ;
        RECT 89.350 192.155 89.730 192.205 ;
        RECT 94.970 192.155 95.350 192.205 ;
        RECT 121.800 192.485 122.180 192.535 ;
        RECT 127.420 192.485 127.800 192.535 ;
        RECT 121.800 192.205 127.800 192.485 ;
        RECT 121.800 192.155 122.180 192.205 ;
        RECT 127.420 192.155 127.800 192.205 ;
        RECT 154.250 192.485 154.630 192.535 ;
        RECT 159.870 192.485 160.250 192.535 ;
        RECT 154.250 192.205 160.250 192.485 ;
        RECT 154.250 192.155 154.630 192.205 ;
        RECT 159.870 192.155 160.250 192.205 ;
        RECT 25.200 191.725 25.580 192.105 ;
        RECT 29.120 191.725 29.500 192.105 ;
        RECT 31.920 191.595 34.160 191.975 ;
        RECT 64.370 191.595 66.610 191.975 ;
        RECT 96.820 191.595 99.060 191.975 ;
        RECT 129.270 191.595 131.510 191.975 ;
        RECT 55.620 190.640 56.000 190.690 ;
        RECT 62.520 190.640 62.900 190.690 ;
        RECT 55.620 190.360 62.900 190.640 ;
        RECT 55.620 190.310 56.000 190.360 ;
        RECT 62.520 190.310 62.900 190.360 ;
        RECT 88.070 190.640 88.450 190.690 ;
        RECT 94.970 190.640 95.350 190.690 ;
        RECT 88.070 190.360 95.350 190.640 ;
        RECT 88.070 190.310 88.450 190.360 ;
        RECT 94.970 190.310 95.350 190.360 ;
        RECT 120.520 190.640 120.900 190.690 ;
        RECT 127.420 190.640 127.800 190.690 ;
        RECT 120.520 190.360 127.800 190.640 ;
        RECT 120.520 190.310 120.900 190.360 ;
        RECT 127.420 190.310 127.800 190.360 ;
        RECT 152.970 190.640 153.350 190.690 ;
        RECT 159.870 190.640 160.250 190.690 ;
        RECT 152.970 190.360 160.250 190.640 ;
        RECT 152.970 190.310 153.350 190.360 ;
        RECT 159.870 190.310 160.250 190.360 ;
        RECT 162.315 190.225 162.695 190.605 ;
        RECT 164.355 190.225 164.735 190.605 ;
        RECT 166.140 190.225 166.520 190.605 ;
        RECT 31.920 189.750 34.160 190.130 ;
        RECT 64.370 189.750 66.610 190.130 ;
        RECT 96.820 189.750 99.060 190.130 ;
        RECT 129.270 189.750 131.510 190.130 ;
        RECT 25.200 188.725 25.580 189.105 ;
        RECT 29.120 188.725 29.500 189.105 ;
        RECT 31.925 188.990 34.165 189.370 ;
        RECT 64.375 188.990 66.615 189.370 ;
        RECT 96.825 188.990 99.065 189.370 ;
        RECT 129.275 188.990 131.515 189.370 ;
        RECT 54.340 188.000 54.720 188.050 ;
        RECT 62.520 188.000 62.900 188.050 ;
        RECT 54.340 187.720 62.900 188.000 ;
        RECT 54.340 187.670 54.720 187.720 ;
        RECT 62.520 187.670 62.900 187.720 ;
        RECT 86.790 188.000 87.170 188.050 ;
        RECT 94.970 188.000 95.350 188.050 ;
        RECT 86.790 187.720 95.350 188.000 ;
        RECT 86.790 187.670 87.170 187.720 ;
        RECT 94.970 187.670 95.350 187.720 ;
        RECT 119.240 188.000 119.620 188.050 ;
        RECT 127.420 188.000 127.800 188.050 ;
        RECT 119.240 187.720 127.800 188.000 ;
        RECT 119.240 187.670 119.620 187.720 ;
        RECT 127.420 187.670 127.800 187.720 ;
        RECT 151.690 188.000 152.070 188.050 ;
        RECT 159.870 188.000 160.250 188.050 ;
        RECT 151.690 187.720 160.250 188.000 ;
        RECT 151.690 187.670 152.070 187.720 ;
        RECT 159.870 187.670 160.250 187.720 ;
        RECT 31.920 187.110 34.160 187.490 ;
        RECT 64.370 187.110 66.610 187.490 ;
        RECT 96.820 187.110 99.060 187.490 ;
        RECT 129.270 187.110 131.510 187.490 ;
        RECT 162.315 187.225 162.695 187.605 ;
        RECT 164.355 187.225 164.735 187.605 ;
        RECT 166.140 187.225 166.520 187.605 ;
        RECT 53.060 186.160 53.440 186.210 ;
        RECT 62.520 186.160 62.900 186.210 ;
        RECT 25.200 185.725 25.580 186.105 ;
        RECT 29.120 185.725 29.500 186.105 ;
        RECT 53.060 185.880 62.900 186.160 ;
        RECT 53.060 185.830 53.440 185.880 ;
        RECT 62.520 185.830 62.900 185.880 ;
        RECT 85.510 186.160 85.890 186.210 ;
        RECT 94.970 186.160 95.350 186.210 ;
        RECT 85.510 185.880 95.350 186.160 ;
        RECT 85.510 185.830 85.890 185.880 ;
        RECT 94.970 185.830 95.350 185.880 ;
        RECT 117.960 186.160 118.340 186.210 ;
        RECT 127.420 186.160 127.800 186.210 ;
        RECT 117.960 185.880 127.800 186.160 ;
        RECT 117.960 185.830 118.340 185.880 ;
        RECT 127.420 185.830 127.800 185.880 ;
        RECT 150.410 186.160 150.790 186.210 ;
        RECT 159.870 186.160 160.250 186.210 ;
        RECT 150.410 185.880 160.250 186.160 ;
        RECT 150.410 185.830 150.790 185.880 ;
        RECT 159.870 185.830 160.250 185.880 ;
        RECT 31.920 185.270 34.160 185.650 ;
        RECT 64.370 185.270 66.610 185.650 ;
        RECT 96.820 185.270 99.060 185.650 ;
        RECT 129.270 185.270 131.510 185.650 ;
        RECT 31.920 184.550 34.160 184.930 ;
        RECT 64.370 184.550 66.610 184.930 ;
        RECT 96.820 184.550 99.060 184.930 ;
        RECT 129.270 184.550 131.510 184.930 ;
        RECT 53.700 184.320 54.080 184.370 ;
        RECT 62.520 184.320 62.900 184.370 ;
        RECT 53.700 184.040 62.900 184.320 ;
        RECT 53.700 183.990 54.080 184.040 ;
        RECT 62.520 183.990 62.900 184.040 ;
        RECT 86.150 184.320 86.530 184.370 ;
        RECT 94.970 184.320 95.350 184.370 ;
        RECT 86.150 184.040 95.350 184.320 ;
        RECT 86.150 183.990 86.530 184.040 ;
        RECT 94.970 183.990 95.350 184.040 ;
        RECT 118.600 184.320 118.980 184.370 ;
        RECT 127.420 184.320 127.800 184.370 ;
        RECT 118.600 184.040 127.800 184.320 ;
        RECT 118.600 183.990 118.980 184.040 ;
        RECT 127.420 183.990 127.800 184.040 ;
        RECT 151.050 184.320 151.430 184.370 ;
        RECT 159.870 184.320 160.250 184.370 ;
        RECT 151.050 184.040 160.250 184.320 ;
        RECT 151.050 183.990 151.430 184.040 ;
        RECT 159.870 183.990 160.250 184.040 ;
        RECT 25.200 182.340 25.580 182.720 ;
        RECT 29.120 182.340 29.500 182.720 ;
        RECT 31.920 182.710 34.160 183.090 ;
        RECT 64.370 182.710 66.610 183.090 ;
        RECT 96.820 182.710 99.060 183.090 ;
        RECT 129.270 182.710 131.510 183.090 ;
        RECT 54.980 182.480 55.360 182.530 ;
        RECT 62.520 182.480 62.900 182.530 ;
        RECT 54.980 182.200 62.900 182.480 ;
        RECT 54.980 182.150 55.360 182.200 ;
        RECT 62.520 182.150 62.900 182.200 ;
        RECT 87.430 182.480 87.810 182.530 ;
        RECT 94.970 182.480 95.350 182.530 ;
        RECT 87.430 182.200 95.350 182.480 ;
        RECT 87.430 182.150 87.810 182.200 ;
        RECT 94.970 182.150 95.350 182.200 ;
        RECT 119.880 182.480 120.260 182.530 ;
        RECT 127.420 182.480 127.800 182.530 ;
        RECT 119.880 182.200 127.800 182.480 ;
        RECT 119.880 182.150 120.260 182.200 ;
        RECT 127.420 182.150 127.800 182.200 ;
        RECT 152.330 182.480 152.710 182.530 ;
        RECT 159.870 182.480 160.250 182.530 ;
        RECT 152.330 182.200 160.250 182.480 ;
        RECT 152.330 182.150 152.710 182.200 ;
        RECT 159.870 182.150 160.250 182.200 ;
        RECT 31.925 180.825 34.165 181.205 ;
        RECT 64.375 180.825 66.615 181.205 ;
        RECT 96.825 180.825 99.065 181.205 ;
        RECT 129.275 180.825 131.515 181.205 ;
        RECT 162.315 180.840 162.695 181.220 ;
        RECT 164.355 180.840 164.735 181.220 ;
        RECT 166.140 180.840 166.520 181.220 ;
        RECT 31.920 180.065 34.160 180.445 ;
        RECT 64.370 180.065 66.610 180.445 ;
        RECT 96.820 180.065 99.060 180.445 ;
        RECT 129.270 180.065 131.510 180.445 ;
        RECT 56.260 179.835 56.640 179.885 ;
        RECT 62.520 179.835 62.900 179.885 ;
        RECT 25.200 179.340 25.580 179.720 ;
        RECT 29.120 179.340 29.500 179.720 ;
        RECT 56.260 179.555 62.900 179.835 ;
        RECT 56.260 179.505 56.640 179.555 ;
        RECT 62.520 179.505 62.900 179.555 ;
        RECT 88.710 179.835 89.090 179.885 ;
        RECT 94.970 179.835 95.350 179.885 ;
        RECT 88.710 179.555 95.350 179.835 ;
        RECT 88.710 179.505 89.090 179.555 ;
        RECT 94.970 179.505 95.350 179.555 ;
        RECT 121.160 179.835 121.540 179.885 ;
        RECT 127.420 179.835 127.800 179.885 ;
        RECT 121.160 179.555 127.800 179.835 ;
        RECT 121.160 179.505 121.540 179.555 ;
        RECT 127.420 179.505 127.800 179.555 ;
        RECT 153.610 179.835 153.990 179.885 ;
        RECT 159.870 179.835 160.250 179.885 ;
        RECT 153.610 179.555 160.250 179.835 ;
        RECT 153.610 179.505 153.990 179.555 ;
        RECT 159.870 179.505 160.250 179.555 ;
        RECT 31.920 178.225 34.160 178.605 ;
        RECT 64.370 178.225 66.610 178.605 ;
        RECT 96.820 178.225 99.060 178.605 ;
        RECT 129.270 178.225 131.510 178.605 ;
        RECT 57.540 177.995 57.920 178.045 ;
        RECT 62.520 177.995 62.900 178.045 ;
        RECT 57.540 177.715 62.900 177.995 ;
        RECT 57.540 177.665 57.920 177.715 ;
        RECT 62.520 177.665 62.900 177.715 ;
        RECT 89.990 177.995 90.370 178.045 ;
        RECT 94.970 177.995 95.350 178.045 ;
        RECT 89.990 177.715 95.350 177.995 ;
        RECT 89.990 177.665 90.370 177.715 ;
        RECT 94.970 177.665 95.350 177.715 ;
        RECT 122.440 177.995 122.820 178.045 ;
        RECT 127.420 177.995 127.800 178.045 ;
        RECT 122.440 177.715 127.800 177.995 ;
        RECT 122.440 177.665 122.820 177.715 ;
        RECT 127.420 177.665 127.800 177.715 ;
        RECT 154.890 177.995 155.270 178.045 ;
        RECT 159.870 177.995 160.250 178.045 ;
        RECT 154.890 177.715 160.250 177.995 ;
        RECT 162.315 177.840 162.695 178.220 ;
        RECT 164.355 177.840 164.735 178.220 ;
        RECT 166.140 177.840 166.520 178.220 ;
        RECT 154.890 177.665 155.270 177.715 ;
        RECT 159.870 177.665 160.250 177.715 ;
        RECT 25.200 176.340 25.580 176.720 ;
        RECT 29.120 176.340 29.500 176.720 ;
        RECT 31.920 176.385 34.160 176.765 ;
        RECT 64.370 176.385 66.610 176.765 ;
        RECT 96.820 176.385 99.060 176.765 ;
        RECT 129.270 176.385 131.510 176.765 ;
        RECT 58.820 176.155 59.200 176.205 ;
        RECT 62.520 176.155 62.900 176.205 ;
        RECT 58.820 175.875 62.900 176.155 ;
        RECT 58.820 175.825 59.200 175.875 ;
        RECT 62.520 175.825 62.900 175.875 ;
        RECT 91.270 176.155 91.650 176.205 ;
        RECT 94.970 176.155 95.350 176.205 ;
        RECT 91.270 175.875 95.350 176.155 ;
        RECT 91.270 175.825 91.650 175.875 ;
        RECT 94.970 175.825 95.350 175.875 ;
        RECT 123.720 176.155 124.100 176.205 ;
        RECT 127.420 176.155 127.800 176.205 ;
        RECT 123.720 175.875 127.800 176.155 ;
        RECT 123.720 175.825 124.100 175.875 ;
        RECT 127.420 175.825 127.800 175.875 ;
        RECT 156.170 176.155 156.550 176.205 ;
        RECT 159.870 176.155 160.250 176.205 ;
        RECT 156.170 175.875 160.250 176.155 ;
        RECT 156.170 175.825 156.550 175.875 ;
        RECT 159.870 175.825 160.250 175.875 ;
        RECT 31.925 174.500 34.165 174.880 ;
        RECT 64.375 174.500 66.615 174.880 ;
        RECT 96.825 174.500 99.065 174.880 ;
        RECT 129.275 174.500 131.515 174.880 ;
        RECT 162.315 174.840 162.695 175.220 ;
        RECT 164.355 174.840 164.735 175.220 ;
        RECT 166.140 174.840 166.520 175.220 ;
        RECT 31.920 173.740 34.160 174.120 ;
        RECT 64.370 173.740 66.610 174.120 ;
        RECT 96.820 173.740 99.060 174.120 ;
        RECT 129.270 173.740 131.510 174.120 ;
        RECT 25.200 173.340 25.580 173.720 ;
        RECT 29.120 173.340 29.500 173.720 ;
        RECT 60.100 173.510 60.480 173.560 ;
        RECT 62.520 173.510 62.900 173.560 ;
        RECT 60.100 173.230 62.900 173.510 ;
        RECT 60.100 173.180 60.480 173.230 ;
        RECT 62.520 173.180 62.900 173.230 ;
        RECT 92.550 173.510 92.930 173.560 ;
        RECT 94.970 173.510 95.350 173.560 ;
        RECT 92.550 173.230 95.350 173.510 ;
        RECT 92.550 173.180 92.930 173.230 ;
        RECT 94.970 173.180 95.350 173.230 ;
        RECT 125.000 173.510 125.380 173.560 ;
        RECT 127.420 173.510 127.800 173.560 ;
        RECT 125.000 173.230 127.800 173.510 ;
        RECT 125.000 173.180 125.380 173.230 ;
        RECT 127.420 173.180 127.800 173.230 ;
        RECT 157.450 173.510 157.830 173.560 ;
        RECT 159.870 173.510 160.250 173.560 ;
        RECT 157.450 173.230 160.250 173.510 ;
        RECT 157.450 173.180 157.830 173.230 ;
        RECT 159.870 173.180 160.250 173.230 ;
        RECT 31.920 171.900 34.160 172.280 ;
        RECT 64.370 171.900 66.610 172.280 ;
        RECT 96.820 171.900 99.060 172.280 ;
        RECT 129.270 171.900 131.510 172.280 ;
        RECT 162.315 171.840 162.695 172.220 ;
        RECT 164.355 171.840 164.735 172.220 ;
        RECT 166.140 171.840 166.520 172.220 ;
        RECT 61.380 171.670 61.760 171.720 ;
        RECT 62.520 171.670 62.900 171.720 ;
        RECT 61.380 171.390 62.900 171.670 ;
        RECT 61.380 171.340 61.760 171.390 ;
        RECT 62.520 171.340 62.900 171.390 ;
        RECT 93.830 171.670 94.210 171.720 ;
        RECT 94.970 171.670 95.350 171.720 ;
        RECT 93.830 171.390 95.350 171.670 ;
        RECT 93.830 171.340 94.210 171.390 ;
        RECT 94.970 171.340 95.350 171.390 ;
        RECT 126.280 171.670 126.660 171.720 ;
        RECT 127.420 171.670 127.800 171.720 ;
        RECT 126.280 171.390 127.800 171.670 ;
        RECT 126.280 171.340 126.660 171.390 ;
        RECT 127.420 171.340 127.800 171.390 ;
        RECT 158.730 171.670 159.110 171.720 ;
        RECT 159.870 171.670 160.250 171.720 ;
        RECT 158.730 171.390 160.250 171.670 ;
        RECT 158.730 171.340 159.110 171.390 ;
        RECT 159.870 171.340 160.250 171.390 ;
        RECT 25.200 170.340 25.580 170.720 ;
        RECT 29.120 170.340 29.500 170.720 ;
        RECT 31.920 170.060 34.160 170.440 ;
        RECT 64.370 170.060 66.610 170.440 ;
        RECT 96.820 170.060 99.060 170.440 ;
        RECT 129.270 170.060 131.510 170.440 ;
        RECT 62.520 169.500 63.040 169.880 ;
        RECT 94.970 169.500 95.490 169.880 ;
        RECT 127.420 169.500 127.940 169.880 ;
        RECT 159.870 169.500 160.390 169.880 ;
        RECT 162.315 168.840 162.695 169.220 ;
        RECT 164.355 168.840 164.735 169.220 ;
        RECT 166.140 168.840 166.520 169.220 ;
        RECT 25.200 167.340 25.580 167.720 ;
        RECT 29.120 167.340 29.500 167.720 ;
        RECT 25.200 164.340 25.580 164.720 ;
        RECT 162.315 162.840 162.695 163.220 ;
        RECT 164.355 162.840 164.735 163.220 ;
        RECT 166.140 162.840 166.520 163.220 ;
        RECT 25.200 161.340 25.580 161.720 ;
        RECT 29.120 161.340 29.500 161.720 ;
        RECT 62.020 160.935 62.900 161.315 ;
        RECT 94.470 160.935 95.350 161.315 ;
        RECT 126.920 160.935 127.800 161.315 ;
        RECT 159.370 160.935 160.250 161.315 ;
        RECT 31.920 160.375 34.160 160.755 ;
        RECT 64.370 160.375 66.610 160.755 ;
        RECT 96.820 160.375 99.060 160.755 ;
        RECT 129.270 160.375 131.510 160.755 ;
        RECT 162.315 159.840 162.695 160.220 ;
        RECT 164.355 159.840 164.735 160.220 ;
        RECT 166.140 159.840 166.520 160.220 ;
        RECT 60.740 159.425 61.120 159.475 ;
        RECT 62.520 159.425 62.900 159.475 ;
        RECT 60.740 159.145 62.900 159.425 ;
        RECT 60.740 159.095 61.120 159.145 ;
        RECT 62.520 159.095 62.900 159.145 ;
        RECT 93.190 159.425 93.570 159.475 ;
        RECT 94.970 159.425 95.350 159.475 ;
        RECT 93.190 159.145 95.350 159.425 ;
        RECT 93.190 159.095 93.570 159.145 ;
        RECT 94.970 159.095 95.350 159.145 ;
        RECT 125.640 159.425 126.020 159.475 ;
        RECT 127.420 159.425 127.800 159.475 ;
        RECT 125.640 159.145 127.800 159.425 ;
        RECT 125.640 159.095 126.020 159.145 ;
        RECT 127.420 159.095 127.800 159.145 ;
        RECT 158.090 159.425 158.470 159.475 ;
        RECT 159.870 159.425 160.250 159.475 ;
        RECT 158.090 159.145 160.250 159.425 ;
        RECT 158.090 159.095 158.470 159.145 ;
        RECT 159.870 159.095 160.250 159.145 ;
        RECT 25.200 158.340 25.580 158.720 ;
        RECT 29.120 158.340 29.500 158.720 ;
        RECT 31.920 158.535 34.160 158.915 ;
        RECT 64.370 158.535 66.610 158.915 ;
        RECT 96.820 158.535 99.060 158.915 ;
        RECT 129.270 158.535 131.510 158.915 ;
        RECT 59.460 157.580 59.840 157.630 ;
        RECT 62.520 157.580 62.900 157.630 ;
        RECT 59.460 157.300 62.900 157.580 ;
        RECT 59.460 157.250 59.840 157.300 ;
        RECT 62.520 157.250 62.900 157.300 ;
        RECT 91.910 157.580 92.290 157.630 ;
        RECT 94.970 157.580 95.350 157.630 ;
        RECT 91.910 157.300 95.350 157.580 ;
        RECT 91.910 157.250 92.290 157.300 ;
        RECT 94.970 157.250 95.350 157.300 ;
        RECT 124.360 157.580 124.740 157.630 ;
        RECT 127.420 157.580 127.800 157.630 ;
        RECT 124.360 157.300 127.800 157.580 ;
        RECT 124.360 157.250 124.740 157.300 ;
        RECT 127.420 157.250 127.800 157.300 ;
        RECT 156.810 157.580 157.190 157.630 ;
        RECT 159.870 157.580 160.250 157.630 ;
        RECT 156.810 157.300 160.250 157.580 ;
        RECT 156.810 157.250 157.190 157.300 ;
        RECT 159.870 157.250 160.250 157.300 ;
        RECT 31.920 156.690 34.160 157.070 ;
        RECT 64.370 156.690 66.610 157.070 ;
        RECT 96.820 156.690 99.060 157.070 ;
        RECT 129.270 156.690 131.510 157.070 ;
        RECT 162.315 156.840 162.695 157.220 ;
        RECT 164.355 156.840 164.735 157.220 ;
        RECT 166.140 156.840 166.520 157.220 ;
        RECT 31.925 155.930 34.165 156.310 ;
        RECT 64.375 155.930 66.615 156.310 ;
        RECT 96.825 155.930 99.065 156.310 ;
        RECT 129.275 155.930 131.515 156.310 ;
        RECT 25.200 155.340 25.580 155.720 ;
        RECT 29.120 155.340 29.500 155.720 ;
        RECT 58.180 154.940 58.560 154.990 ;
        RECT 62.520 154.940 62.900 154.990 ;
        RECT 58.180 154.660 62.900 154.940 ;
        RECT 58.180 154.610 58.560 154.660 ;
        RECT 62.520 154.610 62.900 154.660 ;
        RECT 90.630 154.940 91.010 154.990 ;
        RECT 94.970 154.940 95.350 154.990 ;
        RECT 90.630 154.660 95.350 154.940 ;
        RECT 90.630 154.610 91.010 154.660 ;
        RECT 94.970 154.610 95.350 154.660 ;
        RECT 123.080 154.940 123.460 154.990 ;
        RECT 127.420 154.940 127.800 154.990 ;
        RECT 123.080 154.660 127.800 154.940 ;
        RECT 123.080 154.610 123.460 154.660 ;
        RECT 127.420 154.610 127.800 154.660 ;
        RECT 155.530 154.940 155.910 154.990 ;
        RECT 159.870 154.940 160.250 154.990 ;
        RECT 155.530 154.660 160.250 154.940 ;
        RECT 155.530 154.610 155.910 154.660 ;
        RECT 159.870 154.610 160.250 154.660 ;
        RECT 31.920 154.050 34.160 154.430 ;
        RECT 64.370 154.050 66.610 154.430 ;
        RECT 96.820 154.050 99.060 154.430 ;
        RECT 129.270 154.050 131.510 154.430 ;
        RECT 162.315 153.840 162.695 154.220 ;
        RECT 164.355 153.840 164.735 154.220 ;
        RECT 166.140 153.840 166.520 154.220 ;
        RECT 56.900 153.100 57.280 153.150 ;
        RECT 62.520 153.100 62.900 153.150 ;
        RECT 56.900 152.820 62.900 153.100 ;
        RECT 56.900 152.770 57.280 152.820 ;
        RECT 62.520 152.770 62.900 152.820 ;
        RECT 89.350 153.100 89.730 153.150 ;
        RECT 94.970 153.100 95.350 153.150 ;
        RECT 89.350 152.820 95.350 153.100 ;
        RECT 89.350 152.770 89.730 152.820 ;
        RECT 94.970 152.770 95.350 152.820 ;
        RECT 121.800 153.100 122.180 153.150 ;
        RECT 127.420 153.100 127.800 153.150 ;
        RECT 121.800 152.820 127.800 153.100 ;
        RECT 121.800 152.770 122.180 152.820 ;
        RECT 127.420 152.770 127.800 152.820 ;
        RECT 154.250 153.100 154.630 153.150 ;
        RECT 159.870 153.100 160.250 153.150 ;
        RECT 154.250 152.820 160.250 153.100 ;
        RECT 154.250 152.770 154.630 152.820 ;
        RECT 159.870 152.770 160.250 152.820 ;
        RECT 25.200 152.340 25.580 152.720 ;
        RECT 29.120 152.340 29.500 152.720 ;
        RECT 31.920 152.210 34.160 152.590 ;
        RECT 64.370 152.210 66.610 152.590 ;
        RECT 96.820 152.210 99.060 152.590 ;
        RECT 129.270 152.210 131.510 152.590 ;
        RECT 55.620 151.255 56.000 151.305 ;
        RECT 62.520 151.255 62.900 151.305 ;
        RECT 55.620 150.975 62.900 151.255 ;
        RECT 55.620 150.925 56.000 150.975 ;
        RECT 62.520 150.925 62.900 150.975 ;
        RECT 88.070 151.255 88.450 151.305 ;
        RECT 94.970 151.255 95.350 151.305 ;
        RECT 88.070 150.975 95.350 151.255 ;
        RECT 88.070 150.925 88.450 150.975 ;
        RECT 94.970 150.925 95.350 150.975 ;
        RECT 120.520 151.255 120.900 151.305 ;
        RECT 127.420 151.255 127.800 151.305 ;
        RECT 120.520 150.975 127.800 151.255 ;
        RECT 120.520 150.925 120.900 150.975 ;
        RECT 127.420 150.925 127.800 150.975 ;
        RECT 152.970 151.255 153.350 151.305 ;
        RECT 159.870 151.255 160.250 151.305 ;
        RECT 152.970 150.975 160.250 151.255 ;
        RECT 152.970 150.925 153.350 150.975 ;
        RECT 159.870 150.925 160.250 150.975 ;
        RECT 162.315 150.840 162.695 151.220 ;
        RECT 164.355 150.840 164.735 151.220 ;
        RECT 166.140 150.840 166.520 151.220 ;
        RECT 31.920 150.365 34.160 150.745 ;
        RECT 64.370 150.365 66.610 150.745 ;
        RECT 96.820 150.365 99.060 150.745 ;
        RECT 129.270 150.365 131.510 150.745 ;
        RECT 25.200 149.340 25.580 149.720 ;
        RECT 29.120 149.340 29.500 149.720 ;
        RECT 31.925 149.605 34.165 149.985 ;
        RECT 64.375 149.605 66.615 149.985 ;
        RECT 96.825 149.605 99.065 149.985 ;
        RECT 129.275 149.605 131.515 149.985 ;
        RECT 54.340 148.615 54.720 148.665 ;
        RECT 62.520 148.615 62.900 148.665 ;
        RECT 54.340 148.335 62.900 148.615 ;
        RECT 54.340 148.285 54.720 148.335 ;
        RECT 62.520 148.285 62.900 148.335 ;
        RECT 86.790 148.615 87.170 148.665 ;
        RECT 94.970 148.615 95.350 148.665 ;
        RECT 86.790 148.335 95.350 148.615 ;
        RECT 86.790 148.285 87.170 148.335 ;
        RECT 94.970 148.285 95.350 148.335 ;
        RECT 119.240 148.615 119.620 148.665 ;
        RECT 127.420 148.615 127.800 148.665 ;
        RECT 119.240 148.335 127.800 148.615 ;
        RECT 119.240 148.285 119.620 148.335 ;
        RECT 127.420 148.285 127.800 148.335 ;
        RECT 151.690 148.615 152.070 148.665 ;
        RECT 159.870 148.615 160.250 148.665 ;
        RECT 151.690 148.335 160.250 148.615 ;
        RECT 151.690 148.285 152.070 148.335 ;
        RECT 159.870 148.285 160.250 148.335 ;
        RECT 31.920 147.725 34.160 148.105 ;
        RECT 64.370 147.725 66.610 148.105 ;
        RECT 96.820 147.725 99.060 148.105 ;
        RECT 129.270 147.725 131.510 148.105 ;
        RECT 162.315 147.840 162.695 148.220 ;
        RECT 164.355 147.840 164.735 148.220 ;
        RECT 166.140 147.840 166.520 148.220 ;
        RECT 53.060 146.775 53.440 146.825 ;
        RECT 62.520 146.775 62.900 146.825 ;
        RECT 25.200 146.340 25.580 146.720 ;
        RECT 29.120 146.340 29.500 146.720 ;
        RECT 53.060 146.495 62.900 146.775 ;
        RECT 53.060 146.445 53.440 146.495 ;
        RECT 62.520 146.445 62.900 146.495 ;
        RECT 85.510 146.775 85.890 146.825 ;
        RECT 94.970 146.775 95.350 146.825 ;
        RECT 85.510 146.495 95.350 146.775 ;
        RECT 85.510 146.445 85.890 146.495 ;
        RECT 94.970 146.445 95.350 146.495 ;
        RECT 117.960 146.775 118.340 146.825 ;
        RECT 127.420 146.775 127.800 146.825 ;
        RECT 117.960 146.495 127.800 146.775 ;
        RECT 117.960 146.445 118.340 146.495 ;
        RECT 127.420 146.445 127.800 146.495 ;
        RECT 150.410 146.775 150.790 146.825 ;
        RECT 159.870 146.775 160.250 146.825 ;
        RECT 150.410 146.495 160.250 146.775 ;
        RECT 150.410 146.445 150.790 146.495 ;
        RECT 159.870 146.445 160.250 146.495 ;
        RECT 31.920 145.885 34.160 146.265 ;
        RECT 64.370 145.885 66.610 146.265 ;
        RECT 96.820 145.885 99.060 146.265 ;
        RECT 129.270 145.885 131.510 146.265 ;
        RECT 31.920 145.165 34.160 145.545 ;
        RECT 64.370 145.165 66.610 145.545 ;
        RECT 96.820 145.165 99.060 145.545 ;
        RECT 129.270 145.165 131.510 145.545 ;
        RECT 53.700 144.935 54.080 144.985 ;
        RECT 62.520 144.935 62.900 144.985 ;
        RECT 53.700 144.655 62.900 144.935 ;
        RECT 53.700 144.605 54.080 144.655 ;
        RECT 62.520 144.605 62.900 144.655 ;
        RECT 86.150 144.935 86.530 144.985 ;
        RECT 94.970 144.935 95.350 144.985 ;
        RECT 86.150 144.655 95.350 144.935 ;
        RECT 86.150 144.605 86.530 144.655 ;
        RECT 94.970 144.605 95.350 144.655 ;
        RECT 118.600 144.935 118.980 144.985 ;
        RECT 127.420 144.935 127.800 144.985 ;
        RECT 118.600 144.655 127.800 144.935 ;
        RECT 118.600 144.605 118.980 144.655 ;
        RECT 127.420 144.605 127.800 144.655 ;
        RECT 151.050 144.935 151.430 144.985 ;
        RECT 159.870 144.935 160.250 144.985 ;
        RECT 151.050 144.655 160.250 144.935 ;
        RECT 151.050 144.605 151.430 144.655 ;
        RECT 159.870 144.605 160.250 144.655 ;
        RECT 25.200 142.955 25.580 143.335 ;
        RECT 29.120 142.955 29.500 143.335 ;
        RECT 31.920 143.325 34.160 143.705 ;
        RECT 64.370 143.325 66.610 143.705 ;
        RECT 96.820 143.325 99.060 143.705 ;
        RECT 129.270 143.325 131.510 143.705 ;
        RECT 54.980 143.095 55.360 143.145 ;
        RECT 62.520 143.095 62.900 143.145 ;
        RECT 54.980 142.815 62.900 143.095 ;
        RECT 54.980 142.765 55.360 142.815 ;
        RECT 62.520 142.765 62.900 142.815 ;
        RECT 87.430 143.095 87.810 143.145 ;
        RECT 94.970 143.095 95.350 143.145 ;
        RECT 87.430 142.815 95.350 143.095 ;
        RECT 87.430 142.765 87.810 142.815 ;
        RECT 94.970 142.765 95.350 142.815 ;
        RECT 119.880 143.095 120.260 143.145 ;
        RECT 127.420 143.095 127.800 143.145 ;
        RECT 119.880 142.815 127.800 143.095 ;
        RECT 119.880 142.765 120.260 142.815 ;
        RECT 127.420 142.765 127.800 142.815 ;
        RECT 152.330 143.095 152.710 143.145 ;
        RECT 159.870 143.095 160.250 143.145 ;
        RECT 152.330 142.815 160.250 143.095 ;
        RECT 152.330 142.765 152.710 142.815 ;
        RECT 159.870 142.765 160.250 142.815 ;
        RECT 31.925 141.440 34.165 141.820 ;
        RECT 64.375 141.440 66.615 141.820 ;
        RECT 96.825 141.440 99.065 141.820 ;
        RECT 129.275 141.440 131.515 141.820 ;
        RECT 162.315 141.455 162.695 141.835 ;
        RECT 164.355 141.455 164.735 141.835 ;
        RECT 166.140 141.455 166.520 141.835 ;
        RECT 31.920 140.680 34.160 141.060 ;
        RECT 64.370 140.680 66.610 141.060 ;
        RECT 96.820 140.680 99.060 141.060 ;
        RECT 129.270 140.680 131.510 141.060 ;
        RECT 56.260 140.450 56.640 140.500 ;
        RECT 62.520 140.450 62.900 140.500 ;
        RECT 25.200 139.955 25.580 140.335 ;
        RECT 29.120 139.955 29.500 140.335 ;
        RECT 56.260 140.170 62.900 140.450 ;
        RECT 56.260 140.120 56.640 140.170 ;
        RECT 62.520 140.120 62.900 140.170 ;
        RECT 88.710 140.450 89.090 140.500 ;
        RECT 94.970 140.450 95.350 140.500 ;
        RECT 88.710 140.170 95.350 140.450 ;
        RECT 88.710 140.120 89.090 140.170 ;
        RECT 94.970 140.120 95.350 140.170 ;
        RECT 121.160 140.450 121.540 140.500 ;
        RECT 127.420 140.450 127.800 140.500 ;
        RECT 121.160 140.170 127.800 140.450 ;
        RECT 121.160 140.120 121.540 140.170 ;
        RECT 127.420 140.120 127.800 140.170 ;
        RECT 153.610 140.450 153.990 140.500 ;
        RECT 159.870 140.450 160.250 140.500 ;
        RECT 153.610 140.170 160.250 140.450 ;
        RECT 153.610 140.120 153.990 140.170 ;
        RECT 159.870 140.120 160.250 140.170 ;
        RECT 31.920 138.840 34.160 139.220 ;
        RECT 64.370 138.840 66.610 139.220 ;
        RECT 96.820 138.840 99.060 139.220 ;
        RECT 129.270 138.840 131.510 139.220 ;
        RECT 57.540 138.610 57.920 138.660 ;
        RECT 62.520 138.610 62.900 138.660 ;
        RECT 57.540 138.330 62.900 138.610 ;
        RECT 57.540 138.280 57.920 138.330 ;
        RECT 62.520 138.280 62.900 138.330 ;
        RECT 89.990 138.610 90.370 138.660 ;
        RECT 94.970 138.610 95.350 138.660 ;
        RECT 89.990 138.330 95.350 138.610 ;
        RECT 89.990 138.280 90.370 138.330 ;
        RECT 94.970 138.280 95.350 138.330 ;
        RECT 122.440 138.610 122.820 138.660 ;
        RECT 127.420 138.610 127.800 138.660 ;
        RECT 122.440 138.330 127.800 138.610 ;
        RECT 122.440 138.280 122.820 138.330 ;
        RECT 127.420 138.280 127.800 138.330 ;
        RECT 154.890 138.610 155.270 138.660 ;
        RECT 159.870 138.610 160.250 138.660 ;
        RECT 154.890 138.330 160.250 138.610 ;
        RECT 162.315 138.455 162.695 138.835 ;
        RECT 164.355 138.455 164.735 138.835 ;
        RECT 166.140 138.455 166.520 138.835 ;
        RECT 154.890 138.280 155.270 138.330 ;
        RECT 159.870 138.280 160.250 138.330 ;
        RECT 25.200 136.955 25.580 137.335 ;
        RECT 29.120 136.955 29.500 137.335 ;
        RECT 31.920 137.000 34.160 137.380 ;
        RECT 64.370 137.000 66.610 137.380 ;
        RECT 96.820 137.000 99.060 137.380 ;
        RECT 129.270 137.000 131.510 137.380 ;
        RECT 58.820 136.770 59.200 136.820 ;
        RECT 62.520 136.770 62.900 136.820 ;
        RECT 58.820 136.490 62.900 136.770 ;
        RECT 58.820 136.440 59.200 136.490 ;
        RECT 62.520 136.440 62.900 136.490 ;
        RECT 91.270 136.770 91.650 136.820 ;
        RECT 94.970 136.770 95.350 136.820 ;
        RECT 91.270 136.490 95.350 136.770 ;
        RECT 91.270 136.440 91.650 136.490 ;
        RECT 94.970 136.440 95.350 136.490 ;
        RECT 123.720 136.770 124.100 136.820 ;
        RECT 127.420 136.770 127.800 136.820 ;
        RECT 123.720 136.490 127.800 136.770 ;
        RECT 123.720 136.440 124.100 136.490 ;
        RECT 127.420 136.440 127.800 136.490 ;
        RECT 156.170 136.770 156.550 136.820 ;
        RECT 159.870 136.770 160.250 136.820 ;
        RECT 156.170 136.490 160.250 136.770 ;
        RECT 156.170 136.440 156.550 136.490 ;
        RECT 159.870 136.440 160.250 136.490 ;
        RECT 31.925 135.115 34.165 135.495 ;
        RECT 64.375 135.115 66.615 135.495 ;
        RECT 96.825 135.115 99.065 135.495 ;
        RECT 129.275 135.115 131.515 135.495 ;
        RECT 162.315 135.455 162.695 135.835 ;
        RECT 164.355 135.455 164.735 135.835 ;
        RECT 166.140 135.455 166.520 135.835 ;
        RECT 31.920 134.355 34.160 134.735 ;
        RECT 64.370 134.355 66.610 134.735 ;
        RECT 96.820 134.355 99.060 134.735 ;
        RECT 129.270 134.355 131.510 134.735 ;
        RECT 25.200 133.955 25.580 134.335 ;
        RECT 29.120 133.955 29.500 134.335 ;
        RECT 60.100 134.125 60.480 134.175 ;
        RECT 62.520 134.125 62.900 134.175 ;
        RECT 60.100 133.845 62.900 134.125 ;
        RECT 60.100 133.795 60.480 133.845 ;
        RECT 62.520 133.795 62.900 133.845 ;
        RECT 92.550 134.125 92.930 134.175 ;
        RECT 94.970 134.125 95.350 134.175 ;
        RECT 92.550 133.845 95.350 134.125 ;
        RECT 92.550 133.795 92.930 133.845 ;
        RECT 94.970 133.795 95.350 133.845 ;
        RECT 125.000 134.125 125.380 134.175 ;
        RECT 127.420 134.125 127.800 134.175 ;
        RECT 125.000 133.845 127.800 134.125 ;
        RECT 125.000 133.795 125.380 133.845 ;
        RECT 127.420 133.795 127.800 133.845 ;
        RECT 157.450 134.125 157.830 134.175 ;
        RECT 159.870 134.125 160.250 134.175 ;
        RECT 157.450 133.845 160.250 134.125 ;
        RECT 157.450 133.795 157.830 133.845 ;
        RECT 159.870 133.795 160.250 133.845 ;
        RECT 31.920 132.515 34.160 132.895 ;
        RECT 64.370 132.515 66.610 132.895 ;
        RECT 96.820 132.515 99.060 132.895 ;
        RECT 129.270 132.515 131.510 132.895 ;
        RECT 162.315 132.455 162.695 132.835 ;
        RECT 164.355 132.455 164.735 132.835 ;
        RECT 166.140 132.455 166.520 132.835 ;
        RECT 61.380 132.285 61.760 132.335 ;
        RECT 62.520 132.285 62.900 132.335 ;
        RECT 61.380 132.005 62.900 132.285 ;
        RECT 61.380 131.955 61.760 132.005 ;
        RECT 62.520 131.955 62.900 132.005 ;
        RECT 93.830 132.285 94.210 132.335 ;
        RECT 94.970 132.285 95.350 132.335 ;
        RECT 93.830 132.005 95.350 132.285 ;
        RECT 93.830 131.955 94.210 132.005 ;
        RECT 94.970 131.955 95.350 132.005 ;
        RECT 126.280 132.285 126.660 132.335 ;
        RECT 127.420 132.285 127.800 132.335 ;
        RECT 126.280 132.005 127.800 132.285 ;
        RECT 126.280 131.955 126.660 132.005 ;
        RECT 127.420 131.955 127.800 132.005 ;
        RECT 158.730 132.285 159.110 132.335 ;
        RECT 159.870 132.285 160.250 132.335 ;
        RECT 158.730 132.005 160.250 132.285 ;
        RECT 158.730 131.955 159.110 132.005 ;
        RECT 159.870 131.955 160.250 132.005 ;
        RECT 25.200 130.955 25.580 131.335 ;
        RECT 29.120 130.955 29.500 131.335 ;
        RECT 31.920 130.675 34.160 131.055 ;
        RECT 64.370 130.675 66.610 131.055 ;
        RECT 96.820 130.675 99.060 131.055 ;
        RECT 129.270 130.675 131.510 131.055 ;
        RECT 62.520 130.115 63.040 130.495 ;
        RECT 94.970 130.115 95.490 130.495 ;
        RECT 127.420 130.115 127.940 130.495 ;
        RECT 159.870 130.115 160.390 130.495 ;
        RECT 162.315 129.455 162.695 129.835 ;
        RECT 164.355 129.455 164.735 129.835 ;
        RECT 166.140 129.455 166.520 129.835 ;
        RECT 25.200 127.955 25.580 128.335 ;
        RECT 29.120 127.955 29.500 128.335 ;
        RECT 25.200 124.955 25.580 125.335 ;
        RECT 162.315 123.455 162.695 123.835 ;
        RECT 164.355 123.455 164.735 123.835 ;
        RECT 166.140 123.455 166.520 123.835 ;
        RECT 25.200 121.955 25.580 122.335 ;
        RECT 29.120 121.955 29.500 122.335 ;
        RECT 62.020 121.550 62.900 121.930 ;
        RECT 94.470 121.550 95.350 121.930 ;
        RECT 126.920 121.550 127.800 121.930 ;
        RECT 159.370 121.550 160.250 121.930 ;
        RECT 31.920 120.990 34.160 121.370 ;
        RECT 64.370 120.990 66.610 121.370 ;
        RECT 96.820 120.990 99.060 121.370 ;
        RECT 129.270 120.990 131.510 121.370 ;
        RECT 162.315 120.455 162.695 120.835 ;
        RECT 164.355 120.455 164.735 120.835 ;
        RECT 166.140 120.455 166.520 120.835 ;
        RECT 60.740 120.040 61.120 120.090 ;
        RECT 62.520 120.040 62.900 120.090 ;
        RECT 60.740 119.760 62.900 120.040 ;
        RECT 60.740 119.710 61.120 119.760 ;
        RECT 62.520 119.710 62.900 119.760 ;
        RECT 93.190 120.040 93.570 120.090 ;
        RECT 94.970 120.040 95.350 120.090 ;
        RECT 93.190 119.760 95.350 120.040 ;
        RECT 93.190 119.710 93.570 119.760 ;
        RECT 94.970 119.710 95.350 119.760 ;
        RECT 125.640 120.040 126.020 120.090 ;
        RECT 127.420 120.040 127.800 120.090 ;
        RECT 125.640 119.760 127.800 120.040 ;
        RECT 125.640 119.710 126.020 119.760 ;
        RECT 127.420 119.710 127.800 119.760 ;
        RECT 158.090 120.040 158.470 120.090 ;
        RECT 159.870 120.040 160.250 120.090 ;
        RECT 158.090 119.760 160.250 120.040 ;
        RECT 158.090 119.710 158.470 119.760 ;
        RECT 159.870 119.710 160.250 119.760 ;
        RECT 25.200 118.955 25.580 119.335 ;
        RECT 29.120 118.955 29.500 119.335 ;
        RECT 31.920 119.150 34.160 119.530 ;
        RECT 64.370 119.150 66.610 119.530 ;
        RECT 96.820 119.150 99.060 119.530 ;
        RECT 129.270 119.150 131.510 119.530 ;
        RECT 59.460 118.195 59.840 118.245 ;
        RECT 62.520 118.195 62.900 118.245 ;
        RECT 59.460 117.915 62.900 118.195 ;
        RECT 59.460 117.865 59.840 117.915 ;
        RECT 62.520 117.865 62.900 117.915 ;
        RECT 91.910 118.195 92.290 118.245 ;
        RECT 94.970 118.195 95.350 118.245 ;
        RECT 91.910 117.915 95.350 118.195 ;
        RECT 91.910 117.865 92.290 117.915 ;
        RECT 94.970 117.865 95.350 117.915 ;
        RECT 124.360 118.195 124.740 118.245 ;
        RECT 127.420 118.195 127.800 118.245 ;
        RECT 124.360 117.915 127.800 118.195 ;
        RECT 124.360 117.865 124.740 117.915 ;
        RECT 127.420 117.865 127.800 117.915 ;
        RECT 156.810 118.195 157.190 118.245 ;
        RECT 159.870 118.195 160.250 118.245 ;
        RECT 156.810 117.915 160.250 118.195 ;
        RECT 156.810 117.865 157.190 117.915 ;
        RECT 159.870 117.865 160.250 117.915 ;
        RECT 31.920 117.305 34.160 117.685 ;
        RECT 64.370 117.305 66.610 117.685 ;
        RECT 96.820 117.305 99.060 117.685 ;
        RECT 129.270 117.305 131.510 117.685 ;
        RECT 162.315 117.455 162.695 117.835 ;
        RECT 164.355 117.455 164.735 117.835 ;
        RECT 166.140 117.455 166.520 117.835 ;
        RECT 31.925 116.545 34.165 116.925 ;
        RECT 64.375 116.545 66.615 116.925 ;
        RECT 96.825 116.545 99.065 116.925 ;
        RECT 129.275 116.545 131.515 116.925 ;
        RECT 25.200 115.955 25.580 116.335 ;
        RECT 29.120 115.955 29.500 116.335 ;
        RECT 58.180 115.555 58.560 115.605 ;
        RECT 62.520 115.555 62.900 115.605 ;
        RECT 58.180 115.275 62.900 115.555 ;
        RECT 58.180 115.225 58.560 115.275 ;
        RECT 62.520 115.225 62.900 115.275 ;
        RECT 90.630 115.555 91.010 115.605 ;
        RECT 94.970 115.555 95.350 115.605 ;
        RECT 90.630 115.275 95.350 115.555 ;
        RECT 90.630 115.225 91.010 115.275 ;
        RECT 94.970 115.225 95.350 115.275 ;
        RECT 123.080 115.555 123.460 115.605 ;
        RECT 127.420 115.555 127.800 115.605 ;
        RECT 123.080 115.275 127.800 115.555 ;
        RECT 123.080 115.225 123.460 115.275 ;
        RECT 127.420 115.225 127.800 115.275 ;
        RECT 155.530 115.555 155.910 115.605 ;
        RECT 159.870 115.555 160.250 115.605 ;
        RECT 155.530 115.275 160.250 115.555 ;
        RECT 155.530 115.225 155.910 115.275 ;
        RECT 159.870 115.225 160.250 115.275 ;
        RECT 31.920 114.665 34.160 115.045 ;
        RECT 64.370 114.665 66.610 115.045 ;
        RECT 96.820 114.665 99.060 115.045 ;
        RECT 129.270 114.665 131.510 115.045 ;
        RECT 162.315 114.455 162.695 114.835 ;
        RECT 164.355 114.455 164.735 114.835 ;
        RECT 166.140 114.455 166.520 114.835 ;
        RECT 56.900 113.715 57.280 113.765 ;
        RECT 62.520 113.715 62.900 113.765 ;
        RECT 56.900 113.435 62.900 113.715 ;
        RECT 56.900 113.385 57.280 113.435 ;
        RECT 62.520 113.385 62.900 113.435 ;
        RECT 89.350 113.715 89.730 113.765 ;
        RECT 94.970 113.715 95.350 113.765 ;
        RECT 89.350 113.435 95.350 113.715 ;
        RECT 89.350 113.385 89.730 113.435 ;
        RECT 94.970 113.385 95.350 113.435 ;
        RECT 121.800 113.715 122.180 113.765 ;
        RECT 127.420 113.715 127.800 113.765 ;
        RECT 121.800 113.435 127.800 113.715 ;
        RECT 121.800 113.385 122.180 113.435 ;
        RECT 127.420 113.385 127.800 113.435 ;
        RECT 154.250 113.715 154.630 113.765 ;
        RECT 159.870 113.715 160.250 113.765 ;
        RECT 154.250 113.435 160.250 113.715 ;
        RECT 154.250 113.385 154.630 113.435 ;
        RECT 159.870 113.385 160.250 113.435 ;
        RECT 25.200 112.955 25.580 113.335 ;
        RECT 29.120 112.955 29.500 113.335 ;
        RECT 31.920 112.825 34.160 113.205 ;
        RECT 64.370 112.825 66.610 113.205 ;
        RECT 96.820 112.825 99.060 113.205 ;
        RECT 129.270 112.825 131.510 113.205 ;
        RECT 55.620 111.870 56.000 111.920 ;
        RECT 62.520 111.870 62.900 111.920 ;
        RECT 55.620 111.590 62.900 111.870 ;
        RECT 55.620 111.540 56.000 111.590 ;
        RECT 62.520 111.540 62.900 111.590 ;
        RECT 88.070 111.870 88.450 111.920 ;
        RECT 94.970 111.870 95.350 111.920 ;
        RECT 88.070 111.590 95.350 111.870 ;
        RECT 88.070 111.540 88.450 111.590 ;
        RECT 94.970 111.540 95.350 111.590 ;
        RECT 120.520 111.870 120.900 111.920 ;
        RECT 127.420 111.870 127.800 111.920 ;
        RECT 120.520 111.590 127.800 111.870 ;
        RECT 120.520 111.540 120.900 111.590 ;
        RECT 127.420 111.540 127.800 111.590 ;
        RECT 152.970 111.870 153.350 111.920 ;
        RECT 159.870 111.870 160.250 111.920 ;
        RECT 152.970 111.590 160.250 111.870 ;
        RECT 152.970 111.540 153.350 111.590 ;
        RECT 159.870 111.540 160.250 111.590 ;
        RECT 162.315 111.455 162.695 111.835 ;
        RECT 164.355 111.455 164.735 111.835 ;
        RECT 166.140 111.455 166.520 111.835 ;
        RECT 31.920 110.980 34.160 111.360 ;
        RECT 64.370 110.980 66.610 111.360 ;
        RECT 96.820 110.980 99.060 111.360 ;
        RECT 129.270 110.980 131.510 111.360 ;
        RECT 25.200 109.955 25.580 110.335 ;
        RECT 29.120 109.955 29.500 110.335 ;
        RECT 31.925 110.220 34.165 110.600 ;
        RECT 64.375 110.220 66.615 110.600 ;
        RECT 96.825 110.220 99.065 110.600 ;
        RECT 129.275 110.220 131.515 110.600 ;
        RECT 54.340 109.230 54.720 109.280 ;
        RECT 62.520 109.230 62.900 109.280 ;
        RECT 54.340 108.950 62.900 109.230 ;
        RECT 54.340 108.900 54.720 108.950 ;
        RECT 62.520 108.900 62.900 108.950 ;
        RECT 86.790 109.230 87.170 109.280 ;
        RECT 94.970 109.230 95.350 109.280 ;
        RECT 86.790 108.950 95.350 109.230 ;
        RECT 86.790 108.900 87.170 108.950 ;
        RECT 94.970 108.900 95.350 108.950 ;
        RECT 119.240 109.230 119.620 109.280 ;
        RECT 127.420 109.230 127.800 109.280 ;
        RECT 119.240 108.950 127.800 109.230 ;
        RECT 119.240 108.900 119.620 108.950 ;
        RECT 127.420 108.900 127.800 108.950 ;
        RECT 151.690 109.230 152.070 109.280 ;
        RECT 159.870 109.230 160.250 109.280 ;
        RECT 151.690 108.950 160.250 109.230 ;
        RECT 151.690 108.900 152.070 108.950 ;
        RECT 159.870 108.900 160.250 108.950 ;
        RECT 31.920 108.340 34.160 108.720 ;
        RECT 64.370 108.340 66.610 108.720 ;
        RECT 96.820 108.340 99.060 108.720 ;
        RECT 129.270 108.340 131.510 108.720 ;
        RECT 162.315 108.455 162.695 108.835 ;
        RECT 164.355 108.455 164.735 108.835 ;
        RECT 166.140 108.455 166.520 108.835 ;
        RECT 53.060 107.390 53.440 107.440 ;
        RECT 62.520 107.390 62.900 107.440 ;
        RECT 25.200 106.955 25.580 107.335 ;
        RECT 29.120 106.955 29.500 107.335 ;
        RECT 53.060 107.110 62.900 107.390 ;
        RECT 53.060 107.060 53.440 107.110 ;
        RECT 62.520 107.060 62.900 107.110 ;
        RECT 85.510 107.390 85.890 107.440 ;
        RECT 94.970 107.390 95.350 107.440 ;
        RECT 85.510 107.110 95.350 107.390 ;
        RECT 85.510 107.060 85.890 107.110 ;
        RECT 94.970 107.060 95.350 107.110 ;
        RECT 117.960 107.390 118.340 107.440 ;
        RECT 127.420 107.390 127.800 107.440 ;
        RECT 117.960 107.110 127.800 107.390 ;
        RECT 117.960 107.060 118.340 107.110 ;
        RECT 127.420 107.060 127.800 107.110 ;
        RECT 150.410 107.390 150.790 107.440 ;
        RECT 159.870 107.390 160.250 107.440 ;
        RECT 150.410 107.110 160.250 107.390 ;
        RECT 150.410 107.060 150.790 107.110 ;
        RECT 159.870 107.060 160.250 107.110 ;
        RECT 31.920 106.500 34.160 106.880 ;
        RECT 64.370 106.500 66.610 106.880 ;
        RECT 96.820 106.500 99.060 106.880 ;
        RECT 129.270 106.500 131.510 106.880 ;
        RECT 31.920 105.780 34.160 106.160 ;
        RECT 64.370 105.780 66.610 106.160 ;
        RECT 96.820 105.780 99.060 106.160 ;
        RECT 129.270 105.780 131.510 106.160 ;
        RECT 53.700 105.550 54.080 105.600 ;
        RECT 62.520 105.550 62.900 105.600 ;
        RECT 53.700 105.270 62.900 105.550 ;
        RECT 53.700 105.220 54.080 105.270 ;
        RECT 62.520 105.220 62.900 105.270 ;
        RECT 86.150 105.550 86.530 105.600 ;
        RECT 94.970 105.550 95.350 105.600 ;
        RECT 86.150 105.270 95.350 105.550 ;
        RECT 86.150 105.220 86.530 105.270 ;
        RECT 94.970 105.220 95.350 105.270 ;
        RECT 118.600 105.550 118.980 105.600 ;
        RECT 127.420 105.550 127.800 105.600 ;
        RECT 118.600 105.270 127.800 105.550 ;
        RECT 118.600 105.220 118.980 105.270 ;
        RECT 127.420 105.220 127.800 105.270 ;
        RECT 151.050 105.550 151.430 105.600 ;
        RECT 159.870 105.550 160.250 105.600 ;
        RECT 151.050 105.270 160.250 105.550 ;
        RECT 151.050 105.220 151.430 105.270 ;
        RECT 159.870 105.220 160.250 105.270 ;
        RECT 25.200 103.570 25.580 103.950 ;
        RECT 29.120 103.570 29.500 103.950 ;
        RECT 31.920 103.940 34.160 104.320 ;
        RECT 64.370 103.940 66.610 104.320 ;
        RECT 96.820 103.940 99.060 104.320 ;
        RECT 129.270 103.940 131.510 104.320 ;
        RECT 54.980 103.710 55.360 103.760 ;
        RECT 62.520 103.710 62.900 103.760 ;
        RECT 54.980 103.430 62.900 103.710 ;
        RECT 54.980 103.380 55.360 103.430 ;
        RECT 62.520 103.380 62.900 103.430 ;
        RECT 87.430 103.710 87.810 103.760 ;
        RECT 94.970 103.710 95.350 103.760 ;
        RECT 87.430 103.430 95.350 103.710 ;
        RECT 87.430 103.380 87.810 103.430 ;
        RECT 94.970 103.380 95.350 103.430 ;
        RECT 119.880 103.710 120.260 103.760 ;
        RECT 127.420 103.710 127.800 103.760 ;
        RECT 119.880 103.430 127.800 103.710 ;
        RECT 119.880 103.380 120.260 103.430 ;
        RECT 127.420 103.380 127.800 103.430 ;
        RECT 152.330 103.710 152.710 103.760 ;
        RECT 159.870 103.710 160.250 103.760 ;
        RECT 152.330 103.430 160.250 103.710 ;
        RECT 152.330 103.380 152.710 103.430 ;
        RECT 159.870 103.380 160.250 103.430 ;
        RECT 31.925 102.055 34.165 102.435 ;
        RECT 64.375 102.055 66.615 102.435 ;
        RECT 96.825 102.055 99.065 102.435 ;
        RECT 129.275 102.055 131.515 102.435 ;
        RECT 162.315 102.070 162.695 102.450 ;
        RECT 164.355 102.070 164.735 102.450 ;
        RECT 166.140 102.070 166.520 102.450 ;
        RECT 31.920 101.295 34.160 101.675 ;
        RECT 64.370 101.295 66.610 101.675 ;
        RECT 96.820 101.295 99.060 101.675 ;
        RECT 129.270 101.295 131.510 101.675 ;
        RECT 56.260 101.065 56.640 101.115 ;
        RECT 62.520 101.065 62.900 101.115 ;
        RECT 25.200 100.570 25.580 100.950 ;
        RECT 29.120 100.570 29.500 100.950 ;
        RECT 56.260 100.785 62.900 101.065 ;
        RECT 56.260 100.735 56.640 100.785 ;
        RECT 62.520 100.735 62.900 100.785 ;
        RECT 88.710 101.065 89.090 101.115 ;
        RECT 94.970 101.065 95.350 101.115 ;
        RECT 88.710 100.785 95.350 101.065 ;
        RECT 88.710 100.735 89.090 100.785 ;
        RECT 94.970 100.735 95.350 100.785 ;
        RECT 121.160 101.065 121.540 101.115 ;
        RECT 127.420 101.065 127.800 101.115 ;
        RECT 121.160 100.785 127.800 101.065 ;
        RECT 121.160 100.735 121.540 100.785 ;
        RECT 127.420 100.735 127.800 100.785 ;
        RECT 153.610 101.065 153.990 101.115 ;
        RECT 159.870 101.065 160.250 101.115 ;
        RECT 153.610 100.785 160.250 101.065 ;
        RECT 153.610 100.735 153.990 100.785 ;
        RECT 159.870 100.735 160.250 100.785 ;
        RECT 31.920 99.455 34.160 99.835 ;
        RECT 64.370 99.455 66.610 99.835 ;
        RECT 96.820 99.455 99.060 99.835 ;
        RECT 129.270 99.455 131.510 99.835 ;
        RECT 57.540 99.225 57.920 99.275 ;
        RECT 62.520 99.225 62.900 99.275 ;
        RECT 57.540 98.945 62.900 99.225 ;
        RECT 57.540 98.895 57.920 98.945 ;
        RECT 62.520 98.895 62.900 98.945 ;
        RECT 89.990 99.225 90.370 99.275 ;
        RECT 94.970 99.225 95.350 99.275 ;
        RECT 89.990 98.945 95.350 99.225 ;
        RECT 89.990 98.895 90.370 98.945 ;
        RECT 94.970 98.895 95.350 98.945 ;
        RECT 122.440 99.225 122.820 99.275 ;
        RECT 127.420 99.225 127.800 99.275 ;
        RECT 122.440 98.945 127.800 99.225 ;
        RECT 122.440 98.895 122.820 98.945 ;
        RECT 127.420 98.895 127.800 98.945 ;
        RECT 154.890 99.225 155.270 99.275 ;
        RECT 159.870 99.225 160.250 99.275 ;
        RECT 154.890 98.945 160.250 99.225 ;
        RECT 162.315 99.070 162.695 99.450 ;
        RECT 164.355 99.070 164.735 99.450 ;
        RECT 166.140 99.070 166.520 99.450 ;
        RECT 154.890 98.895 155.270 98.945 ;
        RECT 159.870 98.895 160.250 98.945 ;
        RECT 25.200 97.570 25.580 97.950 ;
        RECT 29.120 97.570 29.500 97.950 ;
        RECT 31.920 97.615 34.160 97.995 ;
        RECT 64.370 97.615 66.610 97.995 ;
        RECT 96.820 97.615 99.060 97.995 ;
        RECT 129.270 97.615 131.510 97.995 ;
        RECT 58.820 97.385 59.200 97.435 ;
        RECT 62.520 97.385 62.900 97.435 ;
        RECT 58.820 97.105 62.900 97.385 ;
        RECT 58.820 97.055 59.200 97.105 ;
        RECT 62.520 97.055 62.900 97.105 ;
        RECT 91.270 97.385 91.650 97.435 ;
        RECT 94.970 97.385 95.350 97.435 ;
        RECT 91.270 97.105 95.350 97.385 ;
        RECT 91.270 97.055 91.650 97.105 ;
        RECT 94.970 97.055 95.350 97.105 ;
        RECT 123.720 97.385 124.100 97.435 ;
        RECT 127.420 97.385 127.800 97.435 ;
        RECT 123.720 97.105 127.800 97.385 ;
        RECT 123.720 97.055 124.100 97.105 ;
        RECT 127.420 97.055 127.800 97.105 ;
        RECT 156.170 97.385 156.550 97.435 ;
        RECT 159.870 97.385 160.250 97.435 ;
        RECT 156.170 97.105 160.250 97.385 ;
        RECT 156.170 97.055 156.550 97.105 ;
        RECT 159.870 97.055 160.250 97.105 ;
        RECT 31.925 95.730 34.165 96.110 ;
        RECT 64.375 95.730 66.615 96.110 ;
        RECT 96.825 95.730 99.065 96.110 ;
        RECT 129.275 95.730 131.515 96.110 ;
        RECT 162.315 96.070 162.695 96.450 ;
        RECT 164.355 96.070 164.735 96.450 ;
        RECT 166.140 96.070 166.520 96.450 ;
        RECT 31.920 94.970 34.160 95.350 ;
        RECT 64.370 94.970 66.610 95.350 ;
        RECT 96.820 94.970 99.060 95.350 ;
        RECT 129.270 94.970 131.510 95.350 ;
        RECT 25.200 94.570 25.580 94.950 ;
        RECT 29.120 94.570 29.500 94.950 ;
        RECT 60.100 94.740 60.480 94.790 ;
        RECT 62.520 94.740 62.900 94.790 ;
        RECT 60.100 94.460 62.900 94.740 ;
        RECT 60.100 94.410 60.480 94.460 ;
        RECT 62.520 94.410 62.900 94.460 ;
        RECT 92.550 94.740 92.930 94.790 ;
        RECT 94.970 94.740 95.350 94.790 ;
        RECT 92.550 94.460 95.350 94.740 ;
        RECT 92.550 94.410 92.930 94.460 ;
        RECT 94.970 94.410 95.350 94.460 ;
        RECT 125.000 94.740 125.380 94.790 ;
        RECT 127.420 94.740 127.800 94.790 ;
        RECT 125.000 94.460 127.800 94.740 ;
        RECT 125.000 94.410 125.380 94.460 ;
        RECT 127.420 94.410 127.800 94.460 ;
        RECT 157.450 94.740 157.830 94.790 ;
        RECT 159.870 94.740 160.250 94.790 ;
        RECT 157.450 94.460 160.250 94.740 ;
        RECT 157.450 94.410 157.830 94.460 ;
        RECT 159.870 94.410 160.250 94.460 ;
        RECT 31.920 93.130 34.160 93.510 ;
        RECT 64.370 93.130 66.610 93.510 ;
        RECT 96.820 93.130 99.060 93.510 ;
        RECT 129.270 93.130 131.510 93.510 ;
        RECT 162.315 93.070 162.695 93.450 ;
        RECT 164.355 93.070 164.735 93.450 ;
        RECT 166.140 93.070 166.520 93.450 ;
        RECT 61.380 92.900 61.760 92.950 ;
        RECT 62.520 92.900 62.900 92.950 ;
        RECT 61.380 92.620 62.900 92.900 ;
        RECT 61.380 92.570 61.760 92.620 ;
        RECT 62.520 92.570 62.900 92.620 ;
        RECT 93.830 92.900 94.210 92.950 ;
        RECT 94.970 92.900 95.350 92.950 ;
        RECT 93.830 92.620 95.350 92.900 ;
        RECT 93.830 92.570 94.210 92.620 ;
        RECT 94.970 92.570 95.350 92.620 ;
        RECT 126.280 92.900 126.660 92.950 ;
        RECT 127.420 92.900 127.800 92.950 ;
        RECT 126.280 92.620 127.800 92.900 ;
        RECT 126.280 92.570 126.660 92.620 ;
        RECT 127.420 92.570 127.800 92.620 ;
        RECT 158.730 92.900 159.110 92.950 ;
        RECT 159.870 92.900 160.250 92.950 ;
        RECT 158.730 92.620 160.250 92.900 ;
        RECT 158.730 92.570 159.110 92.620 ;
        RECT 159.870 92.570 160.250 92.620 ;
        RECT 25.200 91.570 25.580 91.950 ;
        RECT 29.120 91.570 29.500 91.950 ;
        RECT 31.920 91.290 34.160 91.670 ;
        RECT 64.370 91.290 66.610 91.670 ;
        RECT 96.820 91.290 99.060 91.670 ;
        RECT 129.270 91.290 131.510 91.670 ;
        RECT 62.520 90.730 63.040 91.110 ;
        RECT 94.970 90.730 95.490 91.110 ;
        RECT 127.420 90.730 127.940 91.110 ;
        RECT 159.870 90.730 160.390 91.110 ;
        RECT 162.315 90.070 162.695 90.450 ;
        RECT 164.355 90.070 164.735 90.450 ;
        RECT 166.140 90.070 166.520 90.450 ;
        RECT 25.200 88.570 25.580 88.950 ;
        RECT 29.120 88.570 29.500 88.950 ;
        RECT 25.200 85.570 25.580 85.950 ;
        RECT 162.315 84.070 162.695 84.450 ;
        RECT 164.355 84.070 164.735 84.450 ;
        RECT 166.140 84.070 166.520 84.450 ;
        RECT 25.200 82.570 25.580 82.950 ;
        RECT 29.120 82.570 29.500 82.950 ;
        RECT 62.020 82.165 62.900 82.545 ;
        RECT 94.470 82.165 95.350 82.545 ;
        RECT 126.920 82.165 127.800 82.545 ;
        RECT 159.370 82.165 160.250 82.545 ;
        RECT 31.920 81.605 34.160 81.985 ;
        RECT 64.370 81.605 66.610 81.985 ;
        RECT 96.820 81.605 99.060 81.985 ;
        RECT 129.270 81.605 131.510 81.985 ;
        RECT 162.315 81.070 162.695 81.450 ;
        RECT 164.355 81.070 164.735 81.450 ;
        RECT 166.140 81.070 166.520 81.450 ;
        RECT 60.740 80.655 61.120 80.705 ;
        RECT 62.520 80.655 62.900 80.705 ;
        RECT 60.740 80.375 62.900 80.655 ;
        RECT 60.740 80.325 61.120 80.375 ;
        RECT 62.520 80.325 62.900 80.375 ;
        RECT 93.190 80.655 93.570 80.705 ;
        RECT 94.970 80.655 95.350 80.705 ;
        RECT 93.190 80.375 95.350 80.655 ;
        RECT 93.190 80.325 93.570 80.375 ;
        RECT 94.970 80.325 95.350 80.375 ;
        RECT 125.640 80.655 126.020 80.705 ;
        RECT 127.420 80.655 127.800 80.705 ;
        RECT 125.640 80.375 127.800 80.655 ;
        RECT 125.640 80.325 126.020 80.375 ;
        RECT 127.420 80.325 127.800 80.375 ;
        RECT 158.090 80.655 158.470 80.705 ;
        RECT 159.870 80.655 160.250 80.705 ;
        RECT 158.090 80.375 160.250 80.655 ;
        RECT 158.090 80.325 158.470 80.375 ;
        RECT 159.870 80.325 160.250 80.375 ;
        RECT 25.200 79.570 25.580 79.950 ;
        RECT 29.120 79.570 29.500 79.950 ;
        RECT 31.920 79.765 34.160 80.145 ;
        RECT 64.370 79.765 66.610 80.145 ;
        RECT 96.820 79.765 99.060 80.145 ;
        RECT 129.270 79.765 131.510 80.145 ;
        RECT 59.460 78.810 59.840 78.860 ;
        RECT 62.520 78.810 62.900 78.860 ;
        RECT 59.460 78.530 62.900 78.810 ;
        RECT 59.460 78.480 59.840 78.530 ;
        RECT 62.520 78.480 62.900 78.530 ;
        RECT 91.910 78.810 92.290 78.860 ;
        RECT 94.970 78.810 95.350 78.860 ;
        RECT 91.910 78.530 95.350 78.810 ;
        RECT 91.910 78.480 92.290 78.530 ;
        RECT 94.970 78.480 95.350 78.530 ;
        RECT 124.360 78.810 124.740 78.860 ;
        RECT 127.420 78.810 127.800 78.860 ;
        RECT 124.360 78.530 127.800 78.810 ;
        RECT 124.360 78.480 124.740 78.530 ;
        RECT 127.420 78.480 127.800 78.530 ;
        RECT 156.810 78.810 157.190 78.860 ;
        RECT 159.870 78.810 160.250 78.860 ;
        RECT 156.810 78.530 160.250 78.810 ;
        RECT 156.810 78.480 157.190 78.530 ;
        RECT 159.870 78.480 160.250 78.530 ;
        RECT 31.920 77.920 34.160 78.300 ;
        RECT 64.370 77.920 66.610 78.300 ;
        RECT 96.820 77.920 99.060 78.300 ;
        RECT 129.270 77.920 131.510 78.300 ;
        RECT 162.315 78.070 162.695 78.450 ;
        RECT 164.355 78.070 164.735 78.450 ;
        RECT 166.140 78.070 166.520 78.450 ;
        RECT 31.925 77.160 34.165 77.540 ;
        RECT 64.375 77.160 66.615 77.540 ;
        RECT 96.825 77.160 99.065 77.540 ;
        RECT 129.275 77.160 131.515 77.540 ;
        RECT 25.200 76.570 25.580 76.950 ;
        RECT 29.120 76.570 29.500 76.950 ;
        RECT 58.180 76.170 58.560 76.220 ;
        RECT 62.520 76.170 62.900 76.220 ;
        RECT 58.180 75.890 62.900 76.170 ;
        RECT 58.180 75.840 58.560 75.890 ;
        RECT 62.520 75.840 62.900 75.890 ;
        RECT 90.630 76.170 91.010 76.220 ;
        RECT 94.970 76.170 95.350 76.220 ;
        RECT 90.630 75.890 95.350 76.170 ;
        RECT 90.630 75.840 91.010 75.890 ;
        RECT 94.970 75.840 95.350 75.890 ;
        RECT 123.080 76.170 123.460 76.220 ;
        RECT 127.420 76.170 127.800 76.220 ;
        RECT 123.080 75.890 127.800 76.170 ;
        RECT 123.080 75.840 123.460 75.890 ;
        RECT 127.420 75.840 127.800 75.890 ;
        RECT 155.530 76.170 155.910 76.220 ;
        RECT 159.870 76.170 160.250 76.220 ;
        RECT 155.530 75.890 160.250 76.170 ;
        RECT 155.530 75.840 155.910 75.890 ;
        RECT 159.870 75.840 160.250 75.890 ;
        RECT 31.920 75.280 34.160 75.660 ;
        RECT 64.370 75.280 66.610 75.660 ;
        RECT 96.820 75.280 99.060 75.660 ;
        RECT 129.270 75.280 131.510 75.660 ;
        RECT 162.315 75.070 162.695 75.450 ;
        RECT 164.355 75.070 164.735 75.450 ;
        RECT 166.140 75.070 166.520 75.450 ;
        RECT 56.900 74.330 57.280 74.380 ;
        RECT 62.520 74.330 62.900 74.380 ;
        RECT 56.900 74.050 62.900 74.330 ;
        RECT 56.900 74.000 57.280 74.050 ;
        RECT 62.520 74.000 62.900 74.050 ;
        RECT 89.350 74.330 89.730 74.380 ;
        RECT 94.970 74.330 95.350 74.380 ;
        RECT 89.350 74.050 95.350 74.330 ;
        RECT 89.350 74.000 89.730 74.050 ;
        RECT 94.970 74.000 95.350 74.050 ;
        RECT 121.800 74.330 122.180 74.380 ;
        RECT 127.420 74.330 127.800 74.380 ;
        RECT 121.800 74.050 127.800 74.330 ;
        RECT 121.800 74.000 122.180 74.050 ;
        RECT 127.420 74.000 127.800 74.050 ;
        RECT 154.250 74.330 154.630 74.380 ;
        RECT 159.870 74.330 160.250 74.380 ;
        RECT 154.250 74.050 160.250 74.330 ;
        RECT 154.250 74.000 154.630 74.050 ;
        RECT 159.870 74.000 160.250 74.050 ;
        RECT 25.200 73.570 25.580 73.950 ;
        RECT 29.120 73.570 29.500 73.950 ;
        RECT 31.920 73.440 34.160 73.820 ;
        RECT 64.370 73.440 66.610 73.820 ;
        RECT 96.820 73.440 99.060 73.820 ;
        RECT 129.270 73.440 131.510 73.820 ;
        RECT 55.620 72.485 56.000 72.535 ;
        RECT 62.520 72.485 62.900 72.535 ;
        RECT 55.620 72.205 62.900 72.485 ;
        RECT 55.620 72.155 56.000 72.205 ;
        RECT 62.520 72.155 62.900 72.205 ;
        RECT 88.070 72.485 88.450 72.535 ;
        RECT 94.970 72.485 95.350 72.535 ;
        RECT 88.070 72.205 95.350 72.485 ;
        RECT 88.070 72.155 88.450 72.205 ;
        RECT 94.970 72.155 95.350 72.205 ;
        RECT 120.520 72.485 120.900 72.535 ;
        RECT 127.420 72.485 127.800 72.535 ;
        RECT 120.520 72.205 127.800 72.485 ;
        RECT 120.520 72.155 120.900 72.205 ;
        RECT 127.420 72.155 127.800 72.205 ;
        RECT 152.970 72.485 153.350 72.535 ;
        RECT 159.870 72.485 160.250 72.535 ;
        RECT 152.970 72.205 160.250 72.485 ;
        RECT 152.970 72.155 153.350 72.205 ;
        RECT 159.870 72.155 160.250 72.205 ;
        RECT 162.315 72.070 162.695 72.450 ;
        RECT 164.355 72.070 164.735 72.450 ;
        RECT 166.140 72.070 166.520 72.450 ;
        RECT 31.920 71.595 34.160 71.975 ;
        RECT 64.370 71.595 66.610 71.975 ;
        RECT 96.820 71.595 99.060 71.975 ;
        RECT 129.270 71.595 131.510 71.975 ;
        RECT 25.200 70.570 25.580 70.950 ;
        RECT 29.120 70.570 29.500 70.950 ;
        RECT 31.925 70.835 34.165 71.215 ;
        RECT 64.375 70.835 66.615 71.215 ;
        RECT 96.825 70.835 99.065 71.215 ;
        RECT 129.275 70.835 131.515 71.215 ;
        RECT 54.340 69.845 54.720 69.895 ;
        RECT 62.520 69.845 62.900 69.895 ;
        RECT 54.340 69.565 62.900 69.845 ;
        RECT 54.340 69.515 54.720 69.565 ;
        RECT 62.520 69.515 62.900 69.565 ;
        RECT 86.790 69.845 87.170 69.895 ;
        RECT 94.970 69.845 95.350 69.895 ;
        RECT 86.790 69.565 95.350 69.845 ;
        RECT 86.790 69.515 87.170 69.565 ;
        RECT 94.970 69.515 95.350 69.565 ;
        RECT 119.240 69.845 119.620 69.895 ;
        RECT 127.420 69.845 127.800 69.895 ;
        RECT 119.240 69.565 127.800 69.845 ;
        RECT 119.240 69.515 119.620 69.565 ;
        RECT 127.420 69.515 127.800 69.565 ;
        RECT 151.690 69.845 152.070 69.895 ;
        RECT 159.870 69.845 160.250 69.895 ;
        RECT 151.690 69.565 160.250 69.845 ;
        RECT 151.690 69.515 152.070 69.565 ;
        RECT 159.870 69.515 160.250 69.565 ;
        RECT 31.920 68.955 34.160 69.335 ;
        RECT 64.370 68.955 66.610 69.335 ;
        RECT 96.820 68.955 99.060 69.335 ;
        RECT 129.270 68.955 131.510 69.335 ;
        RECT 162.315 69.070 162.695 69.450 ;
        RECT 164.355 69.070 164.735 69.450 ;
        RECT 166.140 69.070 166.520 69.450 ;
        RECT 53.060 68.005 53.440 68.055 ;
        RECT 62.520 68.005 62.900 68.055 ;
        RECT 25.200 67.570 25.580 67.950 ;
        RECT 29.120 67.570 29.500 67.950 ;
        RECT 53.060 67.725 62.900 68.005 ;
        RECT 53.060 67.675 53.440 67.725 ;
        RECT 62.520 67.675 62.900 67.725 ;
        RECT 85.510 68.005 85.890 68.055 ;
        RECT 94.970 68.005 95.350 68.055 ;
        RECT 85.510 67.725 95.350 68.005 ;
        RECT 85.510 67.675 85.890 67.725 ;
        RECT 94.970 67.675 95.350 67.725 ;
        RECT 117.960 68.005 118.340 68.055 ;
        RECT 127.420 68.005 127.800 68.055 ;
        RECT 117.960 67.725 127.800 68.005 ;
        RECT 117.960 67.675 118.340 67.725 ;
        RECT 127.420 67.675 127.800 67.725 ;
        RECT 150.410 68.005 150.790 68.055 ;
        RECT 159.870 68.005 160.250 68.055 ;
        RECT 150.410 67.725 160.250 68.005 ;
        RECT 150.410 67.675 150.790 67.725 ;
        RECT 159.870 67.675 160.250 67.725 ;
        RECT 31.920 67.115 34.160 67.495 ;
        RECT 64.370 67.115 66.610 67.495 ;
        RECT 96.820 67.115 99.060 67.495 ;
        RECT 129.270 67.115 131.510 67.495 ;
  END
END efuse_array_64x8
END LIBRARY

