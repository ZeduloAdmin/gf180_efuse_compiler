* NGSPICE file created from efuse_array_64x8.ext - technology: gf180mcuD

.subckt efuse_array_64x8 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3]
+ BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11]
+ BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18]
+ BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25]
+ BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32]
+ BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39]
+ BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46]
+ BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53]
+ BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60]
+ BIT_SEL[61] BIT_SEL[62] BIT_SEL[63] COL_PROG_N[0] OUT[0] COL_PROG_N[1] OUT[1] COL_PROG_N[2]
+ OUT[2] COL_PROG_N[3] OUT[3] COL_PROG_N[4] OUT[4] COL_PROG_N[5] OUT[5] COL_PROG_N[6]
+ OUT[6] COL_PROG_N[7] OUT[7]
X0 a_1340_61431.t1 a_638_58903.t29 efuse
X1 a_7830_61063.t1 a_638_58903.t0 efuse
X2 VSS.t28 BIT_SEL[50].t0 a_20810_20781.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X3 a_20810_3154.t0 BIT_SEL[49].t0 VSS.t426 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X4 a_638_27395.t36 a_1340_25152.t1 efuse
X5 VDD a_110_52624.t1 a_154_52536.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X6 a_638_35272.t13 a_1340_32660.t0 efuse
X7 a_14320_41274.t0 BIT_SEL[39].t0 VSS.t409 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X8 a_638_43149.t5 a_1340_40906.t0 efuse
X9 a_7738_27712.t1 a_638_27395.t52 efuse
X10 a_1340_9029.t1 BIT_SEL[11].t0 VSS.t415 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X11 a_638_11641.t66 a_20810_9398.t1 efuse
X12 a_110_29441.t0 a_154_29353.t1 VSS.t312 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X13 a_7830_25152.t0 BIT_SEL[25].t0 VSS.t278 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X14 VDD a_110_6258.t1 a_154_6170.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 VDD a_110_61397.t1 a_154_61309.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X16 VDD a_110_49568.t2 OUT[6].t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X17 a_7738_43466.t1 a_638_43149.t59 efuse
X18 VSS.t505 BIT_SEL[52].t0 a_20810_36903.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X19 a_638_11641.t29 a_1340_11031.t1 efuse
X20 a_110_16188.t0 a_154_16100.t1 VSS.t424 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X21 VSS.t27 BIT_SEL[50].t1 a_20810_52289.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X22 VSS.t573 BIT_SEL[38].t0 a_14320_13801.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X23 a_638_27395.t1 a_20810_25152.t0 efuse
X24 a_7830_25520.t0 BIT_SEL[23].t0 VSS.t439 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X25 a_20810_7557.t1 a_638_3764.t57 efuse
X26 VDD a_110_434.t1 a_154_346.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X27 a_14320_62328.t1 a_638_58903.t61 efuse
X28 VSS.t357 BIT_SEL[54].t0 a_20810_37432.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X29 VSS.t458 a_110_34710.t6 a_110_33814.t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X30 VSS.t352 BIT_SEL[52].t1 a_20810_52657.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X31 a_1248_59220.t1 a_638_58903.t18 efuse
X32 a_638_27395.t9 a_1340_26785.t1 efuse
X33 a_1340_7557.t0 a_638_3764.t28 efuse
X34 a_638_43149.t17 a_20810_40906.t0 efuse
X35 a_20810_40906.t1 BIT_SEL[57].t0 VSS.t372 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X36 VSS.t381 BIT_SEL[60].t0 a_20810_7189.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X37 a_638_58903.t32 a_20810_55763.t1 efuse
X38 VSS.t320 BIT_SEL[58].t0 a_20810_38168.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X39 a_110_24961.t0 a_154_24873.t1 VSS.t485 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X40 VDD a_110_21116.t1 a_154_21028.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X41 a_1340_1889.t0 BIT_SEL[7].t0 VSS.t517 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X42 a_20810_26417.t0 BIT_SEL[51].t0 VSS.t579 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X43 VSS.t394 a_110_2306.t2 OUT[0].t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X44 VSS.t612 BIT_SEL[38].t1 a_14320_45309.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X45 a_638_43149.t4 a_1340_42539.t0 efuse
X46 VSS.t174 BIT_SEL[62].t0 a_20810_7557.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X47 VDD a_110_10183.t2 a_110_11079.t3 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X48 a_1340_57028.t1 BIT_SEL[7].t1 VSS.t518 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X49 a_638_11641.t2 a_14320_9398.t0 efuse
X50 a_110_40715.t0 a_154_40627.t1 VSS.t464 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X51 VSS.t491 BIT_SEL[14].t0 a_1340_23311.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X52 a_110_5810.t0 a_154_5722.t1 VSS.t69 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X53 a_7830_52657.t1 a_638_51026.t15 efuse
X54 a_20810_26785.t1 BIT_SEL[49].t1 VSS.t152 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X55 a_638_3764.t56 a_14320_1521.t1 efuse
X56 a_638_58903.t13 a_1340_55395.t0 efuse
X57 VSS.t49 BIT_SEL[40].t0 a_14320_45677.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X58 VSS.t80 BIT_SEL[48].t0 a_20718_19835.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X59 a_638_3764.t7 COL_PROG_N[0].t0 VDD.t77 VDD.t76 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X60 a_110_62741.t0 a_154_62653.t1 VSS.t332 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X61 a_1340_23887.t0 BIT_SEL[15].t0 VSS.t242 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X62 a_20810_42539.t1 BIT_SEL[49].t2 VSS.t404 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X63 a_638_27395.t66 a_14320_25152.t1 efuse
X64 a_7830_14169.t0 a_638_11641.t5 efuse
X65 VSS.t50 BIT_SEL[40].t1 a_14320_61431.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X66 VSS.t213 BIT_SEL[22].t0 a_7830_29555.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X67 VSS.t59 BIT_SEL[20].t0 a_7830_44780.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X68 VSS.t353 BIT_SEL[52].t2 a_20810_21149.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X69 a_638_58903.t4 a_20810_57556.t0 efuse
X70 a_14228_4081.t0 a_638_3764.t0 efuse
X71 a_638_58903.t36 a_20810_58293.t1 efuse
X72 a_638_43149.t29 a_14320_40906.t1 efuse
X73 VDD a_110_37318.t1 a_154_37230.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X74 VSS.t116 BIT_SEL[34].t0 a_14320_12904.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X75 a_20810_58293.t0 BIT_SEL[49].t3 VSS.t277 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X76 a_7830_29923.t0 a_638_27395.t2 efuse
X77 a_110_36198.t0 a_154_36110.t1 VSS.t523 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X78 VDD a_110_26833.t6 a_110_25937.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X79 a_1340_55395.t1 BIT_SEL[15].t1 VSS.t243 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X80 VDD a_110_32390.t1 a_154_32302.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X81 a_638_19518.t10 a_7830_16010.t0 efuse
X82 a_7830_45677.t0 a_638_43149.t18 efuse
X83 a_7830_18908.t0 BIT_SEL[17].t0 VSS.t260 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X84 VSS.t335 BIT_SEL[56].t0 a_20810_6292.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X85 a_110_8759.t0 a_154_8671.t1 VSS.t265 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X86 a_638_58903.t1 a_1340_57028.t0 efuse
X87 VSS.t51 BIT_SEL[40].t2 a_14320_14169.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X88 a_1340_55763.t0 BIT_SEL[13].t0 VSS.t345 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X89 VSS.t266 BIT_SEL[16].t0 a_7738_11958.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X90 a_638_35272.t7 a_7830_31764.t0 efuse
X91 a_110_31233.t0 a_154_31145.t1 VSS.t32 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X92 a_14320_20781.t0 a_638_19518.t21 efuse
X93 a_1340_33925.t0 BIT_SEL[5].t0 VSS.t70 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X94 VDD a_110_32838.t1 a_154_32750.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X95 VSS.t532 BIT_SEL[42].t0 a_14320_14537.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X96 VDD a_110_58341.t6 a_110_57445.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X97 a_1340_1521.t0 BIT_SEL[9].t0 VSS.t85 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X98 a_14320_36535.t0 a_638_35272.t8 efuse
X99 a_20810_41274.t0 BIT_SEL[55].t0 VSS.t593 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X100 VSS.t486 BIT_SEL[32].t0 a_14228_4081.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X101 a_1340_13272.t1 a_638_11641.t23 efuse
X102 VSS.t117 BIT_SEL[34].t1 a_14320_60166.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X103 VDD a_110_54864.t1 a_154_54776.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X104 a_638_58903.t31 a_14320_58293.t0 efuse
X105 VDD PRESET_N.t0 a_110_34710.t1 VDD pfet_06v0 ad=0.3172p pd=1.74u as=0.4575p ps=1.97u w=1.22u l=0.5u
X106 VSS.t229 BIT_SEL[12].t0 a_1340_22943.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X107 VDD a_110_48592.t1 a_154_48504.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X108 a_20810_8133.t0 BIT_SEL[63].t0 VSS.t225 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X109 a_638_19518.t5 a_7830_17643.t0 efuse
X110 VSS.t476 BIT_SEL[36].t0 a_14320_60534.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X111 VSS.t267 BIT_SEL[16].t1 a_7738_43466.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X112 VSS.t358 BIT_SEL[54].t1 a_20810_13801.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X113 a_638_3764.t9 a_1340_1889.t1 efuse
X114 VSS.t533 BIT_SEL[42].t1 a_14320_46045.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X115 a_1340_29026.t0 a_638_27395.t4 efuse
X116 VDD a_110_9207.t1 a_154_9119.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X117 VSS.t479 BIT_SEL[18].t0 a_7830_44412.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X118 a_20810_62328.t1 a_638_58903.t14 efuse
X119 a_638_35272.t17 a_7830_33397.t0 efuse
X120 a_1340_24255.t0 BIT_SEL[13].t1 VSS.t346 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X121 VSS.t6 BIT_SEL[0].t0 a_1248_59220.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X122 a_14320_34294.t1 BIT_SEL[35].t0 VSS.t451 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X123 a_7830_6660.t0 a_638_3764.t11 efuse
X124 a_638_58903.t30 SENSE.t0 a_110_58341.t3 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X125 a_1340_44780.t0 a_638_43149.t10 efuse
X126 VSS.t240 a_110_33814.t2 OUT[4].t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X127 a_110_1330.t0 a_154_1242.t1 VSS.t319 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X128 a_14320_34662.t1 BIT_SEL[33].t0 VSS.t585 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X129 a_7830_33397.t1 BIT_SEL[23].t1 VSS.t600 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X130 a_1340_32660.t1 BIT_SEL[11].t1 VSS.t414 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X131 a_14320_53554.t0 a_638_51026.t16 efuse
X132 VDD a_110_23356.t1 a_154_23268.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X133 VSS.t477 BIT_SEL[36].t1 a_14320_13272.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X134 VSS.t359 BIT_SEL[54].t2 a_20810_45309.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X135 VSS.t239 a_110_42587.t6 a_110_41691.t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X136 a_1340_18171.t0 BIT_SEL[5].t1 VSS.t71 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X137 a_7830_18540.t0 BIT_SEL[19].t0 VSS.t407 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X138 a_638_19518.t7 a_14320_16378.t0 efuse
X139 VDD a_110_17084.t1 a_154_16996.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X140 VSS.t336 BIT_SEL[56].t1 a_20810_45677.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X141 a_7830_41802.t0 BIT_SEL[21].t0 VSS.t440 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X142 a_20810_61431.t0 a_638_58903.t62 efuse
X143 a_638_35272.t66 a_14320_32132.t1 efuse
X144 VSS.t14 BIT_SEL[10].t0 a_1340_6660.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X145 a_20810_60534.t0 a_638_58903.t3 efuse
X146 a_110_61845.t0 a_154_61757.t1 VSS.t204 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X147 VSS.t337 BIT_SEL[56].t2 a_20810_61431.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X148 a_638_11641.t0 a_1340_9029.t0 efuse
X149 a_638_51026.t67 a_7830_47886.t1 efuse
X150 VSS.t7 BIT_SEL[0].t1 a_1248_27712.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X151 a_638_27395.t23 SENSE.t1 a_110_26833.t4 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X152 a_110_55573.t0 a_154_55485.t1 VSS.t510 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X153 a_638_51026.t6 a_7830_48783.t0 efuse
X154 a_1340_50048.t1 BIT_SEL[3].t0 VSS.t183 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X155 a_638_35272.t2 COL_PROG_N[4].t0 VDD.t3 VDD.t2 pfet_06v0 ad=16.83p pd=77.38u as=9.945p ps=38.77u w=38.25u l=0.5u
X156 VSS.t26 BIT_SEL[50].t2 a_20810_12904.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X157 VSS.t191 BIT_SEL[2].t0 a_1340_28658.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X158 a_7830_23311.t1 a_638_19518.t17 efuse
X159 a_1340_61799.t1 a_638_58903.t24 efuse
X160 a_14228_51343.t1 a_638_51026.t33 efuse
X161 a_638_43149.t30 SENSE.t2 a_110_42587.t5 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X162 VSS.t110 BIT_SEL[44].t0 a_14320_38697.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X163 VSS.t114 BIT_SEL[34].t2 a_14320_5027.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X164 a_638_35272.t58 COL_PROG_N[4].t1 VDD.t208 VDD.t76 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X165 a_638_27395.t55 a_1340_24783.t1 efuse
X166 VDD a_110_25937.t2 OUT[3].t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X167 a_20810_5924.t0 a_638_3764.t1 efuse
X168 VSS.t58 a_110_11079.t6 a_110_10183.t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X169 a_638_19518.t4 a_14320_18171.t0 efuse
X170 VSS.t172 a_110_18060.t2 OUT[2].t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X171 a_7830_39065.t0 a_638_35272.t0 efuse
X172 VSS.t111 BIT_SEL[44].t1 a_14320_54451.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X173 VSS.t208 BIT_SEL[24].t0 a_7830_37800.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X174 a_110_14583.t0 a_154_14495.t1 VSS.t171 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X175 a_638_43149.t50 a_1340_40537.t1 efuse
X176 a_1340_5924.t0 a_638_3764.t19 efuse
X177 a_7830_10294.t0 BIT_SEL[21].t1 VSS.t441 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X178 VSS.t338 BIT_SEL[56].t3 a_20810_14169.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X179 VDD a_110_60501.t1 a_154_60413.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X180 a_14320_40009.t0 BIT_SEL[45].t0 VSS.t604 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X181 a_638_35272.t42 a_14320_33925.t0 efuse
X182 VSS.t498 BIT_SEL[46].t0 a_14320_54819.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X183 a_110_30337.t0 a_154_30249.t1 VSS.t203 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X184 VDD a_110_28321.t1 a_154_28233.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X185 VDD.t111 COL_PROG_N[0].t1 a_638_3764.t29 VDD.t86 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X186 VSS.t321 BIT_SEL[58].t1 a_20810_14537.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X187 VSS.t490 BIT_SEL[14].t1 a_1340_62696.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X188 a_14320_60534.t1 a_638_58903.t68 efuse
X189 a_1340_33029.t0 BIT_SEL[9].t1 VSS.t86 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X190 a_638_3764.t10 a_1340_624.t0 efuse
X191 VSS.t173 a_110_18060.t3 a_110_18956.t4 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X192 a_7830_60166.t0 a_638_58903.t45 efuse
X193 VSS.t495 BIT_SEL[4].t0 a_1340_5395.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X194 a_638_51026.t3 a_1340_50048.t0 efuse
X195 a_110_24065.t0 a_154_23977.t1 VSS.t530 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X196 a_638_3764.t33 SENSE.t3 a_110_3202.t5 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X197 a_14320_2417.t0 BIT_SEL[37].t0 VSS.t552 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X198 VDD a_110_57445.t2 OUT[7].t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X199 VSS.t613 BIT_SEL[38].t2 a_14320_21678.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X200 a_7830_22414.t0 a_638_19518.t0 efuse
X201 VSS.t25 BIT_SEL[50].t3 a_20810_60166.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X202 a_1340_22046.t0 a_638_19518.t15 efuse
X203 a_7830_21678.t0 a_638_19518.t1 efuse
X204 VDD a_110_53968.t1 a_154_53880.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X205 VSS.t347 BIT_SEL[6].t0 a_1340_5924.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X206 a_110_46091.t0 a_154_46003.t1 VSS.t514 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X207 a_7830_5027.t0 a_638_3764.t35 efuse
X208 VSS.t354 BIT_SEL[52].t3 a_20810_60534.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X209 a_638_58903.t58 a_20810_55395.t1 efuse
X210 a_1340_48783.t0 BIT_SEL[9].t2 VSS.t87 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X211 a_7830_38168.t0 a_638_35272.t1 efuse
X212 a_110_18956.t2 PRESET_N.t1 VDD VDD pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X213 a_638_58903.t5 a_20810_56291.t0 efuse
X214 VDD a_110_47696.t1 a_154_47608.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X215 a_7830_37432.t0 a_638_35272.t6 efuse
X216 VSS.t480 BIT_SEL[18].t1 a_7830_20781.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X217 a_1340_37800.t1 a_638_35272.t60 efuse
X218 VSS.t322 BIT_SEL[58].t2 a_20810_46045.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X219 a_7830_9398.t1 BIT_SEL[25].t1 VSS.t279 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X220 a_14320_49679.t0 BIT_SEL[37].t1 VSS.t553 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X221 a_638_51026.t54 a_20810_50048.t1 efuse
X222 VDD PRESET_N.t2 a_110_42587.t2 VDD pfet_06v0 ad=0.3172p pd=1.74u as=0.4575p ps=1.97u w=1.22u l=0.5u
X223 a_20810_34294.t0 BIT_SEL[51].t1 VSS.t580 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X224 a_110_46539.t0 a_154_46451.t1 VSS.t598 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X225 VSS.t610 BIT_SEL[38].t3 a_14320_53186.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X226 a_7830_9766.t1 BIT_SEL[23].t2 VSS.t599 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X227 a_638_51026.t2 a_14320_49151.t0 efuse
X228 VSS.t468 BIT_SEL[14].t2 a_1340_31188.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X229 a_1340_16010.t0 BIT_SEL[15].t2 VSS.t244 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X230 a_20810_34662.t1 BIT_SEL[49].t4 VSS.t275 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X231 VSS.t52 BIT_SEL[40].t3 a_14320_53554.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X232 a_14320_22943.t1 a_638_19518.t68 efuse
X233 a_110_12567.t0 a_154_12479.t1 VSS.t567 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X234 VSS.t481 BIT_SEL[18].t2 a_7830_52289.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X235 VSS.t60 BIT_SEL[20].t1 a_7830_36903.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X236 a_1248_19835.t1 a_638_19518.t66 efuse
X237 VSS.t355 BIT_SEL[52].t4 a_20810_13272.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X238 a_14320_16906.t0 BIT_SEL[43].t0 VSS.t574 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X239 a_1340_31764.t0 BIT_SEL[15].t3 VSS.t245 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X240 VSS.t496 BIT_SEL[4].t1 a_1340_29026.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X241 VSS.t499 BIT_SEL[46].t1 a_14320_39065.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X242 VSS.t214 BIT_SEL[22].t1 a_7830_37432.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X243 VDD a_110_29441.t1 a_154_29353.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X244 a_638_19518.t49 a_20810_16378.t1 efuse
X245 VSS.t61 BIT_SEL[20].t2 a_7830_52657.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X246 a_14320_38697.t1 a_638_35272.t39 efuse
X247 a_110_11079.t0 PRESET_N.t3 VDD VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X248 a_1340_17275.t0 BIT_SEL[9].t3 VSS.t88 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X249 a_1248_35589.t1 a_638_35272.t68 efuse
X250 a_638_11641.t57 a_7830_8133.t1 efuse
X251 VDD a_110_16188.t1 a_154_16100.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X252 a_638_58903.t21 a_14320_56291.t1 efuse
X253 a_14320_39641.t0 BIT_SEL[47].t0 VSS.t614 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X254 a_7830_54451.t1 a_638_51026.t7 efuse
X255 a_7830_40906.t1 BIT_SEL[25].t2 VSS.t280 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X256 VSS.t129 BIT_SEL[26].t0 a_7830_38168.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X257 a_638_35272.t10 a_20810_32132.t0 efuse
X258 a_1340_17643.t0 BIT_SEL[7].t2 VSS.t519 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X259 a_20810_7189.t0 a_638_3764.t4 efuse
X260 VDD a_110_34710.t7 a_110_33814.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X261 a_7830_26417.t0 BIT_SEL[19].t1 VSS.t408 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X262 a_110_60949.t0 a_154_60861.t1 VSS.t161 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X263 a_638_51026.t0 a_14320_50048.t0 efuse
X264 a_110_44075.t0 a_154_43987.t1 VSS.t566 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X265 a_638_19518.t48 a_1340_16010.t1 efuse
X266 a_14320_12904.t0 a_638_11641.t3 efuse
X267 a_14320_48414.t0 BIT_SEL[43].t1 VSS.t575 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X268 a_638_27395.t11 a_7830_23887.t0 efuse
X269 a_7830_26785.t1 BIT_SEL[17].t1 VSS.t261 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X270 a_20718_51343.t0 a_638_51026.t23 efuse
X271 a_110_42587.t1 PRESET_N.t4 VDD VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X272 VSS.t382 BIT_SEL[60].t1 a_20810_38697.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X273 VDD a_110_24961.t1 a_154_24873.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X274 VSS.t53 BIT_SEL[40].t4 a_14320_22046.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X275 a_7830_8501.t0 BIT_SEL[29].t0 VSS.t307 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X276 a_638_35272.t35 a_1340_31764.t1 efuse
X277 VSS.t268 BIT_SEL[16].t2 a_7738_19835.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X278 a_638_43149.t11 a_7830_39641.t0 efuse
X279 a_14320_28658.t0 a_638_27395.t10 efuse
X280 a_7830_5395.t1 a_638_3764.t26 efuse
X281 a_1340_62696.t1 a_638_58903.t16 efuse
X282 a_7830_42539.t1 BIT_SEL[17].t2 VSS.t262 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X283 a_638_19518.t3 a_20810_18908.t0 efuse
X284 a_638_19518.t2 a_20810_18171.t0 efuse
X285 a_1340_49151.t0 BIT_SEL[7].t3 VSS.t118 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X286 VDD a_110_40715.t1 a_154_40627.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X287 VSS.t534 BIT_SEL[42].t2 a_14320_22414.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X288 VSS.t383 BIT_SEL[60].t2 a_20810_54451.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X289 VSS.t62 BIT_SEL[20].t3 a_7830_21149.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X290 a_14320_9029.t0 BIT_SEL[43].t2 VSS.t576 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X291 a_14320_44412.t0 a_638_43149.t61 efuse
X292 a_638_3764.t6 COL_PROG_N[0].t2 VDD.t75 VDD.t2 pfet_06v0 ad=16.83p pd=77.38u as=9.945p ps=38.77u w=38.25u l=0.5u
X293 a_638_11641.t28 a_7830_9766.t0 efuse
X294 a_638_58903.t15 a_7830_57556.t1 efuse
X295 a_638_35272.t27 a_20810_33925.t0 efuse
X296 a_638_3764.t13 a_1340_2786.t0 efuse
X297 a_110_4690.t0 a_154_4602.t1 VSS.t33 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X298 a_14320_10663.t1 BIT_SEL[35].t1 VSS.t452 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X299 a_110_13687.t0 a_154_13599.t1 VSS.t572 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X300 VDD a_110_62741.t1 a_154_62653.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X301 a_638_58903.t17 a_7830_58293.t0 efuse
X302 a_1340_52289.t0 a_638_51026.t1 efuse
X303 a_20810_40009.t0 BIT_SEL[61].t0 VSS.t303 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X304 a_638_35272.t9 a_20810_34662.t0 efuse
X305 VDD a_110_7602.t1 a_154_7514.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X306 VSS.t175 BIT_SEL[62].t1 a_20810_54819.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X307 a_7830_58293.t1 BIT_SEL[17].t3 VSS.t263 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X308 a_638_19518.t8 a_1340_17643.t1 efuse
X309 a_14320_11031.t1 BIT_SEL[33].t1 VSS.t586 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X310 a_638_51026.t31 SENSE.t4 a_110_50464.t5 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X311 a_638_27395.t67 a_7830_25520.t1 efuse
X312 VSS.t313 BIT_SEL[54].t3 a_20810_21678.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X313 a_638_3764.t17 a_7830_1521.t0 efuse
X314 a_638_51026.t26 a_14320_47518.t0 efuse
X315 a_14320_7557.t0 a_638_3764.t2 efuse
X316 VSS.t535 BIT_SEL[42].t3 a_14320_53922.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X317 a_638_35272.t18 a_1340_33397.t1 efuse
X318 VDD a_110_2306.t3 a_110_3202.t3 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X319 a_638_43149.t3 a_7830_41274.t0 efuse
X320 VDD a_110_36198.t1 a_154_36110.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X321 a_1340_32132.t0 BIT_SEL[13].t2 VSS.t249 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X322 a_110_45195.t0 a_154_45107.t1 VSS.t360 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X323 a_14320_42171.t0 BIT_SEL[35].t2 VSS.t453 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X324 a_1340_61063.t1 a_638_58903.t59 efuse
X325 a_14320_1889.t0 BIT_SEL[39].t1 VSS.t423 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X326 a_110_7154.t0 a_154_7066.t1 VSS.t283 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X327 a_638_11641.t54 a_14320_8501.t1 efuse
X328 a_14320_53922.t0 a_638_51026.t4 efuse
X329 a_20810_49679.t0 BIT_SEL[53].t0 VSS.t288 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X330 a_110_29889.t0 a_154_29801.t1 VSS.t565 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X331 a_638_19518.t67 a_14320_18908.t1 efuse
X332 a_7830_41274.t1 BIT_SEL[23].t3 VSS.t164 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X333 VSS.t314 BIT_SEL[54].t4 a_20810_53186.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X334 VSS.t301 a_110_50464.t6 a_110_49568.t0 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X335 a_110_31942.t0 a_154_31854.t1 VSS.t539 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X336 VDD a_110_31233.t1 a_154_31145.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X337 a_638_51026.t57 a_20810_49151.t1 efuse
X338 a_638_35272.t22 a_14320_34662.t0 efuse
X339 a_110_882.t0 a_154_794.t1 VSS.t181 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X340 a_638_27395.t3 a_14320_24255.t1 efuse
X341 a_7830_1152.t0 BIT_SEL[27].t0 VSS.t547 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X342 VSS.t339 BIT_SEL[56].t4 a_20810_53554.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X343 VSS.t215 BIT_SEL[22].t2 a_7830_13801.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X344 a_20810_22943.t1 a_638_19518.t12 efuse
X345 a_20810_16906.t0 BIT_SEL[59].t0 VSS.t559 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X346 a_638_43149.t48 a_14320_40009.t1 efuse
X347 VSS.t176 BIT_SEL[62].t2 a_20810_39065.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X348 a_7830_15434.t1 a_638_11641.t14 efuse
X349 a_638_51026.t20 a_1340_47886.t0 efuse
X350 a_638_51026.t66 a_7830_48414.t1 efuse
X351 a_20810_38697.t1 a_638_35272.t12 efuse
X352 VSS.t112 BIT_SEL[44].t2 a_14320_30820.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X353 a_1340_2786.t1 BIT_SEL[3].t1 VSS.t184 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X354 a_20810_39641.t0 BIT_SEL[63].t1 VSS.t226 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X355 VSS.t8 BIT_SEL[0].t2 a_1248_35589.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X356 a_638_35272.t32 SENSE.t5 a_110_34710.t5 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X357 a_638_11641.t11 a_14320_10294.t0 efuse
X358 a_1340_57925.t1 BIT_SEL[3].t2 VSS.t185 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X359 a_638_3764.t12 a_1340_2417.t1 efuse
X360 VSS.t192 BIT_SEL[2].t1 a_1340_36535.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X361 a_7830_31188.t1 a_638_27395.t30 efuse
X362 VSS.t9 BIT_SEL[0].t3 a_1248_51343.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X363 VSS.t113 BIT_SEL[44].t3 a_14320_46574.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X364 a_20810_9398.t0 BIT_SEL[57].t1 VSS.t373 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X365 VSS.t536 BIT_SEL[42].t4 a_14320_61799.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X366 VSS.t216 BIT_SEL[22].t3 a_7830_45309.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X367 a_110_58341.t1 PRESET_N.t5 VDD VDD pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X368 a_20810_48414.t0 BIT_SEL[59].t1 VSS.t560 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X369 VDD a_110_33814.t3 OUT[4].t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X370 a_7830_46942.t1 a_638_43149.t15 efuse
X371 a_638_27395.t0 a_14320_26048.t0 efuse
X372 a_20810_9766.t0 BIT_SEL[55].t1 VSS.t594 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X373 a_20810_22046.t0 a_638_19518.t38 efuse
X374 a_14320_47518.t1 BIT_SEL[47].t1 VSS.t615 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X375 a_110_22460.t0 a_154_22372.t1 VSS.t430 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X376 a_20810_21149.t1 a_638_19518.t65 efuse
X377 VSS.t148 BIT_SEL[44].t4 a_14320_62328.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X378 VSS.t209 BIT_SEL[24].t1 a_7830_45677.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X379 VSS.t340 BIT_SEL[56].t5 a_20810_22046.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X380 a_638_3764.t66 a_7830_1152.t1 efuse
X381 a_14320_1521.t0 BIT_SEL[41].t0 VSS.t205 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X382 a_7830_14537.t0 a_638_11641.t4 efuse
X383 a_14320_47886.t0 BIT_SEL[45].t1 VSS.t605 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X384 a_638_43149.t8 a_14320_41802.t0 efuse
X385 VDD a_110_42587.t7 a_110_41691.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X386 a_7830_13801.t0 a_638_11641.t9 efuse
X387 a_1340_14169.t1 a_638_11641.t65 efuse
X388 a_7830_60534.t1 a_638_58903.t11 efuse
X389 a_638_51026.t5 a_1340_49679.t0 efuse
X390 a_20810_36903.t0 a_638_35272.t5 efuse
X391 a_20810_37800.t0 a_638_35272.t57 efuse
X392 VSS.t210 BIT_SEL[24].t2 a_7830_61431.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X393 a_14320_26048.t1 BIT_SEL[37].t2 VSS.t554 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X394 VSS.t323 BIT_SEL[58].t3 a_20810_22414.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X395 a_638_3764.t8 a_7830_256.t0 efuse
X396 a_20810_54819.t1 a_638_51026.t11 efuse
X397 a_1340_22414.t1 a_638_19518.t61 efuse
X398 a_20810_10663.t1 BIT_SEL[51].t2 VSS.t581 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X399 a_110_51952.t0 a_154_51864.t1 VSS.t418 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X400 a_7830_30291.t0 a_638_27395.t6 efuse
X401 a_110_22908.t0 a_154_22820.t1 VSS.t162 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X402 a_7830_29555.t0 a_638_27395.t7 efuse
X403 VSS.t482 BIT_SEL[18].t3 a_7830_12904.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X404 a_1340_29923.t1 a_638_27395.t57 efuse
X405 a_638_3764.t24 a_14320_1889.t1 efuse
X406 VDD a_110_6706.t1 a_154_6618.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X407 VDD a_110_61845.t1 a_154_61757.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X408 a_1340_38168.t1 a_638_35272.t14 efuse
X409 a_20810_11031.t1 BIT_SEL[49].t5 VSS.t272 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X410 VSS.t149 BIT_SEL[44].t5 a_14320_15066.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X411 a_110_16636.t0 a_154_16548.t1 VSS.t398 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X412 a_1340_56660.t0 BIT_SEL[9].t4 VSS.t89 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X413 VSS.t525 BIT_SEL[42].t5 a_14320_30291.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X414 a_110_26833.t1 PRESET_N.t6 VDD VDD pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X415 VDD a_110_55573.t1 a_154_55485.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X416 a_7830_46045.t1 a_638_43149.t65 efuse
X417 a_1340_45677.t0 a_638_43149.t9 efuse
X418 a_7830_45309.t1 a_638_43149.t63 efuse
X419 a_110_38662.t0 a_154_38574.t1 VSS.t494 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X420 a_638_3764.t21 a_14320_256.t0 efuse
X421 VSS.t324 BIT_SEL[58].t4 a_20810_53922.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X422 VSS.t500 BIT_SEL[46].t2 a_14320_15434.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X423 a_14320_57556.t0 BIT_SEL[37].t3 VSS.t555 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X424 a_14320_21149.t1 a_638_19518.t63 efuse
X425 a_14320_15066.t0 a_638_11641.t6 efuse
X426 VSS.t211 BIT_SEL[24].t3 a_7830_14169.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X427 a_110_42587.t0 PRESET_N.t7 VDD VDD pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X428 a_7830_20781.t0 a_638_19518.t6 efuse
X429 VDD PRESET_N.t8 a_110_50464.t2 VDD pfet_06v0 ad=0.3172p pd=1.74u as=0.4575p ps=1.97u w=1.22u l=0.5u
X430 a_20810_42171.t0 BIT_SEL[51].t3 VSS.t582 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X431 a_20810_8501.t1 BIT_SEL[61].t1 VSS.t304 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X432 VDD a_110_11079.t7 a_110_10183.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X433 a_1248_11958.t0 a_638_11641.t1 efuse
X434 a_14320_16378.t1 BIT_SEL[45].t2 VSS.t606 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X435 VSS.t611 BIT_SEL[38].t4 a_14320_61063.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X436 a_110_54416.t0 a_154_54328.t1 VSS.t399 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X437 a_20810_5395.t0 a_638_3764.t59 efuse
X438 VSS.t130 BIT_SEL[26].t1 a_7830_14537.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X439 VDD a_110_18060.t4 OUT[2].t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X440 a_1340_3154.t1 BIT_SEL[1].t0 VSS.t107 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X441 a_110_6258.t0 a_154_6170.t1 VSS.t492 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X442 a_638_11641.t8 a_20810_8501.t0 efuse
X443 a_20810_53922.t1 a_638_51026.t13 efuse
X444 a_110_48144.t0 a_154_48056.t1 VSS.t568 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X445 a_14320_36903.t0 a_638_35272.t11 efuse
X446 VDD a_110_14583.t1 a_154_14495.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X447 a_20810_53186.t0 a_638_51026.t19 efuse
X448 a_7830_36535.t0 a_638_35272.t15 efuse
X449 a_14320_54819.t0 a_638_51026.t24 efuse
X450 a_14320_30820.t1 a_638_27395.t68 efuse
X451 a_110_20444.t0 a_154_20356.t1 VSS.t106 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X452 a_638_11641.t68 COL_PROG_N[1].t0 VDD.t289 VDD.t76 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X453 a_638_19518.t11 a_20810_16010.t0 efuse
X454 VSS.t483 BIT_SEL[18].t4 a_7830_60166.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X455 a_1248_27712.t0 a_638_27395.t5 efuse
X456 a_14320_24783.t0 BIT_SEL[43].t3 VSS.t577 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X457 a_1340_5395.t1 a_638_3764.t23 efuse
X458 a_638_19518.t14 a_20810_16906.t1 efuse
X459 VDD a_110_30337.t1 a_154_30249.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X460 VSS.t501 BIT_SEL[46].t3 a_14320_46942.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X461 a_638_27395.t16 a_20810_24255.t0 efuse
X462 VSS.t526 BIT_SEL[42].t6 a_14320_6660.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X463 VDD a_110_18060.t5 a_110_18956.t3 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X464 VSS.t63 BIT_SEL[20].t4 a_7830_60534.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X465 a_14320_46574.t0 a_638_43149.t0 efuse
X466 a_1340_25152.t0 BIT_SEL[9].t5 VSS.t90 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X467 a_1248_43466.t0 a_638_43149.t6 efuse
X468 a_14320_40537.t0 BIT_SEL[43].t4 VSS.t578 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X469 a_638_35272.t16 a_20810_32660.t1 efuse
X470 a_638_35272.t23 a_20810_31764.t0 efuse
X471 VDD a_110_24065.t1 a_154_23977.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X472 a_638_11641.t52 a_1340_8133.t1 efuse
X473 a_1340_54451.t0 a_638_51026.t12 efuse
X474 a_14320_50416.t0 BIT_SEL[33].t2 VSS.t587 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X475 VSS.t131 BIT_SEL[26].t2 a_7830_46045.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X476 a_638_43149.t58 a_20810_40009.t1 efuse
X477 a_1340_25520.t0 BIT_SEL[7].t4 VSS.t119 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X478 a_638_3764.t25 a_7830_2786.t1 efuse
X479 a_638_51026.t55 a_7830_50048.t1 efuse
X480 VDD a_110_46091.t1 a_154_46003.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X481 VSS.t384 BIT_SEL[60].t3 a_20810_30820.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X482 a_7830_34294.t0 BIT_SEL[19].t2 VSS.t153 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X483 a_7738_4081.t0 a_638_3764.t61 efuse
X484 a_638_27395.t12 a_1340_23887.t1 efuse
X485 a_638_11641.t17 a_20810_10294.t1 efuse
X486 a_14320_56291.t0 BIT_SEL[43].t5 VSS.t54 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X487 a_20810_52289.t1 a_638_51026.t8 efuse
X488 a_638_11641.t18 a_20810_11031.t0 efuse
X489 a_7830_34662.t0 BIT_SEL[17].t4 VSS.t264 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X490 VDD.t140 COL_PROG_N[3].t0 a_638_27395.t25 VDD.t86 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X491 VSS.t230 BIT_SEL[12].t1 a_1340_7189.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X492 a_110_50464.t1 PRESET_N.t9 VDD VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X493 a_14320_53186.t0 a_638_51026.t14 efuse
X494 VSS.t385 BIT_SEL[60].t4 a_20810_46574.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X495 a_638_43149.t13 a_1340_39641.t0 efuse
X496 VSS.t520 BIT_SEL[40].t5 a_14320_29923.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X497 VSS.t64 BIT_SEL[20].t5 a_7830_13272.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X498 VSS.t391 BIT_SEL[58].t5 a_20810_61799.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X499 VDD a_110_46539.t1 a_154_46451.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X500 a_638_27395.t58 a_20810_26048.t1 efuse
X501 VDD.t167 COL_PROG_N[3].t1 a_638_27395.t29 VDD.t6 pfet_06v0 ad=9.945p pd=38.77u as=16.83p ps=77.38u w=38.25u l=0.5u
X502 a_638_19518.t46 a_14320_16906.t1 efuse
X503 a_14320_5924.t1 a_638_3764.t18 efuse
X504 VSS.t467 BIT_SEL[14].t3 a_1340_7557.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X505 a_20810_47518.t0 BIT_SEL[63].t2 VSS.t227 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X506 a_638_27395.t8 a_20810_26785.t0 efuse
X507 VSS.t386 BIT_SEL[60].t5 a_20810_62328.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X508 a_14320_61431.t0 a_638_58903.t12 efuse
X509 VDD.t166 COL_PROG_N[5].t0 a_638_43149.t35 VDD.t86 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X510 a_638_11641.t13 a_1340_9766.t1 efuse
X511 a_7830_6292.t0 a_638_3764.t16 efuse
X512 a_20810_1152.t0 BIT_SEL[59].t2 VSS.t561 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X513 VDD a_110_12567.t1 a_154_12479.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X514 a_110_21564.t0 a_154_21476.t1 VSS.t333 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X515 a_638_3764.t3 a_14320_624.t0 efuse
X516 VSS.t445 BIT_SEL[36].t2 a_14320_5395.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X517 a_20810_47886.t0 BIT_SEL[61].t2 VSS.t305 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X518 a_638_43149.t7 a_20810_42539.t0 efuse
X519 a_638_43149.t2 a_20810_41802.t0 efuse
X520 a_638_35272.t4 a_14320_32660.t0 efuse
X521 VDD.t87 COL_PROG_N[7].t0 a_638_58903.t7 VDD.t86 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X522 VDD.t123 COL_PROG_N[5].t1 a_638_43149.t28 VDD.t6 pfet_06v0 ad=9.945p pd=38.77u as=16.83p ps=77.38u w=38.25u l=0.5u
X523 VDD a_110_5362.t1 a_154_5274.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X524 VSS.t348 BIT_SEL[6].t1 a_1340_29555.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X525 a_20810_26048.t0 BIT_SEL[53].t1 VSS.t289 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X526 VSS.t497 BIT_SEL[4].t2 a_1340_44780.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X527 a_638_27395.t56 a_1340_25520.t1 efuse
X528 VSS.t94 BIT_SEL[16].t3 a_7738_4081.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X529 VSS.t617 BIT_SEL[38].t5 a_14320_5924.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X530 a_638_51026.t22 a_1340_48783.t1 efuse
X531 VDD.t88 COL_PROG_N[7].t1 a_638_58903.t8 VDD.t6 pfet_06v0 ad=9.945p pd=38.77u as=16.83p ps=77.38u w=38.25u l=0.5u
X532 a_1340_23311.t1 a_638_19518.t51 efuse
X533 a_638_11641.t10 a_14320_11031.t0 efuse
X534 a_638_58903.t6 a_7830_55763.t1 efuse
X535 a_7738_51343.t0 a_638_51026.t21 efuse
X536 a_638_43149.t14 a_1340_41274.t1 efuse
X537 a_638_58903.t2 a_7830_56660.t0 efuse
X538 VSS.t38 BIT_SEL[28].t0 a_7830_38697.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X539 a_20810_6660.t0 a_638_3764.t14 efuse
X540 VSS.t387 BIT_SEL[60].t6 a_20810_15066.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X541 VDD a_110_60949.t1 a_154_60861.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X542 VDD a_110_44075.t1 a_154_43987.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X543 VSS.t392 BIT_SEL[58].t6 a_20810_30291.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X544 a_110_53072.t0 a_154_52984.t1 VSS.t493 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X545 a_638_19518.t28 a_7830_18171.t1 efuse
X546 a_14228_59220.t1 a_638_58903.t55 efuse
X547 a_1340_39065.t1 a_638_35272.t34 efuse
X548 a_638_19518.t50 a_7830_18908.t1 efuse
X549 VSS.t177 BIT_SEL[62].t3 a_20810_15434.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X550 VSS.t39 BIT_SEL[28].t1 a_7830_54451.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X551 a_638_27395.t48 a_14320_26785.t1 efuse
X552 a_1340_18908.t1 BIT_SEL[1].t1 VSS.t108 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X553 a_20810_57556.t1 BIT_SEL[53].t2 VSS.t366 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X554 a_110_37766.t0 a_154_37678.t1 VSS.t124 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X555 VSS.t36 BIT_SEL[8].t0 a_1340_6292.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X556 a_20810_15066.t1 a_638_11641.t49 efuse
X557 a_638_51026.t46 a_20810_48783.t1 efuse
X558 a_638_35272.t55 a_7830_33925.t1 efuse
X559 VSS.t10 BIT_SEL[0].t4 a_1248_11958.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X560 a_7830_40009.t0 BIT_SEL[29].t1 VSS.t308 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X561 a_638_35272.t61 a_7830_34662.t1 efuse
X562 a_638_11641.t26 SENSE.t6 a_110_11079.t5 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X563 a_20810_16378.t0 BIT_SEL[61].t3 VSS.t306 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X564 VSS.t315 BIT_SEL[54].t5 a_20810_61063.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X565 VSS.t4 BIT_SEL[30].t0 a_7830_54819.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X566 a_638_43149.t52 a_14320_42539.t1 efuse
X567 a_14320_57028.t0 BIT_SEL[39].t2 VSS.t422 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X568 a_638_51026.t59 a_1340_50416.t0 efuse
X569 a_20810_30820.t1 a_638_27395.t59 efuse
X570 VSS.t472 BIT_SEL[46].t4 a_14320_23311.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X571 VSS.t217 BIT_SEL[22].t4 a_7830_21678.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X572 a_1340_21678.t1 a_638_19518.t60 efuse
X573 a_110_9207.t0 a_154_9119.t1 VSS.t469 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X574 VDD a_110_13687.t1 a_154_13599.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X575 a_20810_24783.t0 BIT_SEL[59].t3 VSS.t562 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X576 VSS.t459 BIT_SEL[62].t4 a_20810_46942.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X577 a_14320_23887.t1 BIT_SEL[47].t2 VSS.t42 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X578 a_638_58903.t19 a_1340_57925.t0 efuse
X579 a_20810_46574.t1 a_638_43149.t57 efuse
X580 a_1340_8133.t0 BIT_SEL[15].t4 VSS.t246 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X581 a_110_50464.t0 PRESET_N.t10 VDD VDD pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X582 VSS.t11 BIT_SEL[0].t5 a_1248_43466.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X583 a_20810_40537.t0 BIT_SEL[59].t4 VSS.t563 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X584 a_1340_37432.t1 a_638_35272.t38 efuse
X585 a_20810_50416.t0 BIT_SEL[49].t6 VSS.t425 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X586 a_20810_14169.t0 a_638_11641.t15 efuse
X587 a_7830_49679.t0 BIT_SEL[21].t2 VSS.t442 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X588 a_20810_13272.t0 a_638_11641.t32 efuse
X589 a_638_3764.t44 a_7830_1889.t0 efuse
X590 VSS.t193 BIT_SEL[2].t2 a_1340_44412.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X591 a_638_51026.t28 a_14320_48783.t0 efuse
X592 VDD a_110_45195.t1 a_154_45107.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X593 a_20810_56291.t1 BIT_SEL[59].t5 VSS.t564 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X594 VSS.t218 BIT_SEL[22].t5 a_7830_53186.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X595 VSS.t484 BIT_SEL[18].t5 a_7830_5027.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X596 a_638_58903.t38 a_20810_57925.t1 efuse
X597 a_14320_55395.t1 BIT_SEL[47].t3 VSS.t43 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X598 VDD a_110_29889.t1 a_154_29801.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X599 a_20810_29026.t0 a_638_27395.t34 efuse
X600 a_20810_29923.t0 a_638_27395.t54 efuse
X601 VSS.t212 BIT_SEL[24].t4 a_7830_53554.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X602 VSS.t341 BIT_SEL[56].t6 a_20810_29923.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X603 a_1340_14537.t1 a_638_11641.t53 efuse
X604 a_638_58903.t65 a_14320_57028.t1 efuse
X605 a_1340_33397.t0 BIT_SEL[7].t5 VSS.t120 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X606 a_7830_16906.t0 BIT_SEL[27].t1 VSS.t548 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X607 a_7830_53554.t1 a_638_51026.t48 efuse
X608 VDD a_110_50464.t7 a_110_49568.t1 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X609 VDD a_110_31942.t1 a_154_31854.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X610 VDD PRESET_N.t11 a_110_11079.t1 VDD pfet_06v0 ad=0.3172p pd=1.74u as=0.4575p ps=1.97u w=1.22u l=0.5u
X611 a_14320_55763.t0 BIT_SEL[45].t3 VSS.t607 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X612 a_20810_45677.t0 a_638_43149.t21 efuse
X613 VSS.t99 BIT_SEL[30].t1 a_7830_39065.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X614 a_20810_44780.t0 a_638_43149.t44 efuse
X615 a_1340_18540.t1 BIT_SEL[3].t3 VSS.t186 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X616 a_14320_33925.t1 BIT_SEL[37].t4 VSS.t556 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X617 a_1340_41802.t0 BIT_SEL[5].t2 VSS.t72 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X618 a_1340_30291.t1 a_638_27395.t44 efuse
X619 a_7830_39641.t1 BIT_SEL[31].t0 VSS.t300 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X620 a_110_3202.t2 PRESET_N.t12 VDD VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X621 a_14320_13272.t1 a_638_11641.t58 efuse
X622 a_110_24513.t0 a_154_24425.t1 VSS.t160 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X623 a_7830_2417.t0 BIT_SEL[21].t3 VSS.t443 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X624 a_7830_62328.t1 a_638_58903.t48 efuse
X625 a_1340_46045.t1 a_638_43149.t26 efuse
X626 VSS.t150 BIT_SEL[44].t6 a_14320_22943.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X627 a_638_3764.t65 a_20810_2786.t1 efuse
X628 a_7830_12904.t0 a_638_11641.t19 efuse
X629 a_7830_48414.t0 BIT_SEL[27].t2 VSS.t549 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X630 a_110_34710.t2 PRESET_N.t13 VDD VDD pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X631 a_20718_4081.t0 a_638_3764.t54 efuse
X632 VDD a_110_8311.t1 a_154_8223.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X633 a_7830_21149.t1 a_638_19518.t29 efuse
X634 a_638_58903.t28 a_14320_57925.t0 efuse
X635 VSS.t103 BIT_SEL[24].t5 a_7830_22046.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X636 a_14320_29026.t1 a_638_27395.t63 efuse
X637 a_7830_28658.t0 a_638_27395.t46 efuse
X638 a_638_11641.t41 a_20810_8133.t1 efuse
X639 a_638_11641.t48 a_20810_9029.t1 efuse
X640 a_14320_24255.t0 BIT_SEL[45].t4 VSS.t608 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X641 VSS.t487 BIT_SEL[32].t1 a_14228_59220.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X642 a_20718_59220.t0 a_638_58903.t49 efuse
X643 a_7830_36903.t1 a_638_35272.t47 efuse
X644 VSS.t132 BIT_SEL[26].t3 a_7830_22414.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X645 a_14320_44780.t1 a_638_43149.t53 efuse
X646 VDD a_110_22460.t1 a_154_22372.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X647 a_110_56021.t0 a_154_55933.t1 VSS.t506 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X648 a_1340_52657.t1 a_638_51026.t44 efuse
X649 a_7830_44412.t1 a_638_43149.t62 efuse
X650 VSS.t405 a_110_41691.t2 OUT[5].t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X651 VSS.t37 BIT_SEL[8].t1 a_1340_37800.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X652 a_1340_10294.t0 BIT_SEL[5].t3 VSS.t73 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X653 a_7830_10663.t0 BIT_SEL[19].t3 VSS.t154 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X654 a_14320_32660.t1 BIT_SEL[43].t6 VSS.t55 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X655 a_638_27395.t18 a_20810_24783.t1 efuse
X656 a_638_27395.t17 a_20810_23887.t0 efuse
X657 a_7830_11031.t0 BIT_SEL[17].t5 VSS.t178 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X658 a_20810_57028.t0 BIT_SEL[55].t2 VSS.t595 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X659 VSS.t460 BIT_SEL[62].t5 a_20810_23311.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X660 a_14320_18171.t1 BIT_SEL[37].t5 VSS.t557 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X661 a_1340_60166.t1 a_638_58903.t57 efuse
X662 a_638_43149.t68 a_20810_39641.t1 efuse
X663 a_638_3764.t22 a_7830_624.t1 efuse
X664 VSS.t81 BIT_SEL[48].t1 a_20718_4081.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X665 VDD a_110_51952.t1 a_154_51864.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X666 a_638_43149.t37 a_20810_40537.t1 efuse
X667 VDD a_110_22908.t1 a_154_22820.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X668 a_14320_2786.t0 BIT_SEL[35].t3 VSS.t454 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X669 a_110_15031.t0 a_154_14943.t1 VSS.t537 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X670 VSS.t235 BIT_SEL[26].t4 a_7830_53922.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X671 a_20810_23887.t1 BIT_SEL[63].t3 VSS.t219 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X672 a_638_3764.t34 a_14320_2417.t1 efuse
X673 VDD.t261 COL_PROG_N[2].t0 a_638_19518.t57 VDD.t86 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X674 VDD a_110_16636.t1 a_154_16548.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X675 a_7830_42171.t0 BIT_SEL[19].t4 VSS.t155 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X676 a_638_58903.t20 a_14320_55395.t0 efuse
X677 VSS.t194 BIT_SEL[2].t3 a_1340_20781.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X678 a_638_11641.t44 a_14320_9029.t1 efuse
X679 VDD a_110_38662.t1 a_154_38574.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X680 VSS.t488 BIT_SEL[32].t2 a_14228_27712.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X681 VSS.t334 a_110_57445.t3 a_110_58341.t4 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X682 VDD.t247 COL_PROG_N[2].t1 a_638_19518.t52 VDD.t6 pfet_06v0 ad=9.945p pd=38.77u as=16.83p ps=77.38u w=38.25u l=0.5u
X683 a_14320_50048.t1 BIT_SEL[35].t4 VSS.t455 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X684 VSS.t515 a_110_10183.t3 OUT[1].t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X685 VSS.t115 BIT_SEL[34].t3 a_14320_28658.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X686 a_14320_61799.t0 a_638_58903.t33 efuse
X687 VDD a_110_54416.t1 a_154_54328.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X688 a_638_27395.t53 a_14320_24783.t1 efuse
X689 a_20810_5027.t1 a_638_3764.t30 efuse
X690 a_20810_55395.t0 BIT_SEL[63].t4 VSS.t220 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X691 VDD a_110_48144.t1 a_154_48056.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X692 VDD.t254 COL_PROG_N[6].t0 a_638_51026.t63 VDD.t86 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X693 a_638_58903.t39 a_20810_57028.t1 efuse
X694 VSS.t166 BIT_SEL[4].t3 a_1340_36903.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X695 VDD a_110_20444.t1 a_154_20356.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X696 VSS.t195 BIT_SEL[2].t4 a_1340_52289.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X697 a_638_43149.t25 a_14320_40537.t1 efuse
X698 a_7830_9029.t0 BIT_SEL[27].t3 VSS.t550 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X699 a_1340_15434.t1 a_638_11641.t30 efuse
X700 a_20810_55763.t0 BIT_SEL[61].t4 VSS.t290 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X701 a_638_51026.t10 a_1340_48414.t0 efuse
X702 VDD.t246 COL_PROG_N[6].t1 a_638_51026.t60 VDD.t6 pfet_06v0 ad=9.945p pd=38.77u as=16.83p ps=77.38u w=38.25u l=0.5u
X703 VSS.t361 BIT_SEL[6].t2 a_1340_37432.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X704 a_20810_33925.t1 BIT_SEL[53].t3 VSS.t367 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X705 VSS.t138 BIT_SEL[28].t2 a_7830_30820.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X706 VSS.t167 BIT_SEL[4].t4 a_1340_52657.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X707 VSS.t473 BIT_SEL[46].t5 a_14320_62696.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X708 a_14320_33029.t1 BIT_SEL[41].t1 VSS.t206 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X709 a_638_11641.t35 a_7830_10294.t1 efuse
X710 a_638_11641.t64 a_7830_11031.t1 efuse
X711 a_638_58903.t26 a_1340_55763.t1 efuse
X712 a_638_58903.t42 a_7830_56291.t1 efuse
X713 a_1340_40906.t1 BIT_SEL[9].t6 VSS.t91 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X714 VSS.t15 BIT_SEL[10].t1 a_1340_38168.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X715 VSS.t311 a_110_25937.t3 a_110_26833.t3 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X716 a_1340_31188.t1 a_638_27395.t60 efuse
X717 VSS.t139 BIT_SEL[28].t3 a_7830_46574.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X718 VSS.t388 BIT_SEL[60].t7 a_20810_22943.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X719 a_14320_22046.t1 a_638_19518.t54 efuse
X720 a_1340_7189.t1 a_638_3764.t55 efuse
X721 VSS.t236 BIT_SEL[26].t5 a_7830_61799.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X722 a_1340_26417.t1 BIT_SEL[3].t4 VSS.t187 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X723 a_638_3764.t48 a_1340_1521.t1 efuse
X724 VSS.t406 a_110_41691.t3 a_110_42587.t4 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X725 a_638_27395.t61 a_7830_26048.t1 efuse
X726 a_14320_48783.t1 BIT_SEL[41].t2 VSS.t207 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X727 a_1340_46942.t0 a_638_43149.t1 efuse
X728 a_638_27395.t15 a_7830_26785.t0 efuse
X729 VSS.t140 BIT_SEL[28].t4 a_7830_62328.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X730 a_7830_47518.t1 BIT_SEL[31].t1 VSS.t284 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X731 a_1340_26785.t0 BIT_SEL[1].t2 VSS.t109 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X732 a_110_45643.t0 a_154_45555.t1 VSS.t57 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X733 a_14320_37800.t1 a_638_35272.t37 efuse
X734 a_14320_3154.t0 BIT_SEL[33].t3 VSS.t588 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X735 a_7830_1889.t1 BIT_SEL[23].t4 VSS.t163 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X736 VDD a_110_882.t1 a_154_794.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X737 a_638_3764.t49 a_7830_3154.t0 efuse
X738 VSS.t24 BIT_SEL[50].t4 a_20810_5027.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X739 a_110_7602.t0 a_154_7514.t1 VSS.t123 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X740 a_7830_47886.t0 BIT_SEL[29].t2 VSS.t309 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X741 a_638_43149.t16 a_7830_42539.t0 efuse
X742 a_638_43149.t40 a_7830_41802.t1 efuse
X743 a_20810_24255.t1 BIT_SEL[61].t5 VSS.t291 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X744 VSS.t12 BIT_SEL[0].t6 a_1248_19835.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X745 a_1340_13801.t1 a_638_11641.t63 efuse
X746 VSS.t82 BIT_SEL[48].t2 a_20718_59220.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X747 a_1340_42539.t1 BIT_SEL[1].t3 VSS.t144 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X748 a_7830_26048.t0 BIT_SEL[21].t4 VSS.t444 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X749 a_14320_5395.t1 a_638_3764.t62 efuse
X750 VSS.t168 BIT_SEL[4].t5 a_1340_21149.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X751 a_638_19518.t42 a_7830_16378.t1 efuse
X752 a_14320_16010.t1 BIT_SEL[47].t4 VSS.t44 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X753 VSS.t474 BIT_SEL[46].t6 a_14320_31188.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X754 a_638_19518.t13 a_7830_17275.t0 efuse
X755 a_638_58903.t37 a_1340_57556.t1 efuse
X756 VDD a_110_21564.t1 a_154_21476.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X757 a_20810_32660.t0 BIT_SEL[59].t6 VSS.t433 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X758 a_1340_29555.t1 a_638_27395.t42 efuse
X759 VSS.t395 a_110_2306.t4 a_110_3202.t4 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X760 a_638_35272.t41 a_7830_32132.t1 efuse
X761 a_14228_19835.t1 a_638_19518.t35 efuse
X762 a_20810_62696.t1 a_638_58903.t35 efuse
X763 a_1340_58293.t1 BIT_SEL[1].t4 VSS.t145 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X764 a_110_39819.t0 a_154_39731.t1 VSS.t417 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X765 a_638_35272.t64 a_7830_33029.t1 efuse
X766 a_14320_31764.t1 BIT_SEL[47].t5 VSS.t45 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X767 VSS.t446 BIT_SEL[36].t3 a_14320_29026.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X768 a_638_11641.t67 COL_PROG_N[1].t1 VDD.t282 VDD.t2 pfet_06v0 ad=16.83p pd=77.38u as=9.945p ps=38.77u w=38.25u l=0.5u
X769 VSS.t141 BIT_SEL[28].t5 a_7830_15066.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X770 VSS.t237 BIT_SEL[26].t6 a_7830_30291.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X771 a_20810_2417.t0 BIT_SEL[53].t4 VSS.t368 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X772 a_20810_18171.t1 BIT_SEL[53].t5 VSS.t369 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X773 a_1340_45309.t1 a_638_43149.t60 efuse
X774 a_14320_17275.t1 BIT_SEL[41].t3 VSS.t198 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X775 a_14228_35589.t1 a_638_35272.t30 efuse
X776 VSS.t100 BIT_SEL[30].t2 a_7830_15434.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X777 a_7830_57556.t0 BIT_SEL[21].t5 VSS.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X778 a_20810_256.t1 BIT_SEL[63].t5 VSS.t221 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X779 VDD.t120 COL_PROG_N[1].t2 a_638_11641.t20 VDD.t6 pfet_06v0 ad=9.945p pd=38.77u as=16.83p ps=77.38u w=38.25u l=0.5u
X780 a_110_14135.t0 a_154_14047.t1 VSS.t402 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X781 VSS.t151 BIT_SEL[44].t7 a_14320_7189.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X782 a_14320_17643.t0 BIT_SEL[39].t3 VSS.t421 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X783 a_20810_6292.t0 a_638_3764.t52 efuse
X784 a_7830_16378.t0 BIT_SEL[29].t3 VSS.t310 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X785 VSS.t34 BIT_SEL[22].t6 a_7830_61063.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X786 VDD a_110_53072.t1 a_154_52984.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X787 a_20810_624.t1 BIT_SEL[61].t6 VSS.t292 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X788 VSS.t83 BIT_SEL[48].t3 a_20718_27712.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X789 a_638_19518.t44 a_1340_18540.t0 efuse
X790 a_638_3764.t37 a_20810_1152.t1 efuse
X791 VSS.t475 BIT_SEL[46].t7 a_14320_7557.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X792 a_20810_50048.t0 BIT_SEL[51].t4 VSS.t583 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X793 VDD a_110_37766.t1 a_154_37678.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X794 a_1340_41274.t0 BIT_SEL[7].t6 VSS.t121 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X795 VSS.t23 BIT_SEL[50].t5 a_20810_28658.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X796 a_7830_24783.t0 BIT_SEL[27].t4 VSS.t542 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X797 VDD a_110_3202.t6 a_110_2306.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X798 a_110_11079.t2 PRESET_N.t14 VDD VDD pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X799 a_20810_61063.t1 a_638_58903.t67 efuse
X800 a_20810_61799.t1 a_638_58903.t40 efuse
X801 VSS.t101 BIT_SEL[30].t3 a_7830_46942.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X802 a_638_3764.t60 a_1340_1152.t1 efuse
X803 a_638_35272.t54 a_1340_34294.t0 efuse
X804 a_14320_62696.t0 a_638_58903.t41 efuse
X805 a_7830_1521.t1 BIT_SEL[25].t3 VSS.t281 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X806 a_638_51026.t32 a_7830_47518.t0 efuse
X807 a_14320_49151.t1 BIT_SEL[39].t4 VSS.t411 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X808 a_7830_40537.t0 BIT_SEL[27].t5 VSS.t543 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X809 a_7830_50416.t1 BIT_SEL[17].t6 VSS.t179 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X810 VSS.t362 BIT_SEL[6].t3 a_1340_13801.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X811 a_7830_13272.t1 a_638_11641.t36 efuse
X812 a_1340_62328.t1 a_638_58903.t60 efuse
X813 a_14320_52289.t0 a_638_51026.t17 efuse
X814 a_638_19518.t27 a_20810_18540.t1 efuse
X815 a_1340_256.t0 BIT_SEL[15].t5 VSS.t247 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X816 VSS.t461 BIT_SEL[62].t6 a_20810_62696.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X817 a_7830_56291.t0 BIT_SEL[27].t6 VSS.t544 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X818 a_20810_33029.t0 BIT_SEL[57].t2 VSS.t374 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X819 a_638_19518.t22 a_14320_17643.t1 efuse
X820 a_1340_5027.t1 a_638_3764.t32 efuse
X821 a_638_58903.t44 a_7830_57925.t1 efuse
X822 a_638_35272.t51 a_20810_34294.t1 efuse
X823 a_1340_624.t1 BIT_SEL[13].t3 VSS.t250 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X824 a_110_59829.t0 a_154_59741.t1 VSS.t428 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X825 a_7830_29026.t1 a_638_27395.t50 efuse
X826 VSS.t104 BIT_SEL[24].t6 a_7830_29923.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X827 a_20810_60166.t1 a_638_58903.t22 efuse
X828 VSS.t363 BIT_SEL[6].t4 a_1340_45309.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X829 a_638_35272.t53 a_14320_33397.t1 efuse
X830 a_1340_9398.t0 BIT_SEL[9].t7 VSS.t92 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X831 a_20810_48783.t0 BIT_SEL[57].t3 VSS.t375 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X832 a_14320_32132.t0 BIT_SEL[45].t5 VSS.t507 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X833 a_110_28993.t0 a_154_28905.t1 VSS.t431 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X834 VSS.t521 BIT_SEL[40].t6 a_14320_6292.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X835 a_14320_61063.t1 a_638_58903.t43 efuse
X836 a_7830_44780.t1 a_638_43149.t66 efuse
X837 a_638_51026.t42 a_7830_49151.t0 efuse
X838 a_1340_9766.t0 BIT_SEL[7].t7 VSS.t122 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X839 VSS.t125 BIT_SEL[8].t2 a_1340_45677.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X840 a_7830_22943.t1 a_638_19518.t16 efuse
X841 a_110_44747.t0 a_154_44659.t1 VSS.t299 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X842 a_110_6706.t0 a_154_6618.t1 VSS.t609 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X843 a_20810_9029.t0 BIT_SEL[59].t7 VSS.t434 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X844 VSS.t126 BIT_SEL[8].t3 a_1340_61431.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X845 a_638_19518.t31 a_14320_18540.t1 efuse
X846 a_20810_16010.t1 BIT_SEL[63].t6 VSS.t222 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X847 a_7830_38697.t1 a_638_35272.t62 efuse
X848 VSS.t462 BIT_SEL[62].t7 a_20810_31188.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X849 VSS.t238 BIT_SEL[26].t7 a_7830_6660.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X850 a_14320_8133.t0 BIT_SEL[47].t6 VSS.t46 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X851 VSS.t196 BIT_SEL[2].t5 a_1340_12904.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X852 a_638_35272.t25 a_14320_34294.t0 efuse
X853 a_20718_19835.t0 a_638_19518.t41 efuse
X854 a_638_58903.t52 a_1340_56660.t1 efuse
X855 a_20810_31764.t1 BIT_SEL[63].t7 VSS.t223 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X856 VSS.t356 BIT_SEL[52].t5 a_20810_29026.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X857 VDD a_110_24513.t1 a_154_24425.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X858 a_638_51026.t65 a_14320_47886.t1 efuse
X859 a_20810_17275.t0 BIT_SEL[57].t4 VSS.t376 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X860 a_7738_59220.t1 a_638_58903.t63 efuse
X861 VSS.t489 BIT_SEL[32].t3 a_14228_35589.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X862 a_20718_35589.t0 a_638_35272.t50 efuse
X863 a_110_26833.t0 PRESET_N.t15 VDD VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X864 VDD PRESET_N.t16 a_110_3202.t1 VDD pfet_06v0 ad=0.3172p pd=1.74u as=0.4575p ps=1.97u w=1.22u l=0.5u
X865 VSS.t127 BIT_SEL[8].t4 a_1340_14169.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X866 a_14320_57925.t1 BIT_SEL[35].t5 VSS.t456 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X867 a_638_3764.t45 a_20810_3154.t1 efuse
X868 a_20810_1889.t0 BIT_SEL[55].t3 VSS.t596 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X869 a_20810_17643.t0 BIT_SEL[55].t4 VSS.t597 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X870 VSS.t273 BIT_SEL[34].t4 a_14320_36535.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X871 a_1340_20781.t1 a_638_19518.t34 efuse
X872 a_110_13239.t0 a_154_13151.t1 VSS.t412 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X873 VSS.t65 BIT_SEL[32].t4 a_14228_51343.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X874 a_1340_8501.t1 BIT_SEL[13].t4 VSS.t251 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X875 VSS.t16 BIT_SEL[10].t2 a_1340_14537.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X876 a_638_58903.t23 a_20810_56660.t1 efuse
X877 a_7830_57028.t1 BIT_SEL[23].t5 VSS.t538 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X878 VDD a_110_56021.t1 a_154_55933.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X879 VDD a_110_41691.t4 OUT[5].t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X880 a_1340_36535.t1 a_638_35272.t56 efuse
X881 VSS.t102 BIT_SEL[30].t4 a_7830_23311.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X882 a_638_3764.t40 a_1340_3154.t0 efuse
X883 a_110_39110.t0 a_154_39022.t1 VSS.t413 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X884 VSS.t197 BIT_SEL[2].t6 a_1340_60166.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X885 a_7830_54819.t0 a_638_51026.t25 efuse
X886 a_638_19518.t30 a_14320_16010.t0 efuse
X887 a_110_58341.t0 PRESET_N.t17 VDD VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X888 a_638_58903.t53 a_1340_58293.t0 efuse
X889 a_7830_23887.t1 BIT_SEL[31].t2 VSS.t285 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X890 a_1340_6292.t1 a_638_3764.t38 efuse
X891 VDD a_110_2306.t5 OUT[0].t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X892 a_14320_14169.t1 a_638_11641.t45 efuse
X893 a_638_51026.t56 a_14320_49679.t1 efuse
X894 VSS.t511 BIT_SEL[20].t6 a_7830_5395.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X895 VSS.t169 BIT_SEL[4].t6 a_1340_60534.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X896 a_20810_49151.t0 BIT_SEL[55].t5 VSS.t269 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X897 a_638_35272.t44 a_14320_31764.t0 efuse
X898 VDD a_110_5810.t1 a_154_5722.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X899 VSS.t17 BIT_SEL[10].t3 a_1340_46045.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X900 VSS.t241 a_110_33814.t4 a_110_34710.t3 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X901 a_14320_22414.t1 a_638_19518.t56 efuse
X902 VSS.t35 BIT_SEL[22].t7 a_7830_5924.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X903 VDD a_110_15031.t1 a_154_14943.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X904 a_110_30785.t0 a_154_30697.t1 VSS.t143 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X905 a_7830_7557.t0 a_638_3764.t15 efuse
X906 a_1340_34294.t1 BIT_SEL[3].t5 VSS.t188 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X907 a_14320_29923.t1 a_638_27395.t24 efuse
X908 a_638_3764.t63 a_14320_2786.t1 efuse
X909 VSS.t142 a_110_18956.t6 a_110_18060.t0 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X910 VSS.t571 a_110_49568.t3 a_110_50464.t4 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X911 a_14320_38168.t1 a_638_35272.t49 efuse
X912 a_638_19518.t53 a_20810_17643.t1 efuse
X913 a_14320_56660.t1 BIT_SEL[41].t4 VSS.t199 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X914 a_110_434.t0 a_154_346.t1 VSS.t380 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X915 VDD a_110_57445.t4 a_110_58341.t5 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X916 a_7830_55395.t1 BIT_SEL[31].t3 VSS.t286 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X917 a_638_11641.t22 a_7830_8501.t1 efuse
X918 a_638_58903.t46 a_14320_56660.t0 efuse
X919 a_7830_53922.t1 a_638_51026.t49 efuse
X920 a_14320_45677.t1 a_638_43149.t45 efuse
X921 a_1340_34662.t1 BIT_SEL[1].t5 VSS.t146 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X922 VDD a_110_10183.t4 OUT[1].t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X923 a_638_11641.t24 a_7830_9398.t0 efuse
X924 a_110_53520.t0 a_154_53432.t1 VSS.t438 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X925 a_7830_53186.t1 a_638_51026.t30 efuse
X926 a_638_35272.t21 a_20810_33397.t1 efuse
X927 VSS.t170 BIT_SEL[4].t7 a_1340_13272.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X928 a_1340_53554.t0 a_638_51026.t9 efuse
X929 a_7830_55763.t0 BIT_SEL[29].t4 VSS.t294 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X930 a_110_40267.t0 a_154_40179.t1 VSS.t463 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X931 a_20810_32132.t1 BIT_SEL[61].t7 VSS.t293 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X932 a_638_19518.t20 a_7830_16906.t1 efuse
X933 a_110_5362.t0 a_154_5274.t1 VSS.t302 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X934 a_14228_11958.t1 a_638_11641.t39 efuse
X935 a_638_19518.t37 a_1340_16378.t1 efuse
X936 a_7830_33925.t0 BIT_SEL[21].t6 VSS.t2 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X937 a_638_27395.t27 a_7830_24255.t1 efuse
X938 a_110_62293.t0 a_154_62205.t1 VSS.t416 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X939 a_7830_61431.t1 a_638_58903.t56 efuse
X940 a_638_27395.t33 a_7830_25152.t1 efuse
X941 a_20810_1521.t0 BIT_SEL[57].t5 VSS.t377 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X942 a_1340_1152.t0 BIT_SEL[11].t2 VSS.t403 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X943 a_638_35272.t45 a_1340_32132.t1 efuse
X944 a_638_35272.t65 a_7830_32660.t1 efuse
X945 VDD a_110_8759.t1 a_154_8671.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X946 a_110_46987.t0 a_154_46899.t1 VSS.t401 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X947 a_638_43149.t41 a_7830_40009.t1 efuse
X948 a_14228_27712.t1 a_638_27395.t35 efuse
X949 VSS.t133 BIT_SEL[28].t6 a_7830_22943.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X950 a_638_43149.t31 a_7830_40906.t0 efuse
X951 a_638_27395.t20 COL_PROG_N[3].t2 VDD.t125 VDD.t2 pfet_06v0 ad=16.83p pd=77.38u as=9.945p ps=38.77u w=38.25u l=0.5u
X952 a_14320_25152.t0 BIT_SEL[41].t5 VSS.t200 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X953 a_14320_54451.t1 a_638_51026.t51 efuse
X954 a_14228_43466.t1 a_638_43149.t67 efuse
X955 VDD a_110_25937.t4 a_110_26833.t5 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X956 a_638_3764.t39 a_20810_1889.t1 efuse
X957 a_638_27395.t19 COL_PROG_N[3].t3 VDD.t124 VDD.t76 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X958 a_638_11641.t25 a_1340_10663.t0 efuse
X959 a_110_56469.t0 a_154_56381.t1 VSS.t570 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X960 a_1248_51343.t1 a_638_51026.t43 efuse
X961 VSS.t231 BIT_SEL[12].t2 a_1340_38697.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X962 a_110_22012.t0 a_154_21924.t1 VSS.t602 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X963 a_638_43149.t32 COL_PROG_N[5].t2 VDD.t141 VDD.t2 pfet_06v0 ad=16.83p pd=77.38u as=9.945p ps=38.77u w=38.25u l=0.5u
X964 a_14320_25520.t0 BIT_SEL[39].t5 VSS.t410 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X965 a_1340_6660.t1 a_638_3764.t42 efuse
X966 a_638_51026.t39 a_20810_47886.t1 efuse
X967 VDD a_110_41691.t5 a_110_42587.t3 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X968 a_7830_24255.t0 BIT_SEL[29].t5 VSS.t295 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X969 a_638_19518.t18 a_1340_18171.t1 efuse
X970 VSS.t95 BIT_SEL[16].t4 a_7738_59220.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X971 VSS.t84 BIT_SEL[48].t4 a_20718_35589.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X972 VSS.t232 BIT_SEL[12].t3 a_1340_54451.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X973 a_20810_57925.t0 BIT_SEL[51].t5 VSS.t584 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X974 VDD a_110_45643.t1 a_154_45555.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X975 a_638_27395.t13 a_1340_26417.t0 efuse
X976 a_20810_23311.t1 a_638_19518.t43 efuse
X977 a_638_58903.t9 COL_PROG_N[7].t2 VDD.t89 VDD.t2 pfet_06v0 ad=16.83p pd=77.38u as=9.945p ps=38.77u w=38.25u l=0.5u
X978 a_638_43149.t24 COL_PROG_N[5].t3 VDD.t122 VDD.t76 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X979 a_1340_40009.t1 BIT_SEL[13].t5 VSS.t252 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X980 VSS.t22 BIT_SEL[50].t6 a_20810_36535.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X981 a_638_35272.t26 a_1340_33925.t1 efuse
X982 a_7830_32660.t0 BIT_SEL[27].t7 VSS.t545 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X983 VDD.t209 COL_PROG_N[4].t2 a_638_35272.t59 VDD.t86 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X984 VSS.t466 BIT_SEL[14].t4 a_1340_54819.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X985 VSS.t502 BIT_SEL[48].t5 a_20718_51343.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X986 a_110_15479.t0 a_154_15391.t1 VSS.t437 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X987 a_1340_60534.t1 a_638_58903.t27 efuse
X988 a_638_43149.t51 a_1340_42171.t0 efuse
X989 a_638_11641.t12 a_20810_10663.t0 efuse
X990 a_638_58903.t10 COL_PROG_N[7].t3 VDD.t90 VDD.t76 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X991 a_638_51026.t27 a_1340_47518.t1 efuse
X992 a_20810_39065.t1 a_638_35272.t29 efuse
X993 a_7830_18171.t0 BIT_SEL[21].t7 VSS.t3 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X994 VDD.t7 COL_PROG_N[4].t3 a_638_35272.t3 VDD.t6 pfet_06v0 ad=9.945p pd=38.77u as=16.83p ps=77.38u w=38.25u l=0.5u
X995 VSS.t364 BIT_SEL[6].t5 a_1340_21678.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X996 a_638_11641.t7 a_14320_9766.t0 efuse
X997 a_110_38214.t0 a_154_38126.t1 VSS.t546 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X998 VDD a_110_1330.t1 a_154_1242.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X999 VSS.t393 BIT_SEL[58].t7 a_20810_6660.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1000 VDD a_110_39819.t1 a_154_39731.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1001 a_638_27395.t31 a_20810_26417.t1 efuse
X1002 a_638_51026.t29 a_20810_49679.t1 efuse
X1003 VDD PRESET_N.t18 a_110_18956.t1 VDD pfet_06v0 ad=0.3172p pd=1.74u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1004 a_638_51026.t50 a_20810_50416.t1 efuse
X1005 VSS.t618 BIT_SEL[38].t6 a_14320_29555.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1006 a_14320_7189.t1 a_638_3764.t58 efuse
X1007 VSS.t447 BIT_SEL[36].t4 a_14320_44780.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1008 VSS.t96 BIT_SEL[16].t5 a_7738_27712.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1009 a_638_27395.t37 a_14320_25520.t1 efuse
X1010 a_20810_22414.t1 a_638_19518.t36 efuse
X1011 a_20810_21678.t0 a_638_19518.t25 efuse
X1012 a_7830_50048.t0 BIT_SEL[19].t5 VSS.t156 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1013 a_1340_49679.t1 BIT_SEL[5].t4 VSS.t74 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1014 a_638_43149.t42 a_20810_42171.t1 efuse
X1015 VDD a_110_14135.t1 a_154_14047.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1016 VSS.t470 BIT_SEL[18].t6 a_7830_28658.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1017 a_14320_23311.t0 a_638_19518.t9 efuse
X1018 a_7830_15066.t1 a_638_11641.t46 efuse
X1019 a_638_43149.t43 a_14320_41274.t1 efuse
X1020 VSS.t165 BIT_SEL[6].t6 a_1340_53186.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1021 a_20810_38168.t1 a_638_35272.t40 efuse
X1022 a_20810_56660.t0 BIT_SEL[57].t6 VSS.t378 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1023 a_638_51026.t58 a_1340_49151.t1 efuse
X1024 a_110_36870.t0 a_154_36782.t1 VSS.t400 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1025 a_20810_37432.t1 a_638_35272.t67 efuse
X1026 a_638_11641.t27 a_14320_10663.t0 efuse
X1027 a_14320_39065.t0 a_638_35272.t46 efuse
X1028 a_1340_22943.t1 a_638_19518.t40 efuse
X1029 a_638_3764.t67 a_20810_1521.t1 efuse
X1030 VSS.t128 BIT_SEL[8].t5 a_1340_53554.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1031 a_14320_18908.t0 BIT_SEL[33].t4 VSS.t589 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1032 a_110_52624.t0 a_154_52536.t1 VSS.t228 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1033 a_7830_30820.t1 a_638_27395.t32 efuse
X1034 a_1340_16906.t0 BIT_SEL[11].t3 VSS.t298 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1035 VSS.t465 BIT_SEL[14].t5 a_1340_39065.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1036 a_20718_11958.t0 a_638_11641.t47 efuse
X1037 VSS.t66 BIT_SEL[32].t5 a_14228_11958.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1038 a_638_19518.t55 a_7830_18540.t1 efuse
X1039 a_1340_38697.t1 a_638_35272.t52 efuse
X1040 a_638_27395.t45 a_14320_26417.t1 efuse
X1041 a_638_3764.t20 a_20810_624.t0 efuse
X1042 VSS.t135 BIT_SEL[30].t5 a_7830_62696.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1043 a_7830_46574.t1 a_638_43149.t38 efuse
X1044 a_7830_33029.t0 BIT_SEL[25].t4 VSS.t282 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1045 VSS.t396 BIT_SEL[52].t6 a_20810_5395.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1046 a_110_8311.t0 a_154_8223.t1 VSS.t328 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1047 a_638_58903.t64 a_1340_56291.t1 efuse
X1048 a_638_51026.t36 a_14320_50416.t1 efuse
X1049 a_1340_39641.t1 BIT_SEL[15].t6 VSS.t248 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1050 a_20810_20781.t1 a_638_19518.t19 efuse
X1051 a_110_61397.t0 a_154_61309.t1 VSS.t318 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1052 VSS.t569 a_110_49568.t4 OUT[6].t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1053 a_638_35272.t36 a_7830_34294.t1 efuse
X1054 a_20718_27712.t0 a_638_27395.t43 efuse
X1055 a_110_18956.t0 PRESET_N.t19 VDD VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1056 a_14320_21678.t1 a_638_19518.t39 efuse
X1057 a_638_43149.t55 a_14320_42171.t1 efuse
X1058 a_7830_2786.t0 BIT_SEL[19].t6 VSS.t157 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1059 VSS.t316 BIT_SEL[54].t6 a_20810_5924.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1060 a_20810_36535.t1 a_638_35272.t48 efuse
X1061 a_1340_12904.t1 a_638_11641.t42 efuse
X1062 a_7830_48783.t1 BIT_SEL[25].t5 VSS.t255 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1063 a_1340_48414.t1 BIT_SEL[11].t4 VSS.t419 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1064 a_20810_25152.t1 BIT_SEL[57].t7 VSS.t379 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1065 a_1248_4081.t1 a_638_3764.t64 efuse
X1066 a_20810_54451.t1 a_638_51026.t35 efuse
X1067 VSS.t67 BIT_SEL[32].t6 a_14228_43466.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1068 a_20718_43466.t0 a_638_43149.t34 efuse
X1069 a_110_34710.t0 PRESET_N.t20 VDD VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1070 a_14320_37432.t1 a_638_35272.t43 efuse
X1071 a_638_3764.t50 a_7830_2417.t1 efuse
X1072 VDD a_110_59829.t1 a_154_59741.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1073 VSS.t325 BIT_SEL[8].t6 a_1340_22046.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1074 a_110_3202.t0 PRESET_N.t21 VDD VDD pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1075 a_20810_25520.t0 BIT_SEL[55].t6 VSS.t270 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1076 a_1340_28658.t1 a_638_27395.t39 efuse
X1077 a_110_21116.t0 a_154_21028.t1 VSS.t48 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1078 a_638_11641.t59 a_14320_8133.t1 efuse
X1079 VSS.t274 BIT_SEL[34].t5 a_14320_44412.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1080 VDD a_110_28993.t1 a_154_28905.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1081 VDD.t121 COL_PROG_N[1].t3 a_638_11641.t21 VDD.t86 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X1082 VSS.t18 BIT_SEL[10].t4 a_1340_22414.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1083 VSS.t76 a_110_10183.t5 a_110_11079.t4 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1084 a_7830_5924.t1 a_638_3764.t41 efuse
X1085 a_638_3764.t46 a_14320_1152.t1 efuse
X1086 a_7830_16010.t1 BIT_SEL[31].t4 VSS.t287 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1087 VSS.t136 BIT_SEL[30].t6 a_7830_31188.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1088 a_638_19518.t33 a_1340_17275.t1 efuse
X1089 a_1340_44412.t1 a_638_43149.t20 efuse
X1090 a_1340_10663.t1 BIT_SEL[3].t6 VSS.t189 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1091 VDD a_110_44747.t1 a_154_44659.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1092 a_638_27395.t26 a_14320_23887.t0 efuse
X1093 a_14320_14537.t1 a_638_11641.t43 efuse
X1094 a_14320_33397.t0 BIT_SEL[39].t6 VSS.t390 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1095 a_7738_19835.t0 a_638_19518.t26 efuse
X1096 a_638_35272.t31 a_1340_33029.t1 efuse
X1097 a_7830_31764.t1 BIT_SEL[31].t5 VSS.t349 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1098 VSS.t512 BIT_SEL[20].t7 a_7830_29026.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1099 a_1340_11031.t0 BIT_SEL[1].t6 VSS.t147 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1100 a_14320_18540.t0 BIT_SEL[35].t6 VSS.t457 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1101 a_638_11641.t51 a_20810_9766.t1 efuse
X1102 a_7830_17275.t1 BIT_SEL[25].t6 VSS.t256 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1103 a_20810_52657.t0 a_638_51026.t37 efuse
X1104 a_20810_53554.t0 a_638_51026.t38 efuse
X1105 a_638_43149.t64 a_14320_39641.t1 efuse
X1106 VSS.t13 BIT_SEL[0].t7 a_1248_4081.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1107 a_14320_41802.t1 BIT_SEL[37].t6 VSS.t540 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1108 a_7738_35589.t0 a_638_35272.t33 efuse
X1109 a_14320_30291.t1 a_638_27395.t62 efuse
X1110 a_14320_5027.t0 a_638_3764.t53 efuse
X1111 VSS.t19 BIT_SEL[10].t5 a_1340_53922.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1112 a_110_37318.t0 a_154_37230.t1 VSS.t40 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1113 a_7830_17643.t1 BIT_SEL[23].t6 VSS.t435 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1114 a_638_19518.t62 a_20810_17275.t1 efuse
X1115 a_1340_42171.t1 BIT_SEL[3].t7 VSS.t478 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1116 VSS.t397 BIT_SEL[52].t7 a_20810_44780.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1117 VSS.t317 BIT_SEL[54].t7 a_20810_29555.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1118 a_638_27395.t21 a_20810_25520.t1 efuse
X1119 VSS.t529 a_110_26833.t7 a_110_25937.t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1120 a_14320_46045.t1 a_638_43149.t46 efuse
X1121 a_638_3764.t27 a_20810_256.t0 efuse
X1122 a_14320_9398.t1 BIT_SEL[41].t6 VSS.t201 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1123 a_638_11641.t33 a_7830_9029.t1 efuse
X1124 a_638_11641.t16 a_1340_8501.t0 efuse
X1125 a_1340_53922.t1 a_638_51026.t68 efuse
X1126 a_638_35272.t28 a_20810_33029.t1 efuse
X1127 a_110_32390.t0 a_154_32302.t1 VSS.t524 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1128 a_638_19518.t23 a_1340_18908.t0 efuse
X1129 a_14320_9766.t1 BIT_SEL[39].t7 VSS.t389 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1130 a_638_43149.t33 a_20810_41274.t1 efuse
X1131 VDD a_110_13239.t1 a_154_13151.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1132 a_638_35272.t19 a_1340_34662.t0 efuse
X1133 a_638_27395.t38 a_1340_24255.t1 efuse
X1134 a_638_27395.t47 a_7830_24783.t1 efuse
X1135 a_7830_3154.t1 BIT_SEL[17].t7 VSS.t180 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1136 a_7830_49151.t1 BIT_SEL[23].t7 VSS.t432 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1137 a_110_32838.t0 a_154_32750.t1 VSS.t513 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1138 a_20810_18908.t1 BIT_SEL[49].t7 VSS.t429 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1139 VSS.t329 a_110_58341.t7 a_110_57445.t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1140 VDD a_110_39110.t1 a_154_39022.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1141 a_638_19518.t58 COL_PROG_N[2].t2 VDD.t262 VDD.t2 pfet_06v0 ad=16.83p pd=77.38u as=9.945p ps=38.77u w=38.25u l=0.5u
X1142 a_14320_52657.t1 a_638_51026.t47 efuse
X1143 a_638_43149.t27 a_7830_40537.t1 efuse
X1144 VSS.t522 BIT_SEL[40].t7 a_14320_37800.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1145 a_14320_10294.t1 BIT_SEL[37].t7 VSS.t541 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1146 a_638_58903.t54 a_7830_55395.t0 efuse
X1147 a_638_43149.t12 a_1340_40009.t0 efuse
X1148 VSS.t503 BIT_SEL[48].t6 a_20718_11958.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1149 a_110_54864.t0 a_154_54776.t1 VSS.t224 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1150 a_7830_52289.t0 a_638_51026.t18 efuse
X1151 VSS.t233 BIT_SEL[12].t4 a_1340_30820.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1152 a_638_19518.t32 a_14320_17275.t0 efuse
X1153 a_638_19518.t59 COL_PROG_N[2].t3 VDD.t263 VDD.t76 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X1154 a_110_48592.t0 a_154_48504.t1 VSS.t182 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1155 a_638_11641.t50 a_1340_10294.t1 efuse
X1156 a_14320_60166.t0 a_638_58903.t34 efuse
X1157 VDD a_110_33814.t5 a_110_34710.t4 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1158 a_638_35272.t20 a_14320_33029.t0 efuse
X1159 a_20810_15434.t1 a_638_11641.t34 efuse
X1160 a_638_51026.t41 a_20810_48414.t1 efuse
X1161 a_638_51026.t64 a_20810_47518.t1 efuse
X1162 VSS.t234 BIT_SEL[12].t5 a_1340_46574.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1163 VDD a_110_30785.t1 a_154_30697.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1164 a_7830_22046.t1 a_638_19518.t45 efuse
X1165 VDD a_110_4690.t1 a_154_4602.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1166 VSS.t29 BIT_SEL[10].t6 a_1340_61799.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1167 VDD a_110_18956.t7 a_110_18060.t1 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1168 VDD a_110_49568.t5 a_110_50464.t3 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1169 a_638_51026.t61 COL_PROG_N[6].t2 VDD.t252 VDD.t2 pfet_06v0 ad=16.83p pd=77.38u as=9.945p ps=38.77u w=38.25u l=0.5u
X1170 a_7830_32132.t0 BIT_SEL[29].t6 VSS.t296 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1171 a_7830_7189.t1 a_638_3764.t68 efuse
X1172 a_638_27395.t51 a_1340_26048.t1 efuse
X1173 a_1340_47518.t0 BIT_SEL[15].t7 VSS.t77 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1174 VSS.t504 BIT_SEL[48].t7 a_20718_43466.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1175 VSS.t78 BIT_SEL[34].t6 a_14320_20781.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1176 VSS.t134 BIT_SEL[28].t7 a_7830_7189.t0 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1177 a_14320_8501.t0 BIT_SEL[45].t6 VSS.t508 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1178 VSS.t330 BIT_SEL[12].t6 a_1340_62328.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1179 a_7830_37800.t0 a_638_35272.t24 efuse
X1180 VSS.t603 BIT_SEL[2].t7 a_1340_5027.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1181 VDD a_110_53520.t1 a_154_53432.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1182 a_638_51026.t62 COL_PROG_N[6].t3 VDD.t253 VDD.t76 pfet_06v0 ad=9.945p pd=38.77u as=9.945p ps=38.77u w=38.25u l=0.5u
X1183 a_20810_31188.t1 a_638_27395.t28 efuse
X1184 VSS.t21 BIT_SEL[50].t7 a_20810_44412.t0 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1185 a_638_43149.t39 a_1340_41802.t1 efuse
X1186 a_638_3764.t43 a_14320_3154.t1 efuse
X1187 VSS.t137 BIT_SEL[30].t7 a_7830_7557.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1188 a_638_58903.t51 a_7830_57028.t0 efuse
X1189 a_1340_47886.t1 BIT_SEL[13].t6 VSS.t253 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1190 VDD a_110_40267.t1 a_154_40179.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1191 a_110_23356.t0 a_154_23268.t1 VSS.t420 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1192 a_1340_26048.t0 BIT_SEL[5].t5 VSS.t75 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1193 a_20810_46942.t1 a_638_43149.t47 efuse
X1194 VDD a_110_62293.t1 a_154_62205.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1195 a_14320_6292.t1 a_638_3764.t51 efuse
X1196 VDD a_110_7154.t1 a_154_7066.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1197 a_110_17084.t0 a_154_16996.t1 VSS.t190 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1198 a_20810_33397.t0 BIT_SEL[55].t7 VSS.t271 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1199 a_20810_14537.t1 a_638_11641.t61 efuse
X1200 a_20810_13801.t1 a_638_11641.t62 efuse
X1201 VDD a_110_46987.t1 a_154_46899.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1202 VSS.t448 BIT_SEL[36].t5 a_14320_36903.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1203 a_7830_256.t1 BIT_SEL[31].t6 VSS.t350 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1204 VSS.t79 BIT_SEL[34].t7 a_14320_52289.t1 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1205 a_14320_15434.t0 a_638_11641.t31 efuse
X1206 VSS.t331 BIT_SEL[12].t7 a_1340_15066.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1207 a_638_51026.t45 a_14320_48414.t1 efuse
X1208 VSS.t30 BIT_SEL[10].t7 a_1340_30291.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1209 VDD PRESET_N.t22 a_110_26833.t2 VDD pfet_06v0 ad=0.3172p pd=1.74u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1210 a_20810_18540.t0 BIT_SEL[51].t6 VSS.t343 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1211 VSS.t616 BIT_SEL[38].t7 a_14320_37432.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1212 a_20810_2786.t0 BIT_SEL[51].t7 VSS.t344 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1213 a_1340_2417.t0 BIT_SEL[5].t6 VSS.t619 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1214 VSS.t449 BIT_SEL[36].t6 a_14320_52657.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1215 VSS.t97 BIT_SEL[16].t6 a_7738_35589.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1216 a_7830_624.t0 BIT_SEL[29].t7 VSS.t297 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1217 a_20810_41802.t1 BIT_SEL[53].t6 VSS.t370 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1218 a_20810_30291.t1 a_638_27395.t49 efuse
X1219 VSS.t259 BIT_SEL[14].t6 a_1340_15434.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1220 a_7830_57925.t0 BIT_SEL[19].t7 VSS.t158 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1221 a_1340_57556.t0 BIT_SEL[5].t7 VSS.t620 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1222 a_20810_29555.t1 a_638_27395.t40 efuse
X1223 a_1340_21149.t1 a_638_19518.t47 efuse
X1224 a_638_3764.t47 a_20810_2417.t1 efuse
X1225 a_1340_15066.t1 a_638_11641.t55 efuse
X1226 a_638_58903.t47 a_14320_55763.t1 efuse
X1227 VDD a_110_56469.t1 a_154_56381.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1228 a_14320_40906.t0 BIT_SEL[41].t7 VSS.t202 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1229 VSS.t527 BIT_SEL[42].t7 a_14320_38168.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1230 VDD a_110_22012.t1 a_154_21924.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1231 VSS.t471 BIT_SEL[18].t7 a_7830_36535.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1232 a_14320_31188.t0 a_638_27395.t14 efuse
X1233 VSS.t558 a_110_3202.t7 a_110_2306.t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1234 a_1340_16378.t0 BIT_SEL[13].t7 VSS.t254 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1235 VSS.t365 BIT_SEL[6].t7 a_1340_61063.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1236 VSS.t98 BIT_SEL[16].t7 a_7738_51343.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1237 a_20810_46045.t1 a_638_43149.t36 efuse
X1238 a_14320_26417.t0 BIT_SEL[35].t7 VSS.t601 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1239 a_20810_45309.t0 a_638_43149.t23 efuse
X1240 VSS.t93 a_110_25937.t5 OUT[3].t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1241 a_638_11641.t56 a_7830_10663.t1 efuse
X1242 a_1340_36903.t1 a_638_35272.t63 efuse
X1243 a_14320_46942.t0 a_638_43149.t19 efuse
X1244 a_14320_256.t1 BIT_SEL[47].t7 VSS.t47 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1245 VSS.t105 BIT_SEL[24].t7 a_7830_6292.t1 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1246 VDD PRESET_N.t23 a_110_58341.t2 VDD pfet_06v0 ad=0.3172p pd=1.74u as=0.4575p ps=1.97u w=1.22u l=0.5u
X1247 a_1340_30820.t1 a_638_27395.t65 efuse
X1248 a_14320_26785.t0 BIT_SEL[33].t5 VSS.t590 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1249 a_20810_12904.t1 a_638_11641.t38 efuse
X1250 a_1340_54819.t1 a_638_51026.t53 efuse
X1251 a_1340_24783.t0 BIT_SEL[11].t5 VSS.t427 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1252 a_110_60501.t0 a_154_60413.t1 VSS.t159 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1253 a_14320_1152.t0 BIT_SEL[43].t7 VSS.t56 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1254 VDD a_110_15479.t1 a_154_15391.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1255 VSS.t258 BIT_SEL[14].t7 a_1340_46942.t1 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1256 a_638_27395.t41 a_7830_26417.t1 efuse
X1257 VSS.t68 BIT_SEL[32].t7 a_14228_19835.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1258 a_14320_624.t1 BIT_SEL[45].t7 VSS.t509 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1259 a_14320_13801.t1 a_638_11641.t60 efuse
X1260 a_638_51026.t52 a_7830_49679.t1 efuse
X1261 a_1340_46574.t1 a_638_43149.t54 efuse
X1262 a_110_28321.t0 a_154_28233.t1 VSS.t531 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1263 a_638_3764.t36 a_1340_256.t1 efuse
X1264 a_7830_62696.t0 a_638_58903.t25 efuse
X1265 a_638_51026.t40 a_7830_50416.t0 efuse
X1266 a_14320_42539.t0 BIT_SEL[33].t6 VSS.t591 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1267 a_1340_40537.t0 BIT_SEL[11].t6 VSS.t276 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1268 a_1340_50416.t1 BIT_SEL[1].t7 VSS.t327 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1269 VSS.t342 BIT_SEL[56].t7 a_20810_37800.t1 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1270 a_20810_28658.t1 a_638_27395.t22 efuse
X1271 VSS.t450 BIT_SEL[36].t7 a_14320_21149.t0 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1272 VDD.t46 COL_PROG_N[0].t3 a_638_3764.t5 VDD.t6 pfet_06v0 ad=9.945p pd=38.77u as=16.83p ps=77.38u w=38.25u l=0.5u
X1273 VDD a_110_38214.t1 a_154_38126.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1274 a_20810_10294.t0 BIT_SEL[53].t7 VSS.t371 VSS.t20 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1275 a_638_58903.t50 a_14320_57556.t1 efuse
X1276 VSS.t516 a_110_57445.t5 OUT[7].t1 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1277 a_638_43149.t49 a_7830_42171.t1 efuse
X1278 a_14320_29555.t1 a_638_27395.t64 efuse
X1279 a_110_53968.t0 a_154_53880.t1 VSS.t551 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1280 a_7830_8133.t0 BIT_SEL[31].t7 VSS.t351 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1281 a_14320_58293.t1 BIT_SEL[33].t7 VSS.t592 VSS.t41 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1282 a_20810_44412.t1 a_638_43149.t56 efuse
X1283 a_7830_56660.t1 BIT_SEL[25].t7 VSS.t257 VSS.t0 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1284 a_1340_56291.t0 BIT_SEL[11].t7 VSS.t436 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1285 a_14320_6660.t0 a_638_3764.t31 efuse
X1286 a_638_19518.t24 SENSE.t7 a_110_18956.t5 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1287 a_110_47696.t0 a_154_47608.t1 VSS.t528 VSS.t31 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1288 a_14320_45309.t1 a_638_43149.t22 efuse
X1289 a_638_11641.t37 a_1340_9398.t1 efuse
X1290 a_1340_53186.t1 a_638_51026.t34 efuse
X1291 VSS.t326 BIT_SEL[8].t7 a_1340_29923.t0 VSS.t5 nfet_06v0 ad=13.42p pd=61.88u as=13.42p ps=61.88u w=30.5u l=0.6u
X1292 a_638_19518.t64 a_1340_16906.t1 efuse
X1293 a_7738_11958.t0 a_638_11641.t40 efuse
X1294 a_7830_61799.t1 a_638_58903.t66 efuse
X1295 VDD a_110_36870.t1 a_154_36782.t0 VDD pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
R0 a_1340_61431.t0 a_1340_61431.t1 5.92611
R1 a_638_58903.t0 a_638_58903.n0 7.71211
R2 a_638_58903.n1 a_638_58903.t18 7.71211
R3 a_638_58903.n2 a_638_58903.t57 7.71211
R4 a_638_58903.n3 a_638_58903.t27 7.71211
R5 a_638_58903.n4 a_638_58903.t59 7.71211
R6 a_638_58903.n5 a_638_58903.t29 7.71211
R7 a_638_58903.n6 a_638_58903.t24 7.71211
R8 a_638_58903.n7 a_638_58903.t60 7.71211
R9 a_638_58903.n8 a_638_58903.t16 7.71211
R10 a_638_58903.n9 a_638_58903.t63 7.71211
R11 a_638_58903.n10 a_638_58903.t45 7.71211
R12 a_638_58903.n11 a_638_58903.t11 7.71211
R13 a_638_58903.n12 a_638_58903.t56 7.71211
R14 a_638_58903.n13 a_638_58903.t66 7.71211
R15 a_638_58903.n14 a_638_58903.t48 7.71211
R16 a_638_58903.n15 a_638_58903.t25 7.71211
R17 a_638_58903.n16 a_638_58903.t55 7.71211
R18 a_638_58903.n17 a_638_58903.t34 7.71211
R19 a_638_58903.n18 a_638_58903.t68 7.71211
R20 a_638_58903.n19 a_638_58903.t43 7.71211
R21 a_638_58903.n20 a_638_58903.t12 7.71211
R22 a_638_58903.n21 a_638_58903.t33 7.71211
R23 a_638_58903.n22 a_638_58903.t61 7.71211
R24 a_638_58903.n23 a_638_58903.t41 7.71211
R25 a_638_58903.n24 a_638_58903.t49 7.71211
R26 a_638_58903.n25 a_638_58903.t22 7.71211
R27 a_638_58903.n26 a_638_58903.t3 7.71211
R28 a_638_58903.n27 a_638_58903.t67 7.71211
R29 a_638_58903.n28 a_638_58903.t62 7.71211
R30 a_638_58903.n29 a_638_58903.t40 7.71211
R31 a_638_58903.n30 a_638_58903.t14 7.71211
R32 a_638_58903.n31 a_638_58903.t35 7.71211
R33 a_638_58903.n2 a_638_58903.n1 0.427167
R34 a_638_58903.n3 a_638_58903.n2 0.427167
R35 a_638_58903.n4 a_638_58903.n3 0.427167
R36 a_638_58903.n5 a_638_58903.n4 0.427167
R37 a_638_58903.n6 a_638_58903.n5 0.427167
R38 a_638_58903.n7 a_638_58903.n6 0.427167
R39 a_638_58903.n8 a_638_58903.n7 0.427167
R40 a_638_58903.n9 a_638_58903.n8 0.619389
R41 a_638_58903.n10 a_638_58903.n9 0.427167
R42 a_638_58903.n11 a_638_58903.n10 0.427167
R43 a_638_58903.n0 a_638_58903.n11 0.427167
R44 a_638_58903.n0 a_638_58903.n12 0.427167
R45 a_638_58903.n12 a_638_58903.n13 0.427167
R46 a_638_58903.n13 a_638_58903.n14 0.427167
R47 a_638_58903.n14 a_638_58903.n15 0.427167
R48 a_638_58903.n15 a_638_58903.n16 0.619389
R49 a_638_58903.n16 a_638_58903.n17 0.427167
R50 a_638_58903.n17 a_638_58903.n18 0.427167
R51 a_638_58903.n18 a_638_58903.n19 0.427167
R52 a_638_58903.n19 a_638_58903.n20 0.427167
R53 a_638_58903.n20 a_638_58903.n21 0.427167
R54 a_638_58903.n21 a_638_58903.n22 0.427167
R55 a_638_58903.n22 a_638_58903.n23 0.427167
R56 a_638_58903.n23 a_638_58903.n24 0.619389
R57 a_638_58903.n24 a_638_58903.n25 0.427167
R58 a_638_58903.n25 a_638_58903.n26 0.427167
R59 a_638_58903.n26 a_638_58903.n27 0.427167
R60 a_638_58903.n27 a_638_58903.n28 0.427167
R61 a_638_58903.n28 a_638_58903.n29 0.427167
R62 a_638_58903.n29 a_638_58903.n30 0.427167
R63 a_638_58903.n30 a_638_58903.n31 0.427167
R64 a_638_58903.n31 a_638_58903.n34 0.548278
R65 a_638_58903.n34 a_638_58903.n70 0.227167
R66 a_638_58903.n1 a_638_58903.n32 0.466493
R67 a_638_58903.n36 a_638_58903.t53 7.71211
R68 a_638_58903.n37 a_638_58903.t19 7.71211
R69 a_638_58903.n38 a_638_58903.t37 7.71211
R70 a_638_58903.n39 a_638_58903.t1 7.71211
R71 a_638_58903.n40 a_638_58903.t52 7.71211
R72 a_638_58903.n41 a_638_58903.t64 7.71211
R73 a_638_58903.n42 a_638_58903.t26 7.71211
R74 a_638_58903.n43 a_638_58903.t13 7.71211
R75 a_638_58903.n44 a_638_58903.t17 7.71211
R76 a_638_58903.n45 a_638_58903.t44 7.71211
R77 a_638_58903.n46 a_638_58903.t15 7.71211
R78 a_638_58903.n47 a_638_58903.t51 7.71211
R79 a_638_58903.n48 a_638_58903.t2 7.71211
R80 a_638_58903.n49 a_638_58903.t42 7.71211
R81 a_638_58903.n50 a_638_58903.t6 7.71211
R82 a_638_58903.n51 a_638_58903.t54 7.71211
R83 a_638_58903.n52 a_638_58903.t31 7.71211
R84 a_638_58903.n53 a_638_58903.t28 7.71211
R85 a_638_58903.n54 a_638_58903.t50 7.71211
R86 a_638_58903.n55 a_638_58903.t65 7.71211
R87 a_638_58903.n56 a_638_58903.t46 7.71211
R88 a_638_58903.n57 a_638_58903.t21 7.71211
R89 a_638_58903.n58 a_638_58903.t47 7.71211
R90 a_638_58903.n59 a_638_58903.t20 7.71211
R91 a_638_58903.n60 a_638_58903.t36 7.71211
R92 a_638_58903.n61 a_638_58903.t38 7.71211
R93 a_638_58903.n62 a_638_58903.t4 7.71211
R94 a_638_58903.n63 a_638_58903.t39 7.71211
R95 a_638_58903.n64 a_638_58903.t23 7.71211
R96 a_638_58903.n65 a_638_58903.t5 7.71211
R97 a_638_58903.n66 a_638_58903.t32 7.71211
R98 a_638_58903.n67 a_638_58903.t58 7.71211
R99 a_638_58903.n32 a_638_58903.n36 0.69448
R100 a_638_58903.n36 a_638_58903.n37 0.427167
R101 a_638_58903.n37 a_638_58903.n38 0.427167
R102 a_638_58903.n38 a_638_58903.n39 0.427167
R103 a_638_58903.n39 a_638_58903.n40 0.427167
R104 a_638_58903.n40 a_638_58903.n41 0.427167
R105 a_638_58903.n41 a_638_58903.n42 0.427167
R106 a_638_58903.n42 a_638_58903.n43 0.427167
R107 a_638_58903.n43 a_638_58903.n44 0.619389
R108 a_638_58903.n44 a_638_58903.n45 0.427167
R109 a_638_58903.n45 a_638_58903.n46 0.427167
R110 a_638_58903.n46 a_638_58903.n47 0.427167
R111 a_638_58903.n47 a_638_58903.n48 0.427167
R112 a_638_58903.n48 a_638_58903.n49 0.427167
R113 a_638_58903.n49 a_638_58903.n50 0.427167
R114 a_638_58903.n50 a_638_58903.n51 0.427167
R115 a_638_58903.n51 a_638_58903.n52 0.619389
R116 a_638_58903.n52 a_638_58903.n53 0.427167
R117 a_638_58903.n53 a_638_58903.n54 0.427167
R118 a_638_58903.n54 a_638_58903.n55 0.427167
R119 a_638_58903.n55 a_638_58903.n56 0.427167
R120 a_638_58903.n56 a_638_58903.n57 0.427167
R121 a_638_58903.n57 a_638_58903.n58 0.427167
R122 a_638_58903.n58 a_638_58903.n59 0.427167
R123 a_638_58903.n59 a_638_58903.n60 0.619389
R124 a_638_58903.n60 a_638_58903.n61 0.427167
R125 a_638_58903.n61 a_638_58903.n62 0.427167
R126 a_638_58903.n62 a_638_58903.n63 0.427167
R127 a_638_58903.n63 a_638_58903.n64 0.427167
R128 a_638_58903.n64 a_638_58903.n65 0.427167
R129 a_638_58903.n65 a_638_58903.n66 0.427167
R130 a_638_58903.n66 a_638_58903.n67 0.427167
R131 a_638_58903.n35 a_638_58903.n67 0.334944
R132 a_638_58903.n35 a_638_58903.n71 0.227167
R133 a_638_58903.n70 a_638_58903.n72 4.96756
R134 a_638_58903.n72 a_638_58903.n71 4.83019
R135 a_638_58903.n72 a_638_58903.t9 0.113082
R136 a_638_58903.n69 a_638_58903.n68 0.0655
R137 a_638_58903.n69 a_638_58903.n71 4.60509
R138 a_638_58903.n70 a_638_58903.n69 4.74618
R139 a_638_58903.n68 a_638_58903.t10 0.0480817
R140 a_638_58903.n68 a_638_58903.t7 0.0480817
R141 a_638_58903.n33 a_638_58903.n35 4.60509
R142 a_638_58903.n34 a_638_58903.n33 4.74618
R143 a_638_58903.n33 a_638_58903.t8 0.113082
R144 a_638_58903.n32 a_638_58903.t30 9.85476
R145 a_7830_61063.t0 a_7830_61063.t1 6.38524
R146 BIT_SEL[50] BIT_SEL[50].n0 1.95318
R147 BIT_SEL[50] BIT_SEL[50].n0 10.6751
R148 BIT_SEL[50] BIT_SEL[50].n1 1.95318
R149 BIT_SEL[50].n1 BIT_SEL[50] 10.6751
R150 BIT_SEL[50] BIT_SEL[50].n2 1.95318
R151 BIT_SEL[50].n2 BIT_SEL[50] 10.6751
R152 BIT_SEL[50] BIT_SEL[50].n3 1.95318
R153 BIT_SEL[50].n3 BIT_SEL[50] 10.6751
R154 BIT_SEL[50] BIT_SEL[50].n4 1.95318
R155 BIT_SEL[50].n4 BIT_SEL[50] 10.6751
R156 BIT_SEL[50] BIT_SEL[50].n5 1.95318
R157 BIT_SEL[50].n5 BIT_SEL[50] 10.6751
R158 BIT_SEL[50] BIT_SEL[50].n6 1.95318
R159 BIT_SEL[50].n6 BIT_SEL[50] 10.6751
R160 BIT_SEL[50].t3 BIT_SEL[50] 117.727
R161 BIT_SEL[50].t1 BIT_SEL[50].n6 115.775
R162 BIT_SEL[50].t7 BIT_SEL[50].n5 115.775
R163 BIT_SEL[50].t6 BIT_SEL[50].n4 115.775
R164 BIT_SEL[50].t5 BIT_SEL[50].n3 115.775
R165 BIT_SEL[50].t0 BIT_SEL[50].n2 115.775
R166 BIT_SEL[50].n1 BIT_SEL[50].t2 115.775
R167 BIT_SEL[50].n0 BIT_SEL[50].t4 115.775
R168 a_20810_20781.t0 a_20810_20781.t1 8.02269
R169 VSS.n0 VSS.n1 4.5005
R170 VSS.n3 VSS.n2 0.0732424
R171 VSS.n1 VSS.n3 2.21488
R172 VSS.n6 VSS.n5 0.0732424
R173 VSS.n1 VSS.n6 2.21488
R174 VSS.n15 VSS.n16 4.5005
R175 VSS.n18 VSS.n17 0.0732424
R176 VSS.n16 VSS.n18 2.21488
R177 VSS.n21 VSS.n20 0.0732424
R178 VSS.n16 VSS.n21 2.21488
R179 VSS.n30 VSS.n31 4.5005
R180 VSS.n32 VSS.n33 0.0732424
R181 VSS.n33 VSS.n31 2.21488
R182 VSS.n2098 VSS.n31 2.21488
R183 VSS.n2097 VSS.n2098 4.57324
R184 VSS.n36 VSS.n37 4.5005
R185 VSS.n39 VSS.n38 0.0732424
R186 VSS.n37 VSS.n39 2.21488
R187 VSS.n42 VSS.n41 0.0732424
R188 VSS.n37 VSS.n42 2.21488
R189 VSS.n51 VSS.n52 4.5005
R190 VSS.n54 VSS.n53 0.0732424
R191 VSS.n52 VSS.n54 2.21488
R192 VSS.n57 VSS.n56 0.0732424
R193 VSS.n52 VSS.n57 2.21488
R194 VSS.n66 VSS.n67 4.5005
R195 VSS.n69 VSS.n68 0.0732424
R196 VSS.n67 VSS.n69 2.21488
R197 VSS.n72 VSS.n71 0.0732424
R198 VSS.n67 VSS.n72 2.21488
R199 VSS.n81 VSS.n82 4.5005
R200 VSS.n83 VSS.n84 0.0732424
R201 VSS.n84 VSS.n82 2.21488
R202 VSS.n2107 VSS.n82 2.21488
R203 VSS.n2106 VSS.n2107 4.57324
R204 VSS.n87 VSS.n88 4.5005
R205 VSS.n90 VSS.n89 0.0732424
R206 VSS.n88 VSS.n90 2.21488
R207 VSS.n93 VSS.n92 0.0732424
R208 VSS.n88 VSS.n93 2.21488
R209 VSS.n102 VSS.n103 4.5005
R210 VSS.n105 VSS.n104 0.0732424
R211 VSS.n103 VSS.n105 2.21488
R212 VSS.n108 VSS.n107 0.0732424
R213 VSS.n103 VSS.n108 2.21488
R214 VSS.n117 VSS.n118 4.5005
R215 VSS.n120 VSS.n119 0.0732424
R216 VSS.n118 VSS.n120 2.21488
R217 VSS.n123 VSS.n122 0.0732424
R218 VSS.n118 VSS.n123 2.21488
R219 VSS.n132 VSS.n133 4.5005
R220 VSS.n135 VSS.n134 0.0732424
R221 VSS.n133 VSS.n135 2.21488
R222 VSS.n138 VSS.n137 0.0732424
R223 VSS.n133 VSS.n138 2.21488
R224 VSS.n147 VSS.n148 4.5005
R225 VSS.n150 VSS.n149 0.0732424
R226 VSS.n148 VSS.n150 2.21488
R227 VSS.n153 VSS.n152 0.0732424
R228 VSS.n148 VSS.n153 2.21488
R229 VSS.n162 VSS.n163 4.5005
R230 VSS.n165 VSS.n164 0.0732424
R231 VSS.n163 VSS.n165 2.21488
R232 VSS.n168 VSS.n167 0.0732424
R233 VSS.n163 VSS.n168 2.21488
R234 VSS.n177 VSS.n178 4.5005
R235 VSS.n179 VSS.n180 0.0732424
R236 VSS.n180 VSS.n178 2.21488
R237 VSS.n2117 VSS.n178 2.21488
R238 VSS.n2116 VSS.n2117 4.57324
R239 VSS.n183 VSS.n184 4.5005
R240 VSS.n186 VSS.n185 0.0732424
R241 VSS.n184 VSS.n186 2.21488
R242 VSS.n189 VSS.n188 0.0732424
R243 VSS.n184 VSS.n189 2.21488
R244 VSS.n198 VSS.n199 4.5005
R245 VSS.n201 VSS.n200 0.0732424
R246 VSS.n199 VSS.n201 2.21488
R247 VSS.n204 VSS.n203 0.0732424
R248 VSS.n199 VSS.n204 2.21488
R249 VSS.n213 VSS.n214 4.5005
R250 VSS.n216 VSS.n215 0.0732424
R251 VSS.n214 VSS.n216 2.21488
R252 VSS.n219 VSS.n218 0.0732424
R253 VSS.n214 VSS.n219 2.21488
R254 VSS.n228 VSS.n229 4.5005
R255 VSS.n230 VSS.n231 0.0732424
R256 VSS.n231 VSS.n229 2.21488
R257 VSS.n2126 VSS.n229 2.21488
R258 VSS.n2125 VSS.n2126 4.57324
R259 VSS.n234 VSS.n235 4.5005
R260 VSS.n237 VSS.n236 0.0732424
R261 VSS.n235 VSS.n237 2.21488
R262 VSS.n240 VSS.n239 0.0732424
R263 VSS.n235 VSS.n240 2.21488
R264 VSS.n249 VSS.n250 4.5005
R265 VSS.n252 VSS.n251 0.0732424
R266 VSS.n250 VSS.n252 2.21488
R267 VSS.n255 VSS.n254 0.0732424
R268 VSS.n250 VSS.n255 2.21488
R269 VSS.n264 VSS.n265 4.5005
R270 VSS.n267 VSS.n266 0.0732424
R271 VSS.n265 VSS.n267 2.21488
R272 VSS.n270 VSS.n269 0.0732424
R273 VSS.n265 VSS.n270 2.21488
R274 VSS.n279 VSS.n280 4.5005
R275 VSS.n282 VSS.n281 0.0732424
R276 VSS.n280 VSS.n282 2.21488
R277 VSS.n285 VSS.n284 0.0732424
R278 VSS.n280 VSS.n285 2.21488
R279 VSS.n294 VSS.n295 4.5005
R280 VSS.n296 VSS.n297 0.0732424
R281 VSS.n297 VSS.n295 2.21488
R282 VSS.n2135 VSS.n295 2.21488
R283 VSS.n2134 VSS.n2135 4.57324
R284 VSS.n300 VSS.n301 4.5005
R285 VSS.n303 VSS.n302 0.0732424
R286 VSS.n301 VSS.n303 2.21488
R287 VSS.n306 VSS.n305 0.0732424
R288 VSS.n301 VSS.n306 2.21488
R289 VSS.n315 VSS.n316 4.5005
R290 VSS.n318 VSS.n317 0.0732424
R291 VSS.n316 VSS.n318 2.21488
R292 VSS.n321 VSS.n320 0.0732424
R293 VSS.n316 VSS.n321 2.21488
R294 VSS.n330 VSS.n331 4.5005
R295 VSS.n333 VSS.n332 0.0732424
R296 VSS.n331 VSS.n333 2.21488
R297 VSS.n336 VSS.n335 0.0732424
R298 VSS.n331 VSS.n336 2.21488
R299 VSS.n345 VSS.n346 4.5005
R300 VSS.n347 VSS.n348 0.0732424
R301 VSS.n348 VSS.n346 2.21488
R302 VSS.n2144 VSS.n346 2.21488
R303 VSS.n2143 VSS.n2144 4.57324
R304 VSS.n351 VSS.n352 4.5005
R305 VSS.n354 VSS.n353 0.0732424
R306 VSS.n352 VSS.n354 2.21488
R307 VSS.n357 VSS.n356 0.0732424
R308 VSS.n352 VSS.n357 2.21488
R309 VSS.n366 VSS.n367 4.5005
R310 VSS.n369 VSS.n368 0.0732424
R311 VSS.n367 VSS.n369 2.21488
R312 VSS.n372 VSS.n371 0.0732424
R313 VSS.n367 VSS.n372 2.21488
R314 VSS.n381 VSS.n382 4.5005
R315 VSS.n384 VSS.n383 0.0732424
R316 VSS.n382 VSS.n384 2.21488
R317 VSS.n387 VSS.n386 0.0732424
R318 VSS.n382 VSS.n387 2.21488
R319 VSS.n396 VSS.n397 4.5005
R320 VSS.n399 VSS.n398 0.0732424
R321 VSS.n397 VSS.n399 2.21488
R322 VSS.n402 VSS.n401 0.0732424
R323 VSS.n397 VSS.n402 2.21488
R324 VSS.n411 VSS.n412 4.5005
R325 VSS.n414 VSS.n413 0.0732424
R326 VSS.n412 VSS.n414 2.21488
R327 VSS.n417 VSS.n416 0.0732424
R328 VSS.n412 VSS.n417 2.21488
R329 VSS.n426 VSS.n427 4.5005
R330 VSS.n429 VSS.n428 0.0732424
R331 VSS.n427 VSS.n429 2.21488
R332 VSS.n432 VSS.n431 0.0732424
R333 VSS.n427 VSS.n432 2.21488
R334 VSS.n441 VSS.n442 4.5005
R335 VSS.n443 VSS.n444 0.0732424
R336 VSS.n444 VSS.n442 2.21488
R337 VSS.n2153 VSS.n442 2.21488
R338 VSS.n2152 VSS.n2153 4.57324
R339 VSS.n447 VSS.n448 4.5005
R340 VSS.n450 VSS.n449 0.0732424
R341 VSS.n448 VSS.n450 2.21488
R342 VSS.n453 VSS.n452 0.0732424
R343 VSS.n448 VSS.n453 2.21488
R344 VSS.n462 VSS.n463 4.5005
R345 VSS.n465 VSS.n464 0.0732424
R346 VSS.n463 VSS.n465 2.21488
R347 VSS.n468 VSS.n467 0.0732424
R348 VSS.n463 VSS.n468 2.21488
R349 VSS.n477 VSS.n478 4.5005
R350 VSS.n480 VSS.n479 0.0732424
R351 VSS.n478 VSS.n480 2.21488
R352 VSS.n483 VSS.n482 0.0732424
R353 VSS.n478 VSS.n483 2.21488
R354 VSS.n492 VSS.n493 4.5005
R355 VSS.n494 VSS.n495 0.0732424
R356 VSS.n495 VSS.n493 2.21488
R357 VSS.n2162 VSS.n493 2.21488
R358 VSS.n2161 VSS.n2162 4.57324
R359 VSS.n498 VSS.n499 4.5005
R360 VSS.n501 VSS.n500 0.0732424
R361 VSS.n499 VSS.n501 2.21488
R362 VSS.n504 VSS.n503 0.0732424
R363 VSS.n499 VSS.n504 2.21488
R364 VSS.n513 VSS.n514 4.5005
R365 VSS.n516 VSS.n515 0.0732424
R366 VSS.n514 VSS.n516 2.21488
R367 VSS.n519 VSS.n518 0.0732424
R368 VSS.n514 VSS.n519 2.21488
R369 VSS.n528 VSS.n529 4.5005
R370 VSS.n531 VSS.n530 0.0732424
R371 VSS.n529 VSS.n531 2.21488
R372 VSS.n534 VSS.n533 0.0732424
R373 VSS.n529 VSS.n534 2.21488
R374 VSS.n543 VSS.n544 4.5005
R375 VSS.n546 VSS.n545 0.0732424
R376 VSS.n544 VSS.n546 2.21488
R377 VSS.n549 VSS.n548 0.0732424
R378 VSS.n544 VSS.n549 2.21488
R379 VSS.n558 VSS.n559 4.5005
R380 VSS.n560 VSS.n561 0.0732424
R381 VSS.n561 VSS.n559 2.21488
R382 VSS.n2171 VSS.n559 2.21488
R383 VSS.n2170 VSS.n2171 4.57324
R384 VSS.n564 VSS.n565 4.5005
R385 VSS.n567 VSS.n566 0.0732424
R386 VSS.n565 VSS.n567 2.21488
R387 VSS.n570 VSS.n569 0.0732424
R388 VSS.n565 VSS.n570 2.21488
R389 VSS.n579 VSS.n580 4.5005
R390 VSS.n582 VSS.n581 0.0732424
R391 VSS.n580 VSS.n582 2.21488
R392 VSS.n585 VSS.n584 0.0732424
R393 VSS.n580 VSS.n585 2.21488
R394 VSS.n594 VSS.n595 4.5005
R395 VSS.n597 VSS.n596 0.0732424
R396 VSS.n595 VSS.n597 2.21488
R397 VSS.n600 VSS.n599 0.0732424
R398 VSS.n595 VSS.n600 2.21488
R399 VSS.n609 VSS.n610 4.5005
R400 VSS.n611 VSS.n612 0.0732424
R401 VSS.n612 VSS.n610 2.21488
R402 VSS.n2180 VSS.n610 2.21488
R403 VSS.n2179 VSS.n2180 4.57324
R404 VSS.n615 VSS.n616 4.5005
R405 VSS.n618 VSS.n617 0.0732424
R406 VSS.n616 VSS.n618 2.21488
R407 VSS.n621 VSS.n620 0.0732424
R408 VSS.n616 VSS.n621 2.21488
R409 VSS.n630 VSS.n631 4.5005
R410 VSS.n633 VSS.n632 0.0732424
R411 VSS.n631 VSS.n633 2.21488
R412 VSS.n636 VSS.n635 0.0732424
R413 VSS.n631 VSS.n636 2.21488
R414 VSS.n645 VSS.n646 4.5005
R415 VSS.n648 VSS.n647 0.0732424
R416 VSS.n646 VSS.n648 2.21488
R417 VSS.n651 VSS.n650 0.0732424
R418 VSS.n646 VSS.n651 2.21488
R419 VSS.n660 VSS.n661 4.5005
R420 VSS.n663 VSS.n662 0.0732424
R421 VSS.n661 VSS.n663 2.21488
R422 VSS.n666 VSS.n665 0.0732424
R423 VSS.n661 VSS.n666 2.21488
R424 VSS.n675 VSS.n676 4.5005
R425 VSS.n678 VSS.n677 0.0732424
R426 VSS.n676 VSS.n678 2.21488
R427 VSS.n681 VSS.n680 0.0732424
R428 VSS.n676 VSS.n681 2.21488
R429 VSS.n690 VSS.n691 4.5005
R430 VSS.n693 VSS.n692 0.0732424
R431 VSS.n691 VSS.n693 2.21488
R432 VSS.n696 VSS.n695 0.0732424
R433 VSS.n691 VSS.n696 2.21488
R434 VSS.n705 VSS.n706 4.5005
R435 VSS.n707 VSS.n708 0.0732424
R436 VSS.n708 VSS.n706 2.21488
R437 VSS.n2189 VSS.n706 2.21488
R438 VSS.n2188 VSS.n2189 4.57324
R439 VSS.n711 VSS.n712 4.5005
R440 VSS.n714 VSS.n713 0.0732424
R441 VSS.n712 VSS.n714 2.21488
R442 VSS.n717 VSS.n716 0.0732424
R443 VSS.n712 VSS.n717 2.21488
R444 VSS.n726 VSS.n727 4.5005
R445 VSS.n729 VSS.n728 0.0732424
R446 VSS.n727 VSS.n729 2.21488
R447 VSS.n732 VSS.n731 0.0732424
R448 VSS.n727 VSS.n732 2.21488
R449 VSS.n741 VSS.n742 4.5005
R450 VSS.n744 VSS.n743 0.0732424
R451 VSS.n742 VSS.n744 2.21488
R452 VSS.n747 VSS.n746 0.0732424
R453 VSS.n742 VSS.n747 2.21488
R454 VSS.n756 VSS.n757 4.5005
R455 VSS.n758 VSS.n759 0.0732424
R456 VSS.n759 VSS.n757 2.21488
R457 VSS.n2198 VSS.n757 2.21488
R458 VSS.n2197 VSS.n2198 4.57324
R459 VSS.n762 VSS.n763 4.5005
R460 VSS.n765 VSS.n764 0.0732424
R461 VSS.n763 VSS.n765 2.21488
R462 VSS.n768 VSS.n767 0.0732424
R463 VSS.n763 VSS.n768 2.21488
R464 VSS.n777 VSS.n778 4.5005
R465 VSS.n780 VSS.n779 0.0732424
R466 VSS.n778 VSS.n780 2.21488
R467 VSS.n783 VSS.n782 0.0732424
R468 VSS.n778 VSS.n783 2.21488
R469 VSS.n792 VSS.n793 4.5005
R470 VSS.n795 VSS.n794 0.0732424
R471 VSS.n793 VSS.n795 2.21488
R472 VSS.n798 VSS.n797 0.0732424
R473 VSS.n793 VSS.n798 2.21488
R474 VSS.n807 VSS.n808 4.5005
R475 VSS.n810 VSS.n809 0.0732424
R476 VSS.n808 VSS.n810 2.21488
R477 VSS.n813 VSS.n812 0.0732424
R478 VSS.n808 VSS.n813 2.21488
R479 VSS.n822 VSS.n823 4.5005
R480 VSS.n824 VSS.n825 0.0732424
R481 VSS.n825 VSS.n823 2.21488
R482 VSS.n2207 VSS.n823 2.21488
R483 VSS.n2206 VSS.n2207 4.57324
R484 VSS.n828 VSS.n829 4.5005
R485 VSS.n831 VSS.n830 0.0732424
R486 VSS.n829 VSS.n831 2.21488
R487 VSS.n834 VSS.n833 0.0732424
R488 VSS.n829 VSS.n834 2.21488
R489 VSS.n843 VSS.n844 4.5005
R490 VSS.n846 VSS.n845 0.0732424
R491 VSS.n844 VSS.n846 2.21488
R492 VSS.n849 VSS.n848 0.0732424
R493 VSS.n844 VSS.n849 2.21488
R494 VSS.n858 VSS.n859 4.5005
R495 VSS.n861 VSS.n860 0.0732424
R496 VSS.n859 VSS.n861 2.21488
R497 VSS.n864 VSS.n863 0.0732424
R498 VSS.n859 VSS.n864 2.21488
R499 VSS.n873 VSS.n874 4.5005
R500 VSS.n875 VSS.n876 0.0732424
R501 VSS.n876 VSS.n874 2.21488
R502 VSS.n2216 VSS.n874 2.21488
R503 VSS.n2215 VSS.n2216 4.57324
R504 VSS.n879 VSS.n880 4.5005
R505 VSS.n882 VSS.n881 0.0732424
R506 VSS.n880 VSS.n882 2.21488
R507 VSS.n885 VSS.n884 0.0732424
R508 VSS.n880 VSS.n885 2.21488
R509 VSS.n894 VSS.n895 4.5005
R510 VSS.n897 VSS.n896 0.0732424
R511 VSS.n895 VSS.n897 2.21488
R512 VSS.n900 VSS.n899 0.0732424
R513 VSS.n895 VSS.n900 2.21488
R514 VSS.n909 VSS.n910 4.5005
R515 VSS.n912 VSS.n911 0.0732424
R516 VSS.n910 VSS.n912 2.21488
R517 VSS.n915 VSS.n914 0.0732424
R518 VSS.n910 VSS.n915 2.21488
R519 VSS.n924 VSS.n925 4.5005
R520 VSS.n927 VSS.n926 0.0732424
R521 VSS.n925 VSS.n927 2.21488
R522 VSS.n930 VSS.n929 0.0732424
R523 VSS.n925 VSS.n930 2.21488
R524 VSS.n939 VSS.n940 4.5005
R525 VSS.n942 VSS.n941 0.0732424
R526 VSS.n940 VSS.n942 2.21488
R527 VSS.n945 VSS.n944 0.0732424
R528 VSS.n940 VSS.n945 2.21488
R529 VSS.n954 VSS.n955 4.5005
R530 VSS.n957 VSS.n956 0.0732424
R531 VSS.n955 VSS.n957 2.21488
R532 VSS.n960 VSS.n959 0.0732424
R533 VSS.n955 VSS.n960 2.21488
R534 VSS.n969 VSS.n970 4.5005
R535 VSS.n971 VSS.n972 0.0732424
R536 VSS.n972 VSS.n970 2.21488
R537 VSS.n2225 VSS.n970 2.21488
R538 VSS.n2224 VSS.n2225 4.57324
R539 VSS.n975 VSS.n976 4.5005
R540 VSS.n978 VSS.n977 0.0732424
R541 VSS.n976 VSS.n978 2.21488
R542 VSS.n981 VSS.n980 0.0732424
R543 VSS.n976 VSS.n981 2.21488
R544 VSS.n990 VSS.n991 4.5005
R545 VSS.n993 VSS.n992 0.0732424
R546 VSS.n991 VSS.n993 2.21488
R547 VSS.n996 VSS.n995 0.0732424
R548 VSS.n991 VSS.n996 2.21488
R549 VSS.n1005 VSS.n1006 4.5005
R550 VSS.n1008 VSS.n1007 0.0732424
R551 VSS.n1006 VSS.n1008 2.21488
R552 VSS.n1011 VSS.n1010 0.0732424
R553 VSS.n1006 VSS.n1011 2.21488
R554 VSS.n1020 VSS.n1021 4.5005
R555 VSS.n1022 VSS.n1023 0.0732424
R556 VSS.n1023 VSS.n1021 2.21488
R557 VSS.n2234 VSS.n1021 2.21488
R558 VSS.n2233 VSS.n2234 4.57324
R559 VSS.n1026 VSS.n1027 4.5005
R560 VSS.n1029 VSS.n1028 0.0732424
R561 VSS.n1027 VSS.n1029 2.21488
R562 VSS.n1032 VSS.n1031 0.0732424
R563 VSS.n1027 VSS.n1032 2.21488
R564 VSS.n1041 VSS.n1042 4.5005
R565 VSS.n1044 VSS.n1043 0.0732424
R566 VSS.n1042 VSS.n1044 2.21488
R567 VSS.n1047 VSS.n1046 0.0732424
R568 VSS.n1042 VSS.n1047 2.21488
R569 VSS.n1056 VSS.n1057 4.5005
R570 VSS.n1059 VSS.n1058 0.0732424
R571 VSS.n1057 VSS.n1059 2.21488
R572 VSS.n1062 VSS.n1061 0.0732424
R573 VSS.n1057 VSS.n1062 2.21488
R574 VSS.n1071 VSS.n1072 4.5005
R575 VSS.n1074 VSS.n1073 0.0732424
R576 VSS.n1072 VSS.n1074 2.21488
R577 VSS.n1077 VSS.n1076 0.0732424
R578 VSS.n1072 VSS.n1077 2.21488
R579 VSS.n1086 VSS.n1087 4.5005
R580 VSS.n1088 VSS.n1089 0.0732424
R581 VSS.n1089 VSS.n1087 2.21488
R582 VSS.n2243 VSS.n1087 2.21488
R583 VSS.n2242 VSS.n2243 4.57324
R584 VSS.n1092 VSS.n1093 4.5005
R585 VSS.n1095 VSS.n1094 0.0732424
R586 VSS.n1093 VSS.n1095 2.21488
R587 VSS.n1098 VSS.n1097 0.0732424
R588 VSS.n1093 VSS.n1098 2.21488
R589 VSS.n1107 VSS.n1108 4.5005
R590 VSS.n1110 VSS.n1109 0.0732424
R591 VSS.n1108 VSS.n1110 2.21488
R592 VSS.n1113 VSS.n1112 0.0732424
R593 VSS.n1108 VSS.n1113 2.21488
R594 VSS.n1122 VSS.n1123 4.5005
R595 VSS.n1125 VSS.n1124 0.0732424
R596 VSS.n1123 VSS.n1125 2.21488
R597 VSS.n1128 VSS.n1127 0.0732424
R598 VSS.n1123 VSS.n1128 2.21488
R599 VSS.n1137 VSS.n1138 4.5005
R600 VSS.n1139 VSS.n1140 0.0732424
R601 VSS.n1140 VSS.n1138 2.21488
R602 VSS.n2252 VSS.n1138 2.21488
R603 VSS.n2251 VSS.n2252 4.57324
R604 VSS.n1143 VSS.n1144 4.5005
R605 VSS.n1146 VSS.n1145 0.0732424
R606 VSS.n1144 VSS.n1146 2.21488
R607 VSS.n1149 VSS.n1148 0.0732424
R608 VSS.n1144 VSS.n1149 2.21488
R609 VSS.n1158 VSS.n1159 4.5005
R610 VSS.n1161 VSS.n1160 0.0732424
R611 VSS.n1159 VSS.n1161 2.21488
R612 VSS.n1164 VSS.n1163 0.0732424
R613 VSS.n1159 VSS.n1164 2.21488
R614 VSS.n1173 VSS.n1174 4.5005
R615 VSS.n1176 VSS.n1175 0.0732424
R616 VSS.n1174 VSS.n1176 2.21488
R617 VSS.n1179 VSS.n1178 0.0732424
R618 VSS.n1174 VSS.n1179 2.21488
R619 VSS.n1188 VSS.n1189 4.5005
R620 VSS.n1191 VSS.n1190 0.0732424
R621 VSS.n1189 VSS.n1191 2.21488
R622 VSS.n1194 VSS.n1193 0.0732424
R623 VSS.n1189 VSS.n1194 2.21488
R624 VSS.n1203 VSS.n1204 4.5005
R625 VSS.n1206 VSS.n1205 0.0732424
R626 VSS.n1204 VSS.n1206 2.21488
R627 VSS.n1209 VSS.n1208 0.0732424
R628 VSS.n1204 VSS.n1209 2.21488
R629 VSS.n1218 VSS.n1219 4.5005
R630 VSS.n1221 VSS.n1220 0.0732424
R631 VSS.n1219 VSS.n1221 2.21488
R632 VSS.n1224 VSS.n1223 0.0732424
R633 VSS.n1219 VSS.n1224 2.21488
R634 VSS.n1233 VSS.n1234 4.5005
R635 VSS.n1235 VSS.n1236 0.0732424
R636 VSS.n1236 VSS.n1234 2.21488
R637 VSS.n2261 VSS.n1234 2.21488
R638 VSS.n2260 VSS.n2261 4.57324
R639 VSS.n1239 VSS.n1240 4.5005
R640 VSS.n1242 VSS.n1241 0.0732424
R641 VSS.n1240 VSS.n1242 2.21488
R642 VSS.n1245 VSS.n1244 0.0732424
R643 VSS.n1240 VSS.n1245 2.21488
R644 VSS.n1254 VSS.n1255 4.5005
R645 VSS.n1257 VSS.n1256 0.0732424
R646 VSS.n1255 VSS.n1257 2.21488
R647 VSS.n1260 VSS.n1259 0.0732424
R648 VSS.n1255 VSS.n1260 2.21488
R649 VSS.n1269 VSS.n1270 4.5005
R650 VSS.n1272 VSS.n1271 0.0732424
R651 VSS.n1270 VSS.n1272 2.21488
R652 VSS.n1275 VSS.n1274 0.0732424
R653 VSS.n1270 VSS.n1275 2.21488
R654 VSS.n1284 VSS.n1285 4.5005
R655 VSS.n1286 VSS.n1287 0.0732424
R656 VSS.n1287 VSS.n1285 2.21488
R657 VSS.n2270 VSS.n1285 2.21488
R658 VSS.n2269 VSS.n2270 4.57324
R659 VSS.n1290 VSS.n1291 4.5005
R660 VSS.n1293 VSS.n1292 0.0732424
R661 VSS.n1291 VSS.n1293 2.21488
R662 VSS.n1296 VSS.n1295 0.0732424
R663 VSS.n1291 VSS.n1296 2.21488
R664 VSS.n1305 VSS.n1306 4.5005
R665 VSS.n1308 VSS.n1307 0.0732424
R666 VSS.n1306 VSS.n1308 2.21488
R667 VSS.n1311 VSS.n1310 0.0732424
R668 VSS.n1306 VSS.n1311 2.21488
R669 VSS.n1320 VSS.n1321 4.5005
R670 VSS.n1323 VSS.n1322 0.0732424
R671 VSS.n1321 VSS.n1323 2.21488
R672 VSS.n1326 VSS.n1325 0.0732424
R673 VSS.n1321 VSS.n1326 2.21488
R674 VSS.n1335 VSS.n1336 4.5005
R675 VSS.n1338 VSS.n1337 0.0732424
R676 VSS.n1336 VSS.n1338 2.21488
R677 VSS.n1341 VSS.n1340 0.0732424
R678 VSS.n1336 VSS.n1341 2.21488
R679 VSS.n1350 VSS.n1351 4.5005
R680 VSS.n1352 VSS.n1353 0.0732424
R681 VSS.n1353 VSS.n1351 2.21488
R682 VSS.n2279 VSS.n1351 2.21488
R683 VSS.n2278 VSS.n2279 4.57324
R684 VSS.n1356 VSS.n1357 4.5005
R685 VSS.n1359 VSS.n1358 0.0732424
R686 VSS.n1357 VSS.n1359 2.21488
R687 VSS.n1362 VSS.n1361 0.0732424
R688 VSS.n1357 VSS.n1362 2.21488
R689 VSS.n1371 VSS.n1372 4.5005
R690 VSS.n1374 VSS.n1373 0.0732424
R691 VSS.n1372 VSS.n1374 2.21488
R692 VSS.n1377 VSS.n1376 0.0732424
R693 VSS.n1372 VSS.n1377 2.21488
R694 VSS.n1386 VSS.n1387 4.5005
R695 VSS.n1389 VSS.n1388 0.0732424
R696 VSS.n1387 VSS.n1389 2.21488
R697 VSS.n1392 VSS.n1391 0.0732424
R698 VSS.n1387 VSS.n1392 2.21488
R699 VSS.n1401 VSS.n1402 4.5005
R700 VSS.n1403 VSS.n1404 0.0732424
R701 VSS.n1404 VSS.n1402 2.21488
R702 VSS.n2288 VSS.n1402 2.21488
R703 VSS.n2287 VSS.n2288 4.57324
R704 VSS.n1407 VSS.n1408 4.5005
R705 VSS.n1410 VSS.n1409 0.0732424
R706 VSS.n1408 VSS.n1410 2.21488
R707 VSS.n1413 VSS.n1412 0.0732424
R708 VSS.n1408 VSS.n1413 2.21488
R709 VSS.n1422 VSS.n1423 4.5005
R710 VSS.n1425 VSS.n1424 0.0732424
R711 VSS.n1423 VSS.n1425 2.21488
R712 VSS.n1428 VSS.n1427 0.0732424
R713 VSS.n1423 VSS.n1428 2.21488
R714 VSS.n1437 VSS.n1438 4.5005
R715 VSS.n1440 VSS.n1439 0.0732424
R716 VSS.n1438 VSS.n1440 2.21488
R717 VSS.n1443 VSS.n1442 0.0732424
R718 VSS.n1438 VSS.n1443 2.21488
R719 VSS.n1452 VSS.n1453 4.5005
R720 VSS.n1455 VSS.n1454 0.0732424
R721 VSS.n1453 VSS.n1455 2.21488
R722 VSS.n1458 VSS.n1457 0.0732424
R723 VSS.n1453 VSS.n1458 2.21488
R724 VSS.n1467 VSS.n1468 4.5005
R725 VSS.n1470 VSS.n1469 0.0732424
R726 VSS.n1468 VSS.n1470 2.21488
R727 VSS.n1473 VSS.n1472 0.0732424
R728 VSS.n1468 VSS.n1473 2.21488
R729 VSS.n1482 VSS.n1483 4.5005
R730 VSS.n1485 VSS.n1484 0.0732424
R731 VSS.n1483 VSS.n1485 2.21488
R732 VSS.n1488 VSS.n1487 0.0732424
R733 VSS.n1483 VSS.n1488 2.21488
R734 VSS.n1497 VSS.n1498 4.5005
R735 VSS.n1500 VSS.n1499 0.0732424
R736 VSS.n1498 VSS.n1500 2.21488
R737 VSS.n1498 VSS.n2297 2.21488
R738 VSS.n2297 VSS.n2296 4.57324
R739 VSS.n1503 VSS.n1504 4.5005
R740 VSS.n1506 VSS.n1505 0.0732424
R741 VSS.n1504 VSS.n1506 2.21488
R742 VSS.n1509 VSS.n1508 0.0732424
R743 VSS.n1504 VSS.n1509 2.21488
R744 VSS.n1518 VSS.n1519 4.5005
R745 VSS.n1521 VSS.n1520 0.0732424
R746 VSS.n1519 VSS.n1521 2.21488
R747 VSS.n1524 VSS.n1523 0.0732424
R748 VSS.n1519 VSS.n1524 2.21488
R749 VSS.n1533 VSS.n1534 4.5005
R750 VSS.n1536 VSS.n1535 0.0732424
R751 VSS.n1534 VSS.n1536 2.21488
R752 VSS.n1539 VSS.n1538 0.0732424
R753 VSS.n1534 VSS.n1539 2.21488
R754 VSS.n1548 VSS.n1549 4.5005
R755 VSS.n1551 VSS.n1550 0.0732424
R756 VSS.n1549 VSS.n1551 2.21488
R757 VSS.n1549 VSS.n2306 2.21488
R758 VSS.n2306 VSS.n2305 4.57324
R759 VSS.n1554 VSS.n1555 4.5005
R760 VSS.n1557 VSS.n1556 0.0732424
R761 VSS.n1555 VSS.n1557 2.21488
R762 VSS.n1560 VSS.n1559 0.0732424
R763 VSS.n1555 VSS.n1560 2.21488
R764 VSS.n1569 VSS.n1570 4.5005
R765 VSS.n1572 VSS.n1571 0.0732424
R766 VSS.n1570 VSS.n1572 2.21488
R767 VSS.n1575 VSS.n1574 0.0732424
R768 VSS.n1570 VSS.n1575 2.21488
R769 VSS.n1584 VSS.n1585 4.5005
R770 VSS.n1587 VSS.n1586 0.0732424
R771 VSS.n1585 VSS.n1587 2.21488
R772 VSS.n1590 VSS.n1589 0.0732424
R773 VSS.n1585 VSS.n1590 2.21488
R774 VSS.n1599 VSS.n1600 4.5005
R775 VSS.n1602 VSS.n1601 0.0732424
R776 VSS.n1600 VSS.n1602 2.21488
R777 VSS.n1605 VSS.n1604 0.0732424
R778 VSS.n1600 VSS.n1605 2.21488
R779 VSS.n1614 VSS.n1615 4.5005
R780 VSS.n1617 VSS.n1616 0.0732424
R781 VSS.n1615 VSS.n1617 2.21488
R782 VSS.n1615 VSS.n2315 2.21488
R783 VSS.n2315 VSS.n2314 4.57324
R784 VSS.n1620 VSS.n1621 4.5005
R785 VSS.n1623 VSS.n1622 0.0732424
R786 VSS.n1621 VSS.n1623 2.21488
R787 VSS.n1626 VSS.n1625 0.0732424
R788 VSS.n1621 VSS.n1626 2.21488
R789 VSS.n1635 VSS.n1636 4.5005
R790 VSS.n1638 VSS.n1637 0.0732424
R791 VSS.n1636 VSS.n1638 2.21488
R792 VSS.n1641 VSS.n1640 0.0732424
R793 VSS.n1636 VSS.n1641 2.21488
R794 VSS.n1650 VSS.n1651 4.5005
R795 VSS.n1653 VSS.n1652 0.0732424
R796 VSS.n1651 VSS.n1653 2.21488
R797 VSS.n1656 VSS.n1655 0.0732424
R798 VSS.n1651 VSS.n1656 2.21488
R799 VSS.n1665 VSS.n1666 4.5005
R800 VSS.n1668 VSS.n1667 0.0732424
R801 VSS.n1666 VSS.n1668 2.21488
R802 VSS.n1666 VSS.n2324 2.21488
R803 VSS.n2324 VSS.n2323 4.57324
R804 VSS.n1671 VSS.n1672 4.5005
R805 VSS.n1674 VSS.n1673 0.0732424
R806 VSS.n1672 VSS.n1674 2.21488
R807 VSS.n1677 VSS.n1676 0.0732424
R808 VSS.n1672 VSS.n1677 2.21488
R809 VSS.n1686 VSS.n1687 4.5005
R810 VSS.n1689 VSS.n1688 0.0732424
R811 VSS.n1687 VSS.n1689 2.21488
R812 VSS.n1692 VSS.n1691 0.0732424
R813 VSS.n1687 VSS.n1692 2.21488
R814 VSS.n1701 VSS.n1702 4.5005
R815 VSS.n1704 VSS.n1703 0.0732424
R816 VSS.n1702 VSS.n1704 2.21488
R817 VSS.n1707 VSS.n1706 0.0732424
R818 VSS.n1702 VSS.n1707 2.21488
R819 VSS.n1716 VSS.n1717 4.5005
R820 VSS.n1719 VSS.n1718 0.0732424
R821 VSS.n1717 VSS.n1719 2.21488
R822 VSS.n1722 VSS.n1721 0.0732424
R823 VSS.n1717 VSS.n1722 2.21488
R824 VSS.n1731 VSS.n1732 4.5005
R825 VSS.n1734 VSS.n1733 0.0732424
R826 VSS.n1732 VSS.n1734 2.21488
R827 VSS.n1737 VSS.n1736 0.0732424
R828 VSS.n1732 VSS.n1737 2.21488
R829 VSS.n1746 VSS.n1747 4.5005
R830 VSS.n1749 VSS.n1748 0.0732424
R831 VSS.n1747 VSS.n1749 2.21488
R832 VSS.n1752 VSS.n1751 0.0732424
R833 VSS.n1747 VSS.n1752 2.21488
R834 VSS.n1761 VSS.n1762 4.5005
R835 VSS.n1764 VSS.n1763 0.0732424
R836 VSS.n1762 VSS.n1764 2.21488
R837 VSS.n1762 VSS.n2333 2.21488
R838 VSS.n2333 VSS.n2332 4.57324
R839 VSS.n1767 VSS.n1768 4.5005
R840 VSS.n1770 VSS.n1769 0.0732424
R841 VSS.n1768 VSS.n1770 2.21488
R842 VSS.n1773 VSS.n1772 0.0732424
R843 VSS.n1768 VSS.n1773 2.21488
R844 VSS.n1782 VSS.n1783 4.5005
R845 VSS.n1785 VSS.n1784 0.0732424
R846 VSS.n1783 VSS.n1785 2.21488
R847 VSS.n1788 VSS.n1787 0.0732424
R848 VSS.n1783 VSS.n1788 2.21488
R849 VSS.n1797 VSS.n1798 4.5005
R850 VSS.n1800 VSS.n1799 0.0732424
R851 VSS.n1798 VSS.n1800 2.21488
R852 VSS.n1803 VSS.n1802 0.0732424
R853 VSS.n1798 VSS.n1803 2.21488
R854 VSS.n1812 VSS.n1813 4.5005
R855 VSS.n1815 VSS.n1814 0.0732424
R856 VSS.n1813 VSS.n1815 2.21488
R857 VSS.n1813 VSS.n2342 2.21488
R858 VSS.n2342 VSS.n2341 4.57324
R859 VSS.n1818 VSS.n1819 4.5005
R860 VSS.n1821 VSS.n1820 0.0732424
R861 VSS.n1819 VSS.n1821 2.21488
R862 VSS.n1824 VSS.n1823 0.0732424
R863 VSS.n1819 VSS.n1824 2.21488
R864 VSS.n1833 VSS.n1834 4.5005
R865 VSS.n1836 VSS.n1835 0.0732424
R866 VSS.n1834 VSS.n1836 2.21488
R867 VSS.n1839 VSS.n1838 0.0732424
R868 VSS.n1834 VSS.n1839 2.21488
R869 VSS.n1848 VSS.n1849 4.5005
R870 VSS.n1851 VSS.n1850 0.0732424
R871 VSS.n1849 VSS.n1851 2.21488
R872 VSS.n1854 VSS.n1853 0.0732424
R873 VSS.n1849 VSS.n1854 2.21488
R874 VSS.n1863 VSS.n1864 4.5005
R875 VSS.n1866 VSS.n1865 0.0732424
R876 VSS.n1864 VSS.n1866 2.21488
R877 VSS.n1869 VSS.n1868 0.0732424
R878 VSS.n1864 VSS.n1869 2.21488
R879 VSS.n1878 VSS.n1879 4.5005
R880 VSS.n1881 VSS.n1880 0.0732424
R881 VSS.n1879 VSS.n1881 2.21488
R882 VSS.n1879 VSS.n2351 2.21488
R883 VSS.n2351 VSS.n2350 4.57324
R884 VSS.n1884 VSS.n1885 4.5005
R885 VSS.n1887 VSS.n1886 0.0732424
R886 VSS.n1885 VSS.n1887 2.21488
R887 VSS.n1890 VSS.n1889 0.0732424
R888 VSS.n1885 VSS.n1890 2.21488
R889 VSS.n1899 VSS.n1900 4.5005
R890 VSS.n1902 VSS.n1901 0.0732424
R891 VSS.n1900 VSS.n1902 2.21488
R892 VSS.n1905 VSS.n1904 0.0732424
R893 VSS.n1900 VSS.n1905 2.21488
R894 VSS.n1914 VSS.n1915 4.5005
R895 VSS.n1917 VSS.n1916 0.0732424
R896 VSS.n1915 VSS.n1917 2.21488
R897 VSS.n1920 VSS.n1919 0.0732424
R898 VSS.n1915 VSS.n1920 2.21488
R899 VSS.n1929 VSS.n1930 4.5005
R900 VSS.n1932 VSS.n1931 0.0732424
R901 VSS.n1930 VSS.n1932 2.21488
R902 VSS.n1930 VSS.n2360 2.21488
R903 VSS.n2360 VSS.n2359 4.57324
R904 VSS.n1935 VSS.n1936 4.5005
R905 VSS.n1938 VSS.n1937 0.0732424
R906 VSS.n1936 VSS.n1938 2.21488
R907 VSS.n1941 VSS.n1940 0.0732424
R908 VSS.n1936 VSS.n1941 2.21488
R909 VSS.n1950 VSS.n1951 4.5005
R910 VSS.n1953 VSS.n1952 0.0732424
R911 VSS.n1951 VSS.n1953 2.21488
R912 VSS.n1956 VSS.n1955 0.0732424
R913 VSS.n1951 VSS.n1956 2.21488
R914 VSS.n1965 VSS.n1966 4.5005
R915 VSS.n1968 VSS.n1967 0.0732424
R916 VSS.n1966 VSS.n1968 2.21488
R917 VSS.n1971 VSS.n1970 0.0732424
R918 VSS.n1966 VSS.n1971 2.21488
R919 VSS.n1980 VSS.n1981 4.5005
R920 VSS.n1983 VSS.n1982 0.0732424
R921 VSS.n1981 VSS.n1983 2.21488
R922 VSS.n1986 VSS.n1985 0.0732424
R923 VSS.n1981 VSS.n1986 2.21488
R924 VSS.n1995 VSS.n1996 4.5005
R925 VSS.n1998 VSS.n1997 0.0732424
R926 VSS.n1996 VSS.n1998 2.21488
R927 VSS.n2001 VSS.n2000 0.0732424
R928 VSS.n1996 VSS.n2001 2.21488
R929 VSS.n2010 VSS.n2011 4.5005
R930 VSS.n2013 VSS.n2012 0.0732424
R931 VSS.n2011 VSS.n2013 2.21488
R932 VSS.n2016 VSS.n2015 0.0732424
R933 VSS.n2011 VSS.n2016 2.21488
R934 VSS.n2025 VSS.n2026 4.5005
R935 VSS.n2027 VSS.n2028 0.0732424
R936 VSS.n2028 VSS.n2026 2.21488
R937 VSS.n2369 VSS.n2026 2.21488
R938 VSS.n2368 VSS.n2369 4.57324
R939 VSS.n2031 VSS.n2032 4.5005
R940 VSS.n2034 VSS.n2033 0.0732424
R941 VSS.n2032 VSS.n2034 2.21488
R942 VSS.n2037 VSS.n2036 0.0732424
R943 VSS.n2032 VSS.n2037 2.21488
R944 VSS.n2046 VSS.n2047 4.5005
R945 VSS.n2049 VSS.n2048 0.0732424
R946 VSS.n2047 VSS.n2049 2.21488
R947 VSS.n2052 VSS.n2051 0.0732424
R948 VSS.n2047 VSS.n2052 2.21488
R949 VSS.n2061 VSS.n2062 4.5005
R950 VSS.n2064 VSS.n2063 0.0732424
R951 VSS.n2062 VSS.n2064 2.21488
R952 VSS.n2067 VSS.n2066 0.0732424
R953 VSS.n2062 VSS.n2067 2.21488
R954 VSS.n2076 VSS.n2077 4.5005
R955 VSS.n2078 VSS.n2079 0.0732424
R956 VSS.n2079 VSS.n2077 2.21488
R957 VSS.n2081 VSS.n2082 0.0732424
R958 VSS.n2082 VSS.n2077 2.21488
R959 VSS.n9895 VSS.n9896 4.5005
R960 VSS.n9898 VSS.n9897 0.0732424
R961 VSS.n9896 VSS.n9898 2.21488
R962 VSS.n9901 VSS.n9900 0.0732424
R963 VSS.n9896 VSS.n9901 2.21488
R964 VSS.n9910 VSS.n9911 4.5005
R965 VSS.n9913 VSS.n9912 0.0732424
R966 VSS.n9911 VSS.n9913 2.21488
R967 VSS.n9916 VSS.n9915 0.0732424
R968 VSS.n9911 VSS.n9916 2.21488
R969 VSS.n9896 VSS.n9911 0.0584021
R970 VSS.n2077 VSS.n9896 0.0596608
R971 VSS.n2077 VSS.n2062 0.0244161
R972 VSS.n2062 VSS.n2047 0.0585594
R973 VSS.n2047 VSS.n2032 0.0584021
R974 VSS.n2026 VSS.n2032 0.0596608
R975 VSS.n2026 VSS.n2011 0.0244161
R976 VSS.n2011 VSS.n1996 0.0585594
R977 VSS.n1996 VSS.n1981 0.0584021
R978 VSS.n1981 VSS 0.16272
R979 VSS VSS.n1966 0.143052
R980 VSS.n1951 VSS.n1966 0.0584021
R981 VSS.n1936 VSS.n1951 0.0584021
R982 VSS.n1930 VSS.n1936 0.0244161
R983 VSS.n1915 VSS.n1930 0.0598182
R984 VSS.n1900 VSS.n1915 0.0584021
R985 VSS.n1885 VSS.n1900 0.0584021
R986 VSS.n1879 VSS.n1885 0.0244161
R987 VSS.n1864 VSS.n1879 0.0598182
R988 VSS.n1849 VSS.n1864 0.0584021
R989 VSS.n1834 VSS.n1849 0.0231573
R990 VSS.n1819 VSS.n1834 0.0584021
R991 VSS.n1813 VSS.n1819 0.0596608
R992 VSS.n1798 VSS.n1813 0.0244161
R993 VSS.n1783 VSS.n1798 0.0585594
R994 VSS.n1768 VSS.n1783 0.0584021
R995 VSS.n1762 VSS.n1768 0.0596608
R996 VSS.n1747 VSS.n1762 0.0244161
R997 VSS.n1732 VSS.n1747 0.0585594
R998 VSS.n1717 VSS.n1732 0.0584021
R999 VSS VSS.n1717 0.16272
R1000 VSS VSS.n1702 0.143052
R1001 VSS.n1702 VSS.n1687 0.0584021
R1002 VSS.n1687 VSS.n1672 0.0584021
R1003 VSS.n1672 VSS.n1666 0.0244161
R1004 VSS.n1666 VSS.n1651 0.0598182
R1005 VSS.n1651 VSS.n1636 0.0584021
R1006 VSS.n1636 VSS.n1621 0.0584021
R1007 VSS.n1621 VSS.n1615 0.0244161
R1008 VSS.n1615 VSS.n1600 0.0598182
R1009 VSS.n1600 VSS.n1585 0.0584021
R1010 VSS.n1585 VSS.n1570 0.0231573
R1011 VSS.n1570 VSS.n1555 0.0584021
R1012 VSS.n1555 VSS.n1549 0.0596608
R1013 VSS.n1549 VSS.n1534 0.0244161
R1014 VSS.n1534 VSS.n1519 0.0585594
R1015 VSS.n1519 VSS.n1504 0.0584021
R1016 VSS.n1504 VSS.n1498 0.0596608
R1017 VSS.n1498 VSS.n1483 0.0244161
R1018 VSS.n1483 VSS.n1468 0.0585594
R1019 VSS.n1468 VSS.n1453 0.0584021
R1020 VSS.n1453 VSS 0.16272
R1021 VSS VSS.n1438 0.143052
R1022 VSS.n1423 VSS.n1438 0.0584021
R1023 VSS.n1408 VSS.n1423 0.0584021
R1024 VSS.n1402 VSS.n1408 0.0244161
R1025 VSS.n1402 VSS.n1387 0.0598182
R1026 VSS.n1387 VSS.n1372 0.0584021
R1027 VSS.n1357 VSS.n1372 0.0584021
R1028 VSS.n1351 VSS.n1357 0.0244161
R1029 VSS.n1351 VSS.n1336 0.0598182
R1030 VSS.n1336 VSS.n1321 0.0584021
R1031 VSS.n1321 VSS.n1306 0.0231573
R1032 VSS.n1291 VSS.n1306 0.0584021
R1033 VSS.n1285 VSS.n1291 0.0596608
R1034 VSS.n1285 VSS.n1270 0.0244161
R1035 VSS.n1270 VSS.n1255 0.0585594
R1036 VSS.n1255 VSS.n1240 0.0584021
R1037 VSS.n1234 VSS.n1240 0.0596608
R1038 VSS.n1234 VSS.n1219 0.0244161
R1039 VSS.n1219 VSS.n1204 0.0585594
R1040 VSS.n1204 VSS.n1189 0.0584021
R1041 VSS.n1189 VSS 0.16272
R1042 VSS VSS.n1174 0.143052
R1043 VSS.n1159 VSS.n1174 0.0584021
R1044 VSS.n1144 VSS.n1159 0.0584021
R1045 VSS.n1138 VSS.n1144 0.0244161
R1046 VSS.n1138 VSS.n1123 0.0598182
R1047 VSS.n1123 VSS.n1108 0.0584021
R1048 VSS.n1093 VSS.n1108 0.0584021
R1049 VSS.n1087 VSS.n1093 0.0244161
R1050 VSS.n1087 VSS.n1072 0.0598182
R1051 VSS.n1072 VSS.n1057 0.0584021
R1052 VSS.n1057 VSS.n1042 0.0231573
R1053 VSS.n1027 VSS.n1042 0.0584021
R1054 VSS.n1021 VSS.n1027 0.0596608
R1055 VSS.n1021 VSS.n1006 0.0244161
R1056 VSS.n1006 VSS.n991 0.0585594
R1057 VSS.n991 VSS.n976 0.0584021
R1058 VSS.n970 VSS.n976 0.0596608
R1059 VSS.n970 VSS.n955 0.0244161
R1060 VSS.n955 VSS.n940 0.0585594
R1061 VSS.n940 VSS.n925 0.0584021
R1062 VSS.n925 VSS 0.16272
R1063 VSS VSS.n910 0.143052
R1064 VSS.n895 VSS.n910 0.0584021
R1065 VSS.n880 VSS.n895 0.0584021
R1066 VSS.n874 VSS.n880 0.0244161
R1067 VSS.n874 VSS.n859 0.0598182
R1068 VSS.n859 VSS.n844 0.0584021
R1069 VSS.n829 VSS.n844 0.0584021
R1070 VSS.n823 VSS.n829 0.0244161
R1071 VSS.n823 VSS.n808 0.0598182
R1072 VSS.n808 VSS.n793 0.0584021
R1073 VSS.n793 VSS.n778 0.0231573
R1074 VSS.n763 VSS.n778 0.0584021
R1075 VSS.n757 VSS.n763 0.0596608
R1076 VSS.n757 VSS.n742 0.0244161
R1077 VSS.n742 VSS.n727 0.0585594
R1078 VSS.n727 VSS.n712 0.0584021
R1079 VSS.n706 VSS.n712 0.0596608
R1080 VSS.n706 VSS.n691 0.0244161
R1081 VSS.n691 VSS.n676 0.0585594
R1082 VSS.n676 VSS.n661 0.0584021
R1083 VSS.n661 VSS 0.16272
R1084 VSS VSS.n646 0.143052
R1085 VSS.n631 VSS.n646 0.0584021
R1086 VSS.n616 VSS.n631 0.0584021
R1087 VSS.n610 VSS.n616 0.0244161
R1088 VSS.n610 VSS.n595 0.0598182
R1089 VSS.n595 VSS.n580 0.0584021
R1090 VSS.n565 VSS.n580 0.0584021
R1091 VSS.n559 VSS.n565 0.0244161
R1092 VSS.n559 VSS.n544 0.0598182
R1093 VSS.n544 VSS.n529 0.0584021
R1094 VSS.n529 VSS.n514 0.0231573
R1095 VSS.n499 VSS.n514 0.0584021
R1096 VSS.n493 VSS.n499 0.0596608
R1097 VSS.n493 VSS.n478 0.0244161
R1098 VSS.n478 VSS.n463 0.0585594
R1099 VSS.n463 VSS.n448 0.0584021
R1100 VSS.n442 VSS.n448 0.0596608
R1101 VSS.n442 VSS.n427 0.0244161
R1102 VSS.n427 VSS.n412 0.0585594
R1103 VSS.n412 VSS.n397 0.0584021
R1104 VSS.n397 VSS 0.16272
R1105 VSS VSS.n382 0.143052
R1106 VSS.n367 VSS.n382 0.0584021
R1107 VSS.n352 VSS.n367 0.0584021
R1108 VSS.n346 VSS.n352 0.0244161
R1109 VSS.n346 VSS.n331 0.0598182
R1110 VSS.n331 VSS.n316 0.0584021
R1111 VSS.n301 VSS.n316 0.0584021
R1112 VSS.n295 VSS.n301 0.0244161
R1113 VSS.n295 VSS.n280 0.0598182
R1114 VSS.n280 VSS.n265 0.0584021
R1115 VSS.n265 VSS.n250 0.0231573
R1116 VSS.n235 VSS.n250 0.0584021
R1117 VSS.n229 VSS.n235 0.0596608
R1118 VSS.n229 VSS.n214 0.0244161
R1119 VSS.n214 VSS.n199 0.0585594
R1120 VSS.n199 VSS.n184 0.0584021
R1121 VSS.n178 VSS.n184 0.0596608
R1122 VSS.n178 VSS.n163 0.0244161
R1123 VSS.n163 VSS.n148 0.0585594
R1124 VSS.n148 VSS.n133 0.0584021
R1125 VSS.n133 VSS 0.16272
R1126 VSS VSS.n118 0.143052
R1127 VSS.n103 VSS.n118 0.0584021
R1128 VSS.n88 VSS.n103 0.0584021
R1129 VSS.n82 VSS.n88 0.0244161
R1130 VSS.n82 VSS.n67 0.0598182
R1131 VSS.n67 VSS.n52 0.0584021
R1132 VSS.n37 VSS.n52 0.0584021
R1133 VSS.n31 VSS.n37 0.0244161
R1134 VSS.n31 VSS.n16 0.0598182
R1135 VSS.n16 VSS.n1 0.0584021
R1136 VSS.n9912 VSS.n9917 4.5005
R1137 VSS.n9914 VSS.n9918 4.5005
R1138 VSS.n9915 VSS.n9919 4.5005
R1139 VSS.n9916 VSS.n9920 4.57324
R1140 VSS.n9912 VSS.n9910 0.147342
R1141 VSS.n9913 VSS.n9914 0.0732424
R1142 VSS.n9914 VSS.n9915 0.147342
R1143 VSS.n9917 VSS.n9921 0.0721009
R1144 VSS.n9922 VSS.n9918 4.5005
R1145 VSS.n9923 VSS.n9919 4.5005
R1146 VSS.n9924 VSS.n9920 4.5005
R1147 VSS.n9910 VSS.n9921 4.57442
R1148 VSS.n9917 VSS.n9918 0.147342
R1149 VSS.n9918 VSS.n9919 0.147342
R1150 VSS.n9919 VSS.n9920 0.147342
R1151 VSS.n9921 VSS.n9922 2.39784
R1152 VSS.n9922 VSS.n9923 0.147342
R1153 VSS.n9923 VSS.n9924 0.147342
R1154 VSS.n9924 VSS.t221 3.13212
R1155 VSS.n9897 VSS.n9902 4.5005
R1156 VSS.n9899 VSS.n9903 4.5005
R1157 VSS.n9900 VSS.n9904 4.5005
R1158 VSS.n9901 VSS.n9905 4.57324
R1159 VSS.n9897 VSS.n9895 0.147342
R1160 VSS.n9898 VSS.n9899 0.0732424
R1161 VSS.n9899 VSS.n9900 0.147342
R1162 VSS.n9902 VSS.n9906 0.0721009
R1163 VSS.n9907 VSS.n9903 4.5005
R1164 VSS.n9908 VSS.n9904 4.5005
R1165 VSS.n9909 VSS.n9905 4.5005
R1166 VSS.n9895 VSS.n9906 4.57442
R1167 VSS.n9902 VSS.n9903 0.147342
R1168 VSS.n9903 VSS.n9904 0.147342
R1169 VSS.n9904 VSS.n9905 0.147342
R1170 VSS.n9906 VSS.n9907 2.39784
R1171 VSS.n9907 VSS.n9908 0.147342
R1172 VSS.n9908 VSS.n9909 0.147342
R1173 VSS.n9909 VSS.t292 3.13212
R1174 VSS.n2083 VSS.n2078 4.5005
R1175 VSS.n2084 VSS.n2080 4.5005
R1176 VSS.n2085 VSS.n2081 4.5005
R1177 VSS.n2086 VSS.n2082 4.57324
R1178 VSS.n2076 VSS.n2078 0.147342
R1179 VSS.n2079 VSS.n2080 0.0732424
R1180 VSS.n2080 VSS.n2081 0.147342
R1181 VSS.n2087 VSS.n2083 0.0722544
R1182 VSS.n2088 VSS.n2084 4.5005
R1183 VSS.n2089 VSS.n2085 4.5005
R1184 VSS.n9894 VSS.n2086 4.5005
R1185 VSS.n2087 VSS.n2076 4.57426
R1186 VSS.n2083 VSS.n2084 0.147342
R1187 VSS.n2084 VSS.n2085 0.147342
R1188 VSS.n2085 VSS.n2086 0.147342
R1189 VSS.n2088 VSS.n2087 2.37296
R1190 VSS.n2089 VSS.n2088 0.127318
R1191 VSS.n9894 VSS.n2089 0.127318
R1192 VSS.t20 VSS.n9894 2.73618
R1193 VSS.n2108 VSS.t31 0.154858
R1194 VSS.t31 VSS 8.59308
R1195 VSS VSS.t5 180.238
R1196 VSS.t0 VSS.t5 333.928
R1197 VSS.t41 VSS.t0 333.928
R1198 VSS.t20 VSS.t41 333.928
R1199 VSS.n2108 VSS.n9893 5.32359
R1200 VSS.n9570 VSS.n9665 13.5005
R1201 VSS.n9571 VSS.n9666 13.5005
R1202 VSS.n9572 VSS.n9667 13.5005
R1203 VSS.n9573 VSS.n9668 13.5005
R1204 VSS.n9574 VSS.n9669 13.5005
R1205 VSS.n9575 VSS.n9670 13.5005
R1206 VSS.n9576 VSS.n9671 13.5005
R1207 VSS.n9577 VSS.n9672 13.5005
R1208 VSS.n9578 VSS.n9673 13.5005
R1209 VSS.n9579 VSS.n9674 13.5005
R1210 VSS.n9580 VSS.n9675 13.5005
R1211 VSS.n9581 VSS.n9676 13.5005
R1212 VSS.n9582 VSS.n9677 13.5005
R1213 VSS.n9583 VSS.n9678 13.5005
R1214 VSS.n9584 VSS.n9679 13.5005
R1215 VSS.n9585 VSS.n9680 13.5005
R1216 VSS.n9586 VSS.n9681 13.5005
R1217 VSS.n9587 VSS.n9682 13.5005
R1218 VSS.n9588 VSS.n9683 13.5005
R1219 VSS.n9589 VSS.n9684 13.5005
R1220 VSS.n9590 VSS.n9685 13.5005
R1221 VSS.n9591 VSS.n9686 13.5005
R1222 VSS.n9592 VSS.n9687 13.5005
R1223 VSS.n9593 VSS.n9688 13.5005
R1224 VSS.n9594 VSS.n9689 13.5005
R1225 VSS.n9595 VSS.n9690 13.5005
R1226 VSS.n9596 VSS.n9691 13.5005
R1227 VSS.n9597 VSS.n9692 13.5005
R1228 VSS.n9598 VSS.n9693 13.5005
R1229 VSS.n9599 VSS.n9694 13.5005
R1230 VSS.n9600 VSS.n9695 13.5005
R1231 VSS.n9601 VSS.n9696 13.5005
R1232 VSS.n9602 VSS.n9697 13.5005
R1233 VSS.n9603 VSS.n9698 13.5005
R1234 VSS.n9604 VSS.n9699 13.5005
R1235 VSS.n9605 VSS.n9700 13.5005
R1236 VSS.n9606 VSS.n9701 13.5005
R1237 VSS.n9607 VSS.n9702 13.5005
R1238 VSS.n9608 VSS.n9703 13.5005
R1239 VSS.n9609 VSS.n9704 13.5005
R1240 VSS.n9610 VSS.n9705 13.5005
R1241 VSS.n9611 VSS.n9706 13.5005
R1242 VSS.n9612 VSS.n9707 13.5005
R1243 VSS.n9613 VSS.n9708 13.5005
R1244 VSS.n9614 VSS.n9709 13.5005
R1245 VSS.n9615 VSS.n9710 13.5005
R1246 VSS.n9616 VSS.n9711 13.5005
R1247 VSS.n9617 VSS.n9712 13.5005
R1248 VSS.n9618 VSS.n9713 13.5005
R1249 VSS.n9619 VSS.n9714 13.5005
R1250 VSS.n9620 VSS.n9715 13.5005
R1251 VSS.n9621 VSS.n9716 13.5005
R1252 VSS.n9622 VSS.n9717 13.5005
R1253 VSS.n9623 VSS.n9718 13.5005
R1254 VSS.n9624 VSS.n9719 13.5005
R1255 VSS.n9625 VSS.n9720 13.5005
R1256 VSS.n9626 VSS.n9721 13.5005
R1257 VSS.n9627 VSS.n9722 13.5005
R1258 VSS.n9628 VSS.n9723 13.5005
R1259 VSS.n9629 VSS.n9724 13.5005
R1260 VSS.n9630 VSS.n9725 13.5005
R1261 VSS.n9631 VSS.n9726 13.5005
R1262 VSS.n9632 VSS.n9727 13.5005
R1263 VSS.n9633 VSS.n9728 13.5005
R1264 VSS.n9634 VSS.n9729 13.5005
R1265 VSS.n9635 VSS.n9730 13.5005
R1266 VSS.n9636 VSS.n9731 13.5005
R1267 VSS.n9637 VSS.n9732 13.5005
R1268 VSS.n9638 VSS.n9733 13.5005
R1269 VSS.n9639 VSS.n9734 13.5005
R1270 VSS.n9640 VSS.n9735 13.5005
R1271 VSS.n9641 VSS.n9736 13.5005
R1272 VSS.n9642 VSS.n9737 13.5005
R1273 VSS.n9643 VSS.n9738 13.5005
R1274 VSS.n9644 VSS.n9739 13.5005
R1275 VSS.n9645 VSS.n9740 13.5005
R1276 VSS.n9646 VSS.n9741 13.5005
R1277 VSS.n9647 VSS.n9742 13.5005
R1278 VSS.n9648 VSS.n9743 13.5005
R1279 VSS.n9649 VSS.n9744 13.5005
R1280 VSS.n9650 VSS.n9745 13.5005
R1281 VSS.n9651 VSS.n9746 13.5005
R1282 VSS.n9652 VSS.n9747 13.5005
R1283 VSS.n9653 VSS.n9748 13.5005
R1284 VSS.n9654 VSS.n9749 13.5005
R1285 VSS.n9655 VSS.n9750 13.5005
R1286 VSS.n9656 VSS.n9751 13.5005
R1287 VSS.n9657 VSS.n9752 13.5005
R1288 VSS.n9658 VSS.n9753 13.5005
R1289 VSS.n9659 VSS.n9754 13.5005
R1290 VSS.n9660 VSS.n9755 13.5005
R1291 VSS.n9661 VSS.n9756 13.5005
R1292 VSS.n9662 VSS.n9757 13.5005
R1293 VSS.n9663 VSS.n9758 13.5005
R1294 VSS.n9665 VSS.n9893 13.7848
R1295 VSS.n9893 VSS.n9759 0.1415
R1296 VSS.n9759 VSS.n9570 0.29525
R1297 VSS.n9570 VSS.n9760 0.04175
R1298 VSS.n9760 VSS.n9761 0.3365
R1299 VSS.n9761 VSS.n9571 0.07325
R1300 VSS.n9571 VSS.n9762 0.29375
R1301 VSS.n9762 VSS.n9572 0.15725
R1302 VSS.n9572 VSS.n9763 0.01175
R1303 VSS.n9763 VSS.n9764 0.3665
R1304 VSS.n9764 VSS.n9573 0.07325
R1305 VSS.n9573 VSS.n9765 0.26375
R1306 VSS.n9765 VSS.n9574 0.18725
R1307 VSS.n9574 VSS.n9766 0.14975
R1308 VSS.n9766 VSS.n9575 0.75125
R1309 VSS.n9575 VSS.n9767 0.19775
R1310 VSS.n9767 VSS.n9576 0.25325
R1311 VSS.n9576 VSS.n9768 0.11375
R1312 VSS.n9768 VSS.n9769 0.1385
R1313 VSS.n9769 VSS.n9577 0.19925
R1314 VSS.n9577 VSS.n9770 0.13775
R1315 VSS.n9770 VSS.n9578 0.31325
R1316 VSS.n9578 VSS.n9771 0.02375
R1317 VSS.n9771 VSS.n9772 0.3365
R1318 VSS.n9772 VSS.n9579 0.09125
R1319 VSS.n9579 VSS.n9773 0.24575
R1320 VSS.n9773 VSS.n9580 0.20525
R1321 VSS.n9580 VSS.n9774 0.13175
R1322 VSS.n9774 VSS.n9581 0.377
R1323 VSS.n9581 VSS.n9775 0.01475
R1324 VSS.n9775 VSS.n9776 0.1415
R1325 VSS.n9776 VSS.n9582 0.29525
R1326 VSS.n9582 VSS.n9777 0.04175
R1327 VSS.n9777 VSS.n9778 0.3365
R1328 VSS.n9778 VSS.n9583 0.07325
R1329 VSS.n9583 VSS.n9779 0.29375
R1330 VSS.n9779 VSS.n9584 0.15725
R1331 VSS.n9584 VSS.n9780 0.01175
R1332 VSS.n9780 VSS.n9781 0.3665
R1333 VSS.n9781 VSS.n9585 0.07325
R1334 VSS.n9585 VSS.n9782 0.26375
R1335 VSS.n9782 VSS.n9586 0.18725
R1336 VSS.n9586 VSS.n9783 0.14975
R1337 VSS.n9783 VSS.n9587 0.75125
R1338 VSS.n9587 VSS.n9784 0.19775
R1339 VSS.n9784 VSS.n9588 0.25325
R1340 VSS.n9588 VSS.n9785 0.11375
R1341 VSS.n9785 VSS.n9786 0.1385
R1342 VSS.n9786 VSS.n9589 0.19925
R1343 VSS.n9589 VSS.n9787 0.13775
R1344 VSS.n9787 VSS.n9590 0.31325
R1345 VSS.n9590 VSS.n9788 0.02375
R1346 VSS.n9788 VSS.n9789 0.3365
R1347 VSS.n9789 VSS.n9591 0.09125
R1348 VSS.n9591 VSS.n9790 0.24575
R1349 VSS.n9790 VSS.n9592 0.20525
R1350 VSS.n9592 VSS.n9791 0.13175
R1351 VSS.n9791 VSS.n9593 0.377
R1352 VSS.n9593 VSS.n9792 0.01475
R1353 VSS.n9792 VSS.n9793 0.1415
R1354 VSS.n9793 VSS.n9594 0.29525
R1355 VSS.n9594 VSS.n9794 0.04175
R1356 VSS.n9794 VSS.n9795 0.3365
R1357 VSS.n9795 VSS.n9595 0.07325
R1358 VSS.n9595 VSS.n9796 0.29375
R1359 VSS.n9796 VSS.n9596 0.15725
R1360 VSS.n9596 VSS.n9797 0.01175
R1361 VSS.n9797 VSS.n9798 0.3665
R1362 VSS.n9798 VSS.n9597 0.07325
R1363 VSS.n9597 VSS.n9799 0.26375
R1364 VSS.n9799 VSS.n9598 0.18725
R1365 VSS.n9598 VSS.n9800 0.14975
R1366 VSS.n9800 VSS.n9599 0.75125
R1367 VSS.n9599 VSS.n9801 0.19775
R1368 VSS.n9801 VSS.n9600 0.25325
R1369 VSS.n9600 VSS.n9802 0.11375
R1370 VSS.n9802 VSS.n9803 0.1385
R1371 VSS.n9803 VSS.n9601 0.19925
R1372 VSS.n9601 VSS.n9804 0.13775
R1373 VSS.n9804 VSS.n9602 0.31325
R1374 VSS.n9602 VSS.n9805 0.02375
R1375 VSS.n9805 VSS.n9806 0.3365
R1376 VSS.n9806 VSS.n9603 0.09125
R1377 VSS.n9603 VSS.n9807 0.24575
R1378 VSS.n9807 VSS.n9604 0.20525
R1379 VSS.n9604 VSS.n9808 0.13175
R1380 VSS.n9808 VSS.n9605 0.377
R1381 VSS.n9605 VSS.n9809 0.01475
R1382 VSS.n9809 VSS.n9810 0.1415
R1383 VSS.n9810 VSS.n9606 0.29525
R1384 VSS.n9606 VSS.n9811 0.04175
R1385 VSS.n9811 VSS.n9812 0.3365
R1386 VSS.n9812 VSS.n9607 0.07325
R1387 VSS.n9607 VSS.n9813 0.29375
R1388 VSS.n9813 VSS.n9608 0.15725
R1389 VSS.n9608 VSS.n9814 0.01175
R1390 VSS.n9814 VSS.n9815 0.3665
R1391 VSS.n9815 VSS.n9609 0.07325
R1392 VSS.n9609 VSS.n9816 0.26375
R1393 VSS.n9816 VSS.n9610 0.18725
R1394 VSS.n9610 VSS.n9817 0.14975
R1395 VSS.n9817 VSS.n9611 0.75125
R1396 VSS.n9611 VSS.n9818 0.19775
R1397 VSS.n9818 VSS.n9612 0.25325
R1398 VSS.n9612 VSS.n9819 0.11375
R1399 VSS.n9819 VSS.n9820 0.1385
R1400 VSS.n9820 VSS.n9613 0.19925
R1401 VSS.n9613 VSS.n9821 0.13775
R1402 VSS.n9821 VSS.n9614 0.31325
R1403 VSS.n9614 VSS.n9822 0.02375
R1404 VSS.n9822 VSS.n9823 0.3365
R1405 VSS.n9823 VSS.n9615 0.09125
R1406 VSS.n9615 VSS.n9824 0.24575
R1407 VSS.n9824 VSS.n9616 0.20525
R1408 VSS.n9616 VSS.n9825 0.13175
R1409 VSS.n9825 VSS.n9617 0.377
R1410 VSS.n9617 VSS.n9826 0.01475
R1411 VSS.n9826 VSS.n9827 0.1415
R1412 VSS.n9827 VSS.n9618 0.29525
R1413 VSS.n9618 VSS.n9828 0.04175
R1414 VSS.n9828 VSS.n9829 0.3365
R1415 VSS.n9829 VSS.n9619 0.07325
R1416 VSS.n9619 VSS.n9830 0.29375
R1417 VSS.n9830 VSS.n9620 0.15725
R1418 VSS.n9620 VSS.n9831 0.01175
R1419 VSS.n9831 VSS.n9832 0.3665
R1420 VSS.n9832 VSS.n9621 0.07325
R1421 VSS.n9621 VSS.n9833 0.26375
R1422 VSS.n9833 VSS.n9622 0.18725
R1423 VSS.n9622 VSS.n9834 0.14975
R1424 VSS.n9834 VSS.n9623 0.75125
R1425 VSS.n9623 VSS.n9835 0.19775
R1426 VSS.n9835 VSS.n9624 0.25325
R1427 VSS.n9624 VSS.n9836 0.11375
R1428 VSS.n9836 VSS.n9837 0.1385
R1429 VSS.n9837 VSS.n9625 0.19925
R1430 VSS.n9625 VSS.n9838 0.13775
R1431 VSS.n9838 VSS.n9626 0.31325
R1432 VSS.n9626 VSS.n9839 0.02375
R1433 VSS.n9839 VSS.n9840 0.3365
R1434 VSS.n9840 VSS.n9627 0.09125
R1435 VSS.n9627 VSS.n9841 0.24575
R1436 VSS.n9841 VSS.n9628 0.20525
R1437 VSS.n9628 VSS.n9842 0.13175
R1438 VSS.n9842 VSS.n9629 0.377
R1439 VSS.n9629 VSS.n9843 0.01475
R1440 VSS.n9843 VSS.n9844 0.1415
R1441 VSS.n9844 VSS.n9630 0.29525
R1442 VSS.n9630 VSS.n9845 0.04175
R1443 VSS.n9845 VSS.n9846 0.3365
R1444 VSS.n9846 VSS.n9631 0.07325
R1445 VSS.n9631 VSS.n9847 0.29375
R1446 VSS.n9847 VSS.n9632 0.15725
R1447 VSS.n9632 VSS.n9848 0.01175
R1448 VSS.n9848 VSS.n9849 0.3665
R1449 VSS.n9849 VSS.n9633 0.07325
R1450 VSS.n9633 VSS.n9850 0.26375
R1451 VSS.n9850 VSS.n9634 0.18725
R1452 VSS.n9634 VSS.n9851 0.14975
R1453 VSS.n9851 VSS.n9635 0.75125
R1454 VSS.n9635 VSS.n9852 0.19775
R1455 VSS.n9852 VSS.n9636 0.25325
R1456 VSS.n9636 VSS.n9853 0.11375
R1457 VSS.n9853 VSS.n9854 0.1385
R1458 VSS.n9854 VSS.n9637 0.19925
R1459 VSS.n9637 VSS.n9855 0.13775
R1460 VSS.n9855 VSS.n9638 0.31325
R1461 VSS.n9638 VSS.n9856 0.02375
R1462 VSS.n9856 VSS.n9857 0.3365
R1463 VSS.n9857 VSS.n9639 0.09125
R1464 VSS.n9639 VSS.n9858 0.24575
R1465 VSS.n9858 VSS.n9640 0.20525
R1466 VSS.n9640 VSS.n9859 0.13175
R1467 VSS.n9859 VSS.n9641 0.377
R1468 VSS.n9641 VSS.n9860 0.01475
R1469 VSS.n9860 VSS.n9861 0.1415
R1470 VSS.n9861 VSS.n9642 0.29525
R1471 VSS.n9642 VSS.n9862 0.04175
R1472 VSS.n9862 VSS.n9863 0.3365
R1473 VSS.n9863 VSS.n9643 0.07325
R1474 VSS.n9643 VSS.n9864 0.29375
R1475 VSS.n9864 VSS.n9644 0.15725
R1476 VSS.n9644 VSS.n9865 0.01175
R1477 VSS.n9865 VSS.n9866 0.3665
R1478 VSS.n9866 VSS.n9645 0.07325
R1479 VSS.n9645 VSS.n9867 0.26375
R1480 VSS.n9867 VSS.n9646 0.18725
R1481 VSS.n9646 VSS.n9868 0.14975
R1482 VSS.n9868 VSS.n9647 0.75125
R1483 VSS.n9647 VSS.n9869 0.19775
R1484 VSS.n9869 VSS.n9648 0.25325
R1485 VSS.n9648 VSS.n9870 0.11375
R1486 VSS.n9870 VSS.n9871 0.1385
R1487 VSS.n9871 VSS.n9649 0.19925
R1488 VSS.n9649 VSS.n9872 0.13775
R1489 VSS.n9872 VSS.n9650 0.31325
R1490 VSS.n9650 VSS.n9873 0.02375
R1491 VSS.n9873 VSS.n9874 0.3365
R1492 VSS.n9874 VSS.n9651 0.09125
R1493 VSS.n9651 VSS.n9875 0.24575
R1494 VSS.n9875 VSS.n9652 0.20525
R1495 VSS.n9652 VSS.n9876 0.13175
R1496 VSS.n9876 VSS.n9653 0.377
R1497 VSS.n9653 VSS.n9877 0.01475
R1498 VSS.n9877 VSS.n9878 0.1415
R1499 VSS.n9878 VSS.n9654 0.29525
R1500 VSS.n9654 VSS.n9879 0.04175
R1501 VSS.n9879 VSS.n9880 0.3365
R1502 VSS.n9880 VSS.n9655 0.07325
R1503 VSS.n9655 VSS.n9881 0.29375
R1504 VSS.n9881 VSS.n9656 0.15725
R1505 VSS.n9656 VSS.n9882 0.01175
R1506 VSS.n9882 VSS.n9883 0.3665
R1507 VSS.n9883 VSS.n9657 0.07325
R1508 VSS.n9657 VSS.n9884 0.26375
R1509 VSS.n9884 VSS.n9658 0.18725
R1510 VSS.n9658 VSS.n9885 0.14975
R1511 VSS.n9885 VSS.n9659 0.75125
R1512 VSS.n9659 VSS.n9886 0.19775
R1513 VSS.n9886 VSS.n9660 0.25325
R1514 VSS.n9660 VSS.n9887 0.11375
R1515 VSS.n9887 VSS.n9888 0.1385
R1516 VSS.n9888 VSS.n9661 0.19925
R1517 VSS.n9661 VSS.n9889 0.13775
R1518 VSS.n9889 VSS.n9662 0.31325
R1519 VSS.n9662 VSS.n9890 0.02375
R1520 VSS.n9890 VSS.n9891 0.3365
R1521 VSS.n9891 VSS.n9663 0.09125
R1522 VSS.n9663 VSS.n9892 0.24575
R1523 VSS.n9892 VSS.n9664 0.20525
R1524 VSS.n9664 VSS.t332 8.64257
R1525 VSS.n9892 VSS.t416 8.51132
R1526 VSS.n9891 VSS.t204 8.51132
R1527 VSS.n9890 VSS.t318 8.51132
R1528 VSS.n9889 VSS.t161 8.51132
R1529 VSS.n9888 VSS.t159 8.51132
R1530 VSS.n2108 VSS.n9887 5.32359
R1531 VSS.n9886 VSS.t428 8.51132
R1532 VSS.t329 VSS.n9885 8.51132
R1533 VSS.t334 VSS.n9884 8.51132
R1534 VSS.t516 VSS.n9883 8.51132
R1535 VSS.n2108 VSS.n9882 5.32359
R1536 VSS.n2108 VSS.n9881 5.32359
R1537 VSS.n9880 VSS.t570 8.51132
R1538 VSS.n9879 VSS.t506 8.51132
R1539 VSS.n9878 VSS.t510 8.51132
R1540 VSS.n2108 VSS.n9877 5.32359
R1541 VSS.n9876 VSS.t224 8.51132
R1542 VSS.n9875 VSS.t399 8.51132
R1543 VSS.n9874 VSS.t551 8.51132
R1544 VSS.n9873 VSS.t438 8.51132
R1545 VSS.n9872 VSS.t493 8.51132
R1546 VSS.n9871 VSS.t228 8.51132
R1547 VSS.n2108 VSS.n9870 5.32359
R1548 VSS.n9869 VSS.t418 8.51132
R1549 VSS.t301 VSS.n9868 8.51132
R1550 VSS.t571 VSS.n9867 8.51132
R1551 VSS.t569 VSS.n9866 8.51132
R1552 VSS.n2108 VSS.n9865 5.32359
R1553 VSS.n2108 VSS.n9864 5.32359
R1554 VSS.n9863 VSS.t182 8.51132
R1555 VSS.n9862 VSS.t568 8.51132
R1556 VSS.n9861 VSS.t528 8.51132
R1557 VSS.n2108 VSS.n9860 5.32359
R1558 VSS.n9859 VSS.t401 8.51132
R1559 VSS.n9858 VSS.t598 8.51132
R1560 VSS.n9857 VSS.t514 8.51132
R1561 VSS.n9856 VSS.t57 8.51132
R1562 VSS.n9855 VSS.t360 8.51132
R1563 VSS.n9854 VSS.t299 8.51132
R1564 VSS.n2108 VSS.n9853 5.32359
R1565 VSS.n9852 VSS.t566 8.51132
R1566 VSS.t239 VSS.n9851 8.51132
R1567 VSS.t406 VSS.n9850 8.51132
R1568 VSS.t405 VSS.n9849 8.51132
R1569 VSS.n2108 VSS.n9848 5.32359
R1570 VSS.n2108 VSS.n9847 5.32359
R1571 VSS.n9846 VSS.t464 8.51132
R1572 VSS.n9845 VSS.t463 8.51132
R1573 VSS.n9844 VSS.t417 8.51132
R1574 VSS.n2108 VSS.n9843 5.32359
R1575 VSS.n9842 VSS.t413 8.51132
R1576 VSS.n9841 VSS.t494 8.51132
R1577 VSS.n9840 VSS.t546 8.51132
R1578 VSS.n9839 VSS.t124 8.51132
R1579 VSS.n9838 VSS.t40 8.51132
R1580 VSS.n9837 VSS.t400 8.51132
R1581 VSS.n2108 VSS.n9836 5.32359
R1582 VSS.n9835 VSS.t523 8.51132
R1583 VSS.t458 VSS.n9834 8.51132
R1584 VSS.t241 VSS.n9833 8.51132
R1585 VSS.t240 VSS.n9832 8.51132
R1586 VSS.n2108 VSS.n9831 5.32359
R1587 VSS.n2108 VSS.n9830 5.32359
R1588 VSS.n9829 VSS.t513 8.51132
R1589 VSS.n9828 VSS.t524 8.51132
R1590 VSS.n9827 VSS.t539 8.51132
R1591 VSS.n2108 VSS.n9826 5.32359
R1592 VSS.n9825 VSS.t32 8.51132
R1593 VSS.n9824 VSS.t143 8.51132
R1594 VSS.n9823 VSS.t203 8.51132
R1595 VSS.n9822 VSS.t565 8.51132
R1596 VSS.n9821 VSS.t312 8.51132
R1597 VSS.n9820 VSS.t431 8.51132
R1598 VSS.n2108 VSS.n9819 5.32359
R1599 VSS.n9818 VSS.t531 8.51132
R1600 VSS.t529 VSS.n9817 8.51132
R1601 VSS.t311 VSS.n9816 8.51132
R1602 VSS.t93 VSS.n9815 8.51132
R1603 VSS.n2108 VSS.n9814 5.32359
R1604 VSS.n2108 VSS.n9813 5.32359
R1605 VSS.n9812 VSS.t485 8.51132
R1606 VSS.n9811 VSS.t160 8.51132
R1607 VSS.n9810 VSS.t530 8.51132
R1608 VSS.n2108 VSS.n9809 5.32359
R1609 VSS.n9808 VSS.t420 8.51132
R1610 VSS.n9807 VSS.t162 8.51132
R1611 VSS.n9806 VSS.t430 8.51132
R1612 VSS.n9805 VSS.t602 8.51132
R1613 VSS.n9804 VSS.t333 8.51132
R1614 VSS.n9803 VSS.t48 8.51132
R1615 VSS.n2108 VSS.n9802 5.32359
R1616 VSS.n9801 VSS.t106 8.51132
R1617 VSS.t142 VSS.n9800 8.51132
R1618 VSS.t173 VSS.n9799 8.51132
R1619 VSS.t172 VSS.n9798 8.51132
R1620 VSS.n2108 VSS.n9797 5.32359
R1621 VSS.n2108 VSS.n9796 5.32359
R1622 VSS.n9795 VSS.t190 8.51132
R1623 VSS.n9794 VSS.t398 8.51132
R1624 VSS.n9793 VSS.t424 8.51132
R1625 VSS.n2108 VSS.n9792 5.32359
R1626 VSS.n9791 VSS.t437 8.51132
R1627 VSS.n9790 VSS.t537 8.51132
R1628 VSS.n9789 VSS.t171 8.51132
R1629 VSS.n9788 VSS.t402 8.51132
R1630 VSS.n9787 VSS.t572 8.51132
R1631 VSS.n9786 VSS.t412 8.51132
R1632 VSS.n2108 VSS.n9785 5.32359
R1633 VSS.n9784 VSS.t567 8.51132
R1634 VSS.t58 VSS.n9783 8.51132
R1635 VSS.t76 VSS.n9782 8.51132
R1636 VSS.t515 VSS.n9781 8.51132
R1637 VSS.n2108 VSS.n9780 5.32359
R1638 VSS.n2108 VSS.n9779 5.32359
R1639 VSS.n9778 VSS.t469 8.51132
R1640 VSS.n9777 VSS.t265 8.51132
R1641 VSS.n9776 VSS.t328 8.51132
R1642 VSS.n2108 VSS.n9775 5.32359
R1643 VSS.n9774 VSS.t123 8.51132
R1644 VSS.n9773 VSS.t283 8.51132
R1645 VSS.n9772 VSS.t609 8.51132
R1646 VSS.n9771 VSS.t492 8.51132
R1647 VSS.n9770 VSS.t69 8.51132
R1648 VSS.n9769 VSS.t302 8.51132
R1649 VSS.n2108 VSS.n9768 5.32359
R1650 VSS.n9767 VSS.t33 8.51132
R1651 VSS.t558 VSS.n9766 8.51132
R1652 VSS.t395 VSS.n9765 8.51132
R1653 VSS.t394 VSS.n9764 8.51132
R1654 VSS.n2108 VSS.n9763 5.32359
R1655 VSS.n2108 VSS.n9762 5.32359
R1656 VSS.n9761 VSS.t319 8.51132
R1657 VSS.n9760 VSS.t181 8.51132
R1658 VSS.n9759 VSS.t380 8.51132
R1659 VSS.n9665 VSS.n9666 0.2705
R1660 VSS.n9666 VSS.n9667 0.2705
R1661 VSS.n9667 VSS.n9668 0.2705
R1662 VSS.n9668 VSS.n9669 0.2705
R1663 VSS.n9669 VSS 0.3776
R1664 VSS VSS.n9670 0.1634
R1665 VSS.n9670 VSS.n9671 0.2705
R1666 VSS.n9671 VSS.n9672 0.2705
R1667 VSS.n9672 VSS.n9673 0.2705
R1668 VSS.n9673 VSS.n9674 0.2705
R1669 VSS.n9674 VSS.n9675 0.2705
R1670 VSS.n9675 VSS.n9676 0.30515
R1671 VSS.n9676 VSS.n9677 0.2705
R1672 VSS.n9677 VSS.n9678 0.2705
R1673 VSS.n9678 VSS.n9679 0.2705
R1674 VSS.n9679 VSS.n9680 0.2705
R1675 VSS.n9680 VSS.n9681 0.2705
R1676 VSS.n9681 VSS 0.3776
R1677 VSS VSS.n9682 0.1634
R1678 VSS.n9682 VSS.n9683 0.2705
R1679 VSS.n9683 VSS.n9684 0.2705
R1680 VSS.n9684 VSS.n9685 0.2705
R1681 VSS.n9685 VSS.n9686 0.2705
R1682 VSS.n9686 VSS.n9687 0.2705
R1683 VSS.n9687 VSS.n9688 0.30515
R1684 VSS.n9688 VSS.n9689 0.2705
R1685 VSS.n9689 VSS.n9690 0.2705
R1686 VSS.n9690 VSS.n9691 0.2705
R1687 VSS.n9691 VSS.n9692 0.2705
R1688 VSS.n9692 VSS.n9693 0.2705
R1689 VSS.n9693 VSS 0.3776
R1690 VSS VSS.n9694 0.1634
R1691 VSS.n9694 VSS.n9695 0.2705
R1692 VSS.n9695 VSS.n9696 0.2705
R1693 VSS.n9696 VSS.n9697 0.2705
R1694 VSS.n9697 VSS.n9698 0.2705
R1695 VSS.n9698 VSS.n9699 0.2705
R1696 VSS.n9699 VSS.n9700 0.30515
R1697 VSS.n9700 VSS.n9701 0.2705
R1698 VSS.n9701 VSS.n9702 0.2705
R1699 VSS.n9702 VSS.n9703 0.2705
R1700 VSS.n9703 VSS.n9704 0.2705
R1701 VSS.n9704 VSS.n9705 0.2705
R1702 VSS.n9705 VSS 0.3776
R1703 VSS VSS.n9706 0.1634
R1704 VSS.n9706 VSS.n9707 0.2705
R1705 VSS.n9707 VSS.n9708 0.2705
R1706 VSS.n9708 VSS.n9709 0.2705
R1707 VSS.n9709 VSS.n9710 0.2705
R1708 VSS.n9710 VSS.n9711 0.2705
R1709 VSS.n9711 VSS.n9712 0.30515
R1710 VSS.n9712 VSS.n9713 0.2705
R1711 VSS.n9713 VSS.n9714 0.2705
R1712 VSS.n9714 VSS.n9715 0.2705
R1713 VSS.n9715 VSS.n9716 0.2705
R1714 VSS.n9716 VSS.n9717 0.2705
R1715 VSS.n9717 VSS 0.3776
R1716 VSS VSS.n9718 0.1634
R1717 VSS.n9718 VSS.n9719 0.2705
R1718 VSS.n9719 VSS.n9720 0.2705
R1719 VSS.n9720 VSS.n9721 0.2705
R1720 VSS.n9721 VSS.n9722 0.2705
R1721 VSS.n9722 VSS.n9723 0.2705
R1722 VSS.n9723 VSS.n9724 0.30515
R1723 VSS.n9724 VSS.n9725 0.2705
R1724 VSS.n9725 VSS.n9726 0.2705
R1725 VSS.n9726 VSS.n9727 0.2705
R1726 VSS.n9727 VSS.n9728 0.2705
R1727 VSS.n9728 VSS.n9729 0.2705
R1728 VSS.n9729 VSS 0.3776
R1729 VSS VSS.n9730 0.1634
R1730 VSS.n9730 VSS.n9731 0.2705
R1731 VSS.n9731 VSS.n9732 0.2705
R1732 VSS.n9732 VSS.n9733 0.2705
R1733 VSS.n9733 VSS.n9734 0.2705
R1734 VSS.n9734 VSS.n9735 0.2705
R1735 VSS.n9735 VSS.n9736 0.30515
R1736 VSS.n9736 VSS.n9737 0.2705
R1737 VSS.n9737 VSS.n9738 0.2705
R1738 VSS.n9738 VSS.n9739 0.2705
R1739 VSS.n9739 VSS.n9740 0.2705
R1740 VSS.n9740 VSS.n9741 0.2705
R1741 VSS.n9741 VSS 0.3776
R1742 VSS VSS.n9742 0.1634
R1743 VSS.n9742 VSS.n9743 0.2705
R1744 VSS.n9743 VSS.n9744 0.2705
R1745 VSS.n9744 VSS.n9745 0.2705
R1746 VSS.n9745 VSS.n9746 0.2705
R1747 VSS.n9746 VSS.n9747 0.2705
R1748 VSS.n9747 VSS.n9748 0.30515
R1749 VSS.n9748 VSS.n9749 0.2705
R1750 VSS.n9749 VSS.n9750 0.2705
R1751 VSS.n9750 VSS.n9751 0.2705
R1752 VSS.n9751 VSS.n9752 0.2705
R1753 VSS.n9752 VSS.n9753 0.2705
R1754 VSS.n9753 VSS 0.3776
R1755 VSS VSS.n9754 0.1634
R1756 VSS.n9754 VSS.n9755 0.2705
R1757 VSS.n9755 VSS.n9756 0.2705
R1758 VSS.n9756 VSS.n9757 0.2705
R1759 VSS.n9757 VSS.n9758 0.2705
R1760 VSS.n9758 VSS.n9664 13.7705
R1761 VSS.n7170 VSS.n7171 0.0722544
R1762 VSS.n7172 VSS.n7173 4.5005
R1763 VSS.n7174 VSS.n7175 4.5005
R1764 VSS.n7176 VSS.n7177 4.5005
R1765 VSS.n7172 VSS.n7170 2.37296
R1766 VSS.n7174 VSS.n7172 0.127318
R1767 VSS.n7176 VSS.n7174 0.127318
R1768 VSS.t41 VSS.n7176 2.73618
R1769 VSS.n7171 VSS.n7178 4.5005
R1770 VSS.n7173 VSS.n7179 4.5005
R1771 VSS.n7175 VSS.n7180 4.5005
R1772 VSS.n7177 VSS.n7181 4.5005
R1773 VSS.n7183 VSS.n7170 4.647
R1774 VSS.n7171 VSS.n7173 0.147342
R1775 VSS.n7173 VSS.n7175 0.147342
R1776 VSS.n7175 VSS.n7177 0.147342
R1777 VSS.n7183 VSS.n7184 2.21488
R1778 VSS.n7178 VSS.n7183 0.0732424
R1779 VSS.n7182 VSS.n7184 2.21488
R1780 VSS.n7182 VSS.n7180 0.0732424
R1781 VSS.n7181 VSS.n7184 4.5005
R1782 VSS.n7178 VSS.n7179 0.147342
R1783 VSS.n7179 VSS.n7182 0.0732424
R1784 VSS.n7180 VSS.n7181 0.147342
R1785 VSS.n7185 VSS.n7186 4.5005
R1786 VSS.n7188 VSS.n7187 0.0732424
R1787 VSS.n7186 VSS.n7188 2.21488
R1788 VSS.n7191 VSS.n7190 0.0732424
R1789 VSS.n7186 VSS.n7191 2.21488
R1790 VSS.n7200 VSS.n7201 4.5005
R1791 VSS.n7203 VSS.n7202 0.0732424
R1792 VSS.n7201 VSS.n7203 2.21488
R1793 VSS.n7206 VSS.n7205 0.0732424
R1794 VSS.n7201 VSS.n7206 2.21488
R1795 VSS.n7215 VSS.n7216 4.5005
R1796 VSS.n7217 VSS.n7218 0.0732424
R1797 VSS.n7218 VSS.n7216 2.21488
R1798 VSS.n7220 VSS.n7221 0.0732424
R1799 VSS.n7221 VSS.n7216 2.21488
R1800 VSS.n7230 VSS.n7231 4.5005
R1801 VSS.n7233 VSS.n7232 0.0732424
R1802 VSS.n7231 VSS.n7233 2.21488
R1803 VSS.n7236 VSS.n7235 0.0732424
R1804 VSS.n7231 VSS.n7236 2.21488
R1805 VSS.n7245 VSS.n7246 4.5005
R1806 VSS.n7248 VSS.n7247 0.0732424
R1807 VSS.n7246 VSS.n7248 2.21488
R1808 VSS.n7251 VSS.n7250 0.0732424
R1809 VSS.n7246 VSS.n7251 2.21488
R1810 VSS.n7260 VSS.n7261 4.5005
R1811 VSS.n7263 VSS.n7262 0.0732424
R1812 VSS.n7261 VSS.n7263 2.21488
R1813 VSS.n7266 VSS.n7265 0.0732424
R1814 VSS.n7261 VSS.n7266 2.21488
R1815 VSS.n7275 VSS.n7276 4.5005
R1816 VSS.n7277 VSS.n7278 0.0732424
R1817 VSS.n7278 VSS.n7276 2.21488
R1818 VSS.n7280 VSS.n7281 0.0732424
R1819 VSS.n7281 VSS.n7276 2.21488
R1820 VSS.n7290 VSS.n7291 4.5005
R1821 VSS.n7293 VSS.n7292 0.0732424
R1822 VSS.n7291 VSS.n7293 2.21488
R1823 VSS.n7296 VSS.n7295 0.0732424
R1824 VSS.n7291 VSS.n7296 2.21488
R1825 VSS.n7305 VSS.n7306 4.5005
R1826 VSS.n7308 VSS.n7307 0.0732424
R1827 VSS.n7306 VSS.n7308 2.21488
R1828 VSS.n7311 VSS.n7310 0.0732424
R1829 VSS.n7306 VSS.n7311 2.21488
R1830 VSS.n7320 VSS.n7321 4.5005
R1831 VSS.n7323 VSS.n7322 0.0732424
R1832 VSS.n7321 VSS.n7323 2.21488
R1833 VSS.n7326 VSS.n7325 0.0732424
R1834 VSS.n7321 VSS.n7326 2.21488
R1835 VSS.n7335 VSS.n7336 4.5005
R1836 VSS.n7338 VSS.n7337 0.0732424
R1837 VSS.n7336 VSS.n7338 2.21488
R1838 VSS.n7341 VSS.n7340 0.0732424
R1839 VSS.n7336 VSS.n7341 2.21488
R1840 VSS.n7350 VSS.n7351 4.5005
R1841 VSS.n7353 VSS.n7352 0.0732424
R1842 VSS.n7351 VSS.n7353 2.21488
R1843 VSS.n7356 VSS.n7355 0.0732424
R1844 VSS.n7351 VSS.n7356 2.21488
R1845 VSS.n7365 VSS.n7366 4.5005
R1846 VSS.n7368 VSS.n7367 0.0732424
R1847 VSS.n7366 VSS.n7368 2.21488
R1848 VSS.n7371 VSS.n7370 0.0732424
R1849 VSS.n7366 VSS.n7371 2.21488
R1850 VSS.n7380 VSS.n7381 4.5005
R1851 VSS.n7382 VSS.n7383 0.0732424
R1852 VSS.n7383 VSS.n7381 2.21488
R1853 VSS.n7385 VSS.n7386 0.0732424
R1854 VSS.n7386 VSS.n7381 2.21488
R1855 VSS.n7395 VSS.n7396 4.5005
R1856 VSS.n7398 VSS.n7397 0.0732424
R1857 VSS.n7396 VSS.n7398 2.21488
R1858 VSS.n7401 VSS.n7400 0.0732424
R1859 VSS.n7396 VSS.n7401 2.21488
R1860 VSS.n7410 VSS.n7411 4.5005
R1861 VSS.n7413 VSS.n7412 0.0732424
R1862 VSS.n7411 VSS.n7413 2.21488
R1863 VSS.n7416 VSS.n7415 0.0732424
R1864 VSS.n7411 VSS.n7416 2.21488
R1865 VSS.n7425 VSS.n7426 4.5005
R1866 VSS.n7428 VSS.n7427 0.0732424
R1867 VSS.n7426 VSS.n7428 2.21488
R1868 VSS.n7431 VSS.n7430 0.0732424
R1869 VSS.n7426 VSS.n7431 2.21488
R1870 VSS.n7440 VSS.n7441 4.5005
R1871 VSS.n7442 VSS.n7443 0.0732424
R1872 VSS.n7443 VSS.n7441 2.21488
R1873 VSS.n7445 VSS.n7446 0.0732424
R1874 VSS.n7446 VSS.n7441 2.21488
R1875 VSS.n7455 VSS.n7456 4.5005
R1876 VSS.n7458 VSS.n7457 0.0732424
R1877 VSS.n7456 VSS.n7458 2.21488
R1878 VSS.n7461 VSS.n7460 0.0732424
R1879 VSS.n7456 VSS.n7461 2.21488
R1880 VSS.n7470 VSS.n7471 4.5005
R1881 VSS.n7473 VSS.n7472 0.0732424
R1882 VSS.n7471 VSS.n7473 2.21488
R1883 VSS.n7476 VSS.n7475 0.0732424
R1884 VSS.n7471 VSS.n7476 2.21488
R1885 VSS.n7485 VSS.n7486 4.5005
R1886 VSS.n7488 VSS.n7487 0.0732424
R1887 VSS.n7486 VSS.n7488 2.21488
R1888 VSS.n7491 VSS.n7490 0.0732424
R1889 VSS.n7486 VSS.n7491 2.21488
R1890 VSS.n7500 VSS.n7501 4.5005
R1891 VSS.n7503 VSS.n7502 0.0732424
R1892 VSS.n7501 VSS.n7503 2.21488
R1893 VSS.n7506 VSS.n7505 0.0732424
R1894 VSS.n7501 VSS.n7506 2.21488
R1895 VSS.n7515 VSS.n7516 4.5005
R1896 VSS.n7517 VSS.n7518 0.0732424
R1897 VSS.n7518 VSS.n7516 2.21488
R1898 VSS.n7520 VSS.n7521 0.0732424
R1899 VSS.n7521 VSS.n7516 2.21488
R1900 VSS.n7530 VSS.n7531 4.5005
R1901 VSS.n7533 VSS.n7532 0.0732424
R1902 VSS.n7531 VSS.n7533 2.21488
R1903 VSS.n7536 VSS.n7535 0.0732424
R1904 VSS.n7531 VSS.n7536 2.21488
R1905 VSS.n7545 VSS.n7546 4.5005
R1906 VSS.n7548 VSS.n7547 0.0732424
R1907 VSS.n7546 VSS.n7548 2.21488
R1908 VSS.n7551 VSS.n7550 0.0732424
R1909 VSS.n7546 VSS.n7551 2.21488
R1910 VSS.n7560 VSS.n7561 4.5005
R1911 VSS.n7563 VSS.n7562 0.0732424
R1912 VSS.n7561 VSS.n7563 2.21488
R1913 VSS.n7566 VSS.n7565 0.0732424
R1914 VSS.n7561 VSS.n7566 2.21488
R1915 VSS.n7575 VSS.n7576 4.5005
R1916 VSS.n7577 VSS.n7578 0.0732424
R1917 VSS.n7578 VSS.n7576 2.21488
R1918 VSS.n7580 VSS.n7581 0.0732424
R1919 VSS.n7581 VSS.n7576 2.21488
R1920 VSS.n7590 VSS.n7591 4.5005
R1921 VSS.n7593 VSS.n7592 0.0732424
R1922 VSS.n7591 VSS.n7593 2.21488
R1923 VSS.n7596 VSS.n7595 0.0732424
R1924 VSS.n7591 VSS.n7596 2.21488
R1925 VSS.n7605 VSS.n7606 4.5005
R1926 VSS.n7608 VSS.n7607 0.0732424
R1927 VSS.n7606 VSS.n7608 2.21488
R1928 VSS.n7611 VSS.n7610 0.0732424
R1929 VSS.n7606 VSS.n7611 2.21488
R1930 VSS.n7620 VSS.n7621 4.5005
R1931 VSS.n7623 VSS.n7622 0.0732424
R1932 VSS.n7621 VSS.n7623 2.21488
R1933 VSS.n7626 VSS.n7625 0.0732424
R1934 VSS.n7621 VSS.n7626 2.21488
R1935 VSS.n7635 VSS.n7636 4.5005
R1936 VSS.n7638 VSS.n7637 0.0732424
R1937 VSS.n7636 VSS.n7638 2.21488
R1938 VSS.n7641 VSS.n7640 0.0732424
R1939 VSS.n7636 VSS.n7641 2.21488
R1940 VSS.n7650 VSS.n7651 4.5005
R1941 VSS.n7653 VSS.n7652 0.0732424
R1942 VSS.n7651 VSS.n7653 2.21488
R1943 VSS.n7656 VSS.n7655 0.0732424
R1944 VSS.n7651 VSS.n7656 2.21488
R1945 VSS.n7665 VSS.n7666 4.5005
R1946 VSS.n7668 VSS.n7667 0.0732424
R1947 VSS.n7666 VSS.n7668 2.21488
R1948 VSS.n7671 VSS.n7670 0.0732424
R1949 VSS.n7666 VSS.n7671 2.21488
R1950 VSS.n7680 VSS.n7681 4.5005
R1951 VSS.n7682 VSS.n7683 0.0732424
R1952 VSS.n7683 VSS.n7681 2.21488
R1953 VSS.n7685 VSS.n7686 0.0732424
R1954 VSS.n7686 VSS.n7681 2.21488
R1955 VSS.n7695 VSS.n7696 4.5005
R1956 VSS.n7698 VSS.n7697 0.0732424
R1957 VSS.n7696 VSS.n7698 2.21488
R1958 VSS.n7701 VSS.n7700 0.0732424
R1959 VSS.n7696 VSS.n7701 2.21488
R1960 VSS.n7710 VSS.n7711 4.5005
R1961 VSS.n7713 VSS.n7712 0.0732424
R1962 VSS.n7711 VSS.n7713 2.21488
R1963 VSS.n7716 VSS.n7715 0.0732424
R1964 VSS.n7711 VSS.n7716 2.21488
R1965 VSS.n7725 VSS.n7726 4.5005
R1966 VSS.n7728 VSS.n7727 0.0732424
R1967 VSS.n7726 VSS.n7728 2.21488
R1968 VSS.n7731 VSS.n7730 0.0732424
R1969 VSS.n7726 VSS.n7731 2.21488
R1970 VSS.n7740 VSS.n7741 4.5005
R1971 VSS.n7742 VSS.n7743 0.0732424
R1972 VSS.n7743 VSS.n7741 2.21488
R1973 VSS.n7745 VSS.n7746 0.0732424
R1974 VSS.n7746 VSS.n7741 2.21488
R1975 VSS.n7755 VSS.n7756 4.5005
R1976 VSS.n7758 VSS.n7757 0.0732424
R1977 VSS.n7756 VSS.n7758 2.21488
R1978 VSS.n7761 VSS.n7760 0.0732424
R1979 VSS.n7756 VSS.n7761 2.21488
R1980 VSS.n7770 VSS.n7771 4.5005
R1981 VSS.n7773 VSS.n7772 0.0732424
R1982 VSS.n7771 VSS.n7773 2.21488
R1983 VSS.n7776 VSS.n7775 0.0732424
R1984 VSS.n7771 VSS.n7776 2.21488
R1985 VSS.n7785 VSS.n7786 4.5005
R1986 VSS.n7788 VSS.n7787 0.0732424
R1987 VSS.n7786 VSS.n7788 2.21488
R1988 VSS.n7791 VSS.n7790 0.0732424
R1989 VSS.n7786 VSS.n7791 2.21488
R1990 VSS.n7800 VSS.n7801 4.5005
R1991 VSS.n7803 VSS.n7802 0.0732424
R1992 VSS.n7801 VSS.n7803 2.21488
R1993 VSS.n7806 VSS.n7805 0.0732424
R1994 VSS.n7801 VSS.n7806 2.21488
R1995 VSS.n7815 VSS.n7816 4.5005
R1996 VSS.n7817 VSS.n7818 0.0732424
R1997 VSS.n7818 VSS.n7816 2.21488
R1998 VSS.n7820 VSS.n7821 0.0732424
R1999 VSS.n7821 VSS.n7816 2.21488
R2000 VSS.n7830 VSS.n7831 4.5005
R2001 VSS.n7833 VSS.n7832 0.0732424
R2002 VSS.n7831 VSS.n7833 2.21488
R2003 VSS.n7836 VSS.n7835 0.0732424
R2004 VSS.n7831 VSS.n7836 2.21488
R2005 VSS.n7845 VSS.n7846 4.5005
R2006 VSS.n7848 VSS.n7847 0.0732424
R2007 VSS.n7846 VSS.n7848 2.21488
R2008 VSS.n7851 VSS.n7850 0.0732424
R2009 VSS.n7846 VSS.n7851 2.21488
R2010 VSS.n7860 VSS.n7861 4.5005
R2011 VSS.n7863 VSS.n7862 0.0732424
R2012 VSS.n7861 VSS.n7863 2.21488
R2013 VSS.n7866 VSS.n7865 0.0732424
R2014 VSS.n7861 VSS.n7866 2.21488
R2015 VSS.n7875 VSS.n7876 4.5005
R2016 VSS.n7877 VSS.n7878 0.0732424
R2017 VSS.n7878 VSS.n7876 2.21488
R2018 VSS.n7880 VSS.n7881 0.0732424
R2019 VSS.n7881 VSS.n7876 2.21488
R2020 VSS.n7890 VSS.n7891 4.5005
R2021 VSS.n7893 VSS.n7892 0.0732424
R2022 VSS.n7891 VSS.n7893 2.21488
R2023 VSS.n7896 VSS.n7895 0.0732424
R2024 VSS.n7891 VSS.n7896 2.21488
R2025 VSS.n7905 VSS.n7906 4.5005
R2026 VSS.n7908 VSS.n7907 0.0732424
R2027 VSS.n7906 VSS.n7908 2.21488
R2028 VSS.n7911 VSS.n7910 0.0732424
R2029 VSS.n7906 VSS.n7911 2.21488
R2030 VSS.n7920 VSS.n7921 4.5005
R2031 VSS.n7923 VSS.n7922 0.0732424
R2032 VSS.n7921 VSS.n7923 2.21488
R2033 VSS.n7926 VSS.n7925 0.0732424
R2034 VSS.n7921 VSS.n7926 2.21488
R2035 VSS.n7935 VSS.n7936 4.5005
R2036 VSS.n7938 VSS.n7937 0.0732424
R2037 VSS.n7936 VSS.n7938 2.21488
R2038 VSS.n7941 VSS.n7940 0.0732424
R2039 VSS.n7936 VSS.n7941 2.21488
R2040 VSS.n7950 VSS.n7951 4.5005
R2041 VSS.n7953 VSS.n7952 0.0732424
R2042 VSS.n7951 VSS.n7953 2.21488
R2043 VSS.n7956 VSS.n7955 0.0732424
R2044 VSS.n7951 VSS.n7956 2.21488
R2045 VSS.n7965 VSS.n7966 4.5005
R2046 VSS.n7968 VSS.n7967 0.0732424
R2047 VSS.n7966 VSS.n7968 2.21488
R2048 VSS.n7971 VSS.n7970 0.0732424
R2049 VSS.n7966 VSS.n7971 2.21488
R2050 VSS.n7980 VSS.n7981 4.5005
R2051 VSS.n7982 VSS.n7983 0.0732424
R2052 VSS.n7983 VSS.n7981 2.21488
R2053 VSS.n7985 VSS.n7986 0.0732424
R2054 VSS.n7986 VSS.n7981 2.21488
R2055 VSS.n7995 VSS.n7996 4.5005
R2056 VSS.n7998 VSS.n7997 0.0732424
R2057 VSS.n7996 VSS.n7998 2.21488
R2058 VSS.n8001 VSS.n8000 0.0732424
R2059 VSS.n7996 VSS.n8001 2.21488
R2060 VSS.n8010 VSS.n8011 4.5005
R2061 VSS.n8013 VSS.n8012 0.0732424
R2062 VSS.n8011 VSS.n8013 2.21488
R2063 VSS.n8016 VSS.n8015 0.0732424
R2064 VSS.n8011 VSS.n8016 2.21488
R2065 VSS.n8025 VSS.n8026 4.5005
R2066 VSS.n8028 VSS.n8027 0.0732424
R2067 VSS.n8026 VSS.n8028 2.21488
R2068 VSS.n8031 VSS.n8030 0.0732424
R2069 VSS.n8026 VSS.n8031 2.21488
R2070 VSS.n8040 VSS.n8041 4.5005
R2071 VSS.n8042 VSS.n8043 0.0732424
R2072 VSS.n8043 VSS.n8041 2.21488
R2073 VSS.n8045 VSS.n8046 0.0732424
R2074 VSS.n8046 VSS.n8041 2.21488
R2075 VSS.n8055 VSS.n8056 4.5005
R2076 VSS.n8058 VSS.n8057 0.0732424
R2077 VSS.n8056 VSS.n8058 2.21488
R2078 VSS.n8061 VSS.n8060 0.0732424
R2079 VSS.n8056 VSS.n8061 2.21488
R2080 VSS.n8070 VSS.n8071 4.5005
R2081 VSS.n8073 VSS.n8072 0.0732424
R2082 VSS.n8071 VSS.n8073 2.21488
R2083 VSS.n8076 VSS.n8075 0.0732424
R2084 VSS.n8071 VSS.n8076 2.21488
R2085 VSS.n8085 VSS.n8086 4.5005
R2086 VSS.n8088 VSS.n8087 0.0732424
R2087 VSS.n8086 VSS.n8088 2.21488
R2088 VSS.n8091 VSS.n8090 0.0732424
R2089 VSS.n8086 VSS.n8091 2.21488
R2090 VSS.n8100 VSS.n8101 4.5005
R2091 VSS.n8103 VSS.n8102 0.0732424
R2092 VSS.n8101 VSS.n8103 2.21488
R2093 VSS.n8106 VSS.n8105 0.0732424
R2094 VSS.n8101 VSS.n8106 2.21488
R2095 VSS.n8115 VSS.n8116 4.5005
R2096 VSS.n8117 VSS.n8118 0.0732424
R2097 VSS.n8118 VSS.n8116 2.21488
R2098 VSS.n8120 VSS.n8121 0.0732424
R2099 VSS.n8121 VSS.n8116 2.21488
R2100 VSS.n8130 VSS.n8131 4.5005
R2101 VSS.n8133 VSS.n8132 0.0732424
R2102 VSS.n8131 VSS.n8133 2.21488
R2103 VSS.n8136 VSS.n8135 0.0732424
R2104 VSS.n8131 VSS.n8136 2.21488
R2105 VSS.n8145 VSS.n8146 4.5005
R2106 VSS.n8148 VSS.n8147 0.0732424
R2107 VSS.n8146 VSS.n8148 2.21488
R2108 VSS.n8151 VSS.n8150 0.0732424
R2109 VSS.n8146 VSS.n8151 2.21488
R2110 VSS.n8160 VSS.n8161 4.5005
R2111 VSS.n8163 VSS.n8162 0.0732424
R2112 VSS.n8161 VSS.n8163 2.21488
R2113 VSS.n8166 VSS.n8165 0.0732424
R2114 VSS.n8161 VSS.n8166 2.21488
R2115 VSS.n8175 VSS.n8176 4.5005
R2116 VSS.n8177 VSS.n8178 0.0732424
R2117 VSS.n8178 VSS.n8176 2.21488
R2118 VSS.n8180 VSS.n8181 0.0732424
R2119 VSS.n8181 VSS.n8176 2.21488
R2120 VSS.n8190 VSS.n8191 4.5005
R2121 VSS.n8193 VSS.n8192 0.0732424
R2122 VSS.n8191 VSS.n8193 2.21488
R2123 VSS.n8196 VSS.n8195 0.0732424
R2124 VSS.n8191 VSS.n8196 2.21488
R2125 VSS.n8205 VSS.n8206 4.5005
R2126 VSS.n8208 VSS.n8207 0.0732424
R2127 VSS.n8206 VSS.n8208 2.21488
R2128 VSS.n8211 VSS.n8210 0.0732424
R2129 VSS.n8206 VSS.n8211 2.21488
R2130 VSS.n8220 VSS.n8221 4.5005
R2131 VSS.n8223 VSS.n8222 0.0732424
R2132 VSS.n8221 VSS.n8223 2.21488
R2133 VSS.n8226 VSS.n8225 0.0732424
R2134 VSS.n8221 VSS.n8226 2.21488
R2135 VSS.n8235 VSS.n8236 4.5005
R2136 VSS.n8238 VSS.n8237 0.0732424
R2137 VSS.n8236 VSS.n8238 2.21488
R2138 VSS.n8241 VSS.n8240 0.0732424
R2139 VSS.n8236 VSS.n8241 2.21488
R2140 VSS.n8250 VSS.n8251 4.5005
R2141 VSS.n8253 VSS.n8252 0.0732424
R2142 VSS.n8251 VSS.n8253 2.21488
R2143 VSS.n8256 VSS.n8255 0.0732424
R2144 VSS.n8251 VSS.n8256 2.21488
R2145 VSS.n8265 VSS.n8266 4.5005
R2146 VSS.n8268 VSS.n8267 0.0732424
R2147 VSS.n8266 VSS.n8268 2.21488
R2148 VSS.n8271 VSS.n8270 0.0732424
R2149 VSS.n8266 VSS.n8271 2.21488
R2150 VSS.n8280 VSS.n8281 4.5005
R2151 VSS.n8282 VSS.n8283 0.0732424
R2152 VSS.n8283 VSS.n8281 2.21488
R2153 VSS.n8285 VSS.n8286 0.0732424
R2154 VSS.n8286 VSS.n8281 2.21488
R2155 VSS.n8295 VSS.n8296 4.5005
R2156 VSS.n8298 VSS.n8297 0.0732424
R2157 VSS.n8296 VSS.n8298 2.21488
R2158 VSS.n8301 VSS.n8300 0.0732424
R2159 VSS.n8296 VSS.n8301 2.21488
R2160 VSS.n8310 VSS.n8311 4.5005
R2161 VSS.n8313 VSS.n8312 0.0732424
R2162 VSS.n8311 VSS.n8313 2.21488
R2163 VSS.n8316 VSS.n8315 0.0732424
R2164 VSS.n8311 VSS.n8316 2.21488
R2165 VSS.n8325 VSS.n8326 4.5005
R2166 VSS.n8328 VSS.n8327 0.0732424
R2167 VSS.n8326 VSS.n8328 2.21488
R2168 VSS.n8331 VSS.n8330 0.0732424
R2169 VSS.n8326 VSS.n8331 2.21488
R2170 VSS.n8340 VSS.n8341 4.5005
R2171 VSS.n8342 VSS.n8343 0.0732424
R2172 VSS.n8343 VSS.n8341 2.21488
R2173 VSS.n8345 VSS.n8346 0.0732424
R2174 VSS.n8346 VSS.n8341 2.21488
R2175 VSS.n8355 VSS.n8356 4.5005
R2176 VSS.n8358 VSS.n8357 0.0732424
R2177 VSS.n8356 VSS.n8358 2.21488
R2178 VSS.n8361 VSS.n8360 0.0732424
R2179 VSS.n8356 VSS.n8361 2.21488
R2180 VSS.n8370 VSS.n8371 4.5005
R2181 VSS.n8373 VSS.n8372 0.0732424
R2182 VSS.n8371 VSS.n8373 2.21488
R2183 VSS.n8376 VSS.n8375 0.0732424
R2184 VSS.n8371 VSS.n8376 2.21488
R2185 VSS.n8385 VSS.n8386 4.5005
R2186 VSS.n8388 VSS.n8387 0.0732424
R2187 VSS.n8386 VSS.n8388 2.21488
R2188 VSS.n8391 VSS.n8390 0.0732424
R2189 VSS.n8386 VSS.n8391 2.21488
R2190 VSS.n8400 VSS.n8401 4.5005
R2191 VSS.n8403 VSS.n8402 0.0732424
R2192 VSS.n8401 VSS.n8403 2.21488
R2193 VSS.n8406 VSS.n8405 0.0732424
R2194 VSS.n8401 VSS.n8406 2.21488
R2195 VSS.n8415 VSS.n8416 4.5005
R2196 VSS.n8417 VSS.n8418 0.0732424
R2197 VSS.n8418 VSS.n8416 2.21488
R2198 VSS.n8420 VSS.n8421 0.0732424
R2199 VSS.n8421 VSS.n8416 2.21488
R2200 VSS.n8430 VSS.n8431 4.5005
R2201 VSS.n8433 VSS.n8432 0.0732424
R2202 VSS.n8431 VSS.n8433 2.21488
R2203 VSS.n8436 VSS.n8435 0.0732424
R2204 VSS.n8431 VSS.n8436 2.21488
R2205 VSS.n8445 VSS.n8446 4.5005
R2206 VSS.n8448 VSS.n8447 0.0732424
R2207 VSS.n8446 VSS.n8448 2.21488
R2208 VSS.n8451 VSS.n8450 0.0732424
R2209 VSS.n8446 VSS.n8451 2.21488
R2210 VSS.n8460 VSS.n8461 4.5005
R2211 VSS.n8463 VSS.n8462 0.0732424
R2212 VSS.n8461 VSS.n8463 2.21488
R2213 VSS.n8466 VSS.n8465 0.0732424
R2214 VSS.n8461 VSS.n8466 2.21488
R2215 VSS.n8475 VSS.n8476 4.5005
R2216 VSS.n8477 VSS.n8478 0.0732424
R2217 VSS.n8478 VSS.n8476 2.21488
R2218 VSS.n8480 VSS.n8481 0.0732424
R2219 VSS.n8481 VSS.n8476 2.21488
R2220 VSS.n8490 VSS.n8491 4.5005
R2221 VSS.n8493 VSS.n8492 0.0732424
R2222 VSS.n8491 VSS.n8493 2.21488
R2223 VSS.n8496 VSS.n8495 0.0732424
R2224 VSS.n8491 VSS.n8496 2.21488
R2225 VSS.n8505 VSS.n8506 4.5005
R2226 VSS.n8508 VSS.n8507 0.0732424
R2227 VSS.n8506 VSS.n8508 2.21488
R2228 VSS.n8511 VSS.n8510 0.0732424
R2229 VSS.n8506 VSS.n8511 2.21488
R2230 VSS.n8520 VSS.n8521 4.5005
R2231 VSS.n8523 VSS.n8522 0.0732424
R2232 VSS.n8521 VSS.n8523 2.21488
R2233 VSS.n8526 VSS.n8525 0.0732424
R2234 VSS.n8521 VSS.n8526 2.21488
R2235 VSS.n8535 VSS.n8536 4.5005
R2236 VSS.n8538 VSS.n8537 0.0732424
R2237 VSS.n8536 VSS.n8538 2.21488
R2238 VSS.n8541 VSS.n8540 0.0732424
R2239 VSS.n8536 VSS.n8541 2.21488
R2240 VSS.n8550 VSS.n8551 4.5005
R2241 VSS.n8553 VSS.n8552 0.0732424
R2242 VSS.n8551 VSS.n8553 2.21488
R2243 VSS.n8556 VSS.n8555 0.0732424
R2244 VSS.n8551 VSS.n8556 2.21488
R2245 VSS.n8565 VSS.n8566 4.5005
R2246 VSS.n8568 VSS.n8567 0.0732424
R2247 VSS.n8566 VSS.n8568 2.21488
R2248 VSS.n8571 VSS.n8570 0.0732424
R2249 VSS.n8566 VSS.n8571 2.21488
R2250 VSS.n8580 VSS.n8581 4.5005
R2251 VSS.n8582 VSS.n8583 0.0732424
R2252 VSS.n8583 VSS.n8581 2.21488
R2253 VSS.n8585 VSS.n8586 0.0732424
R2254 VSS.n8586 VSS.n8581 2.21488
R2255 VSS.n8595 VSS.n8596 4.5005
R2256 VSS.n8598 VSS.n8597 0.0732424
R2257 VSS.n8596 VSS.n8598 2.21488
R2258 VSS.n8601 VSS.n8600 0.0732424
R2259 VSS.n8596 VSS.n8601 2.21488
R2260 VSS.n8610 VSS.n8611 4.5005
R2261 VSS.n8613 VSS.n8612 0.0732424
R2262 VSS.n8611 VSS.n8613 2.21488
R2263 VSS.n8616 VSS.n8615 0.0732424
R2264 VSS.n8611 VSS.n8616 2.21488
R2265 VSS.n8625 VSS.n8626 4.5005
R2266 VSS.n8628 VSS.n8627 0.0732424
R2267 VSS.n8626 VSS.n8628 2.21488
R2268 VSS.n8631 VSS.n8630 0.0732424
R2269 VSS.n8626 VSS.n8631 2.21488
R2270 VSS.n8640 VSS.n8641 4.5005
R2271 VSS.n8642 VSS.n8643 0.0732424
R2272 VSS.n8643 VSS.n8641 2.21488
R2273 VSS.n8645 VSS.n8646 0.0732424
R2274 VSS.n8646 VSS.n8641 2.21488
R2275 VSS.n8655 VSS.n8656 4.5005
R2276 VSS.n8658 VSS.n8657 0.0732424
R2277 VSS.n8656 VSS.n8658 2.21488
R2278 VSS.n8661 VSS.n8660 0.0732424
R2279 VSS.n8656 VSS.n8661 2.21488
R2280 VSS.n8670 VSS.n8671 4.5005
R2281 VSS.n8673 VSS.n8672 0.0732424
R2282 VSS.n8671 VSS.n8673 2.21488
R2283 VSS.n8676 VSS.n8675 0.0732424
R2284 VSS.n8671 VSS.n8676 2.21488
R2285 VSS.n8685 VSS.n8686 4.5005
R2286 VSS.n8688 VSS.n8687 0.0732424
R2287 VSS.n8686 VSS.n8688 2.21488
R2288 VSS.n8691 VSS.n8690 0.0732424
R2289 VSS.n8686 VSS.n8691 2.21488
R2290 VSS.n8700 VSS.n8701 4.5005
R2291 VSS.n8703 VSS.n8702 0.0732424
R2292 VSS.n8701 VSS.n8703 2.21488
R2293 VSS.n8706 VSS.n8705 0.0732424
R2294 VSS.n8701 VSS.n8706 2.21488
R2295 VSS.n8715 VSS.n8716 4.5005
R2296 VSS.n8717 VSS.n8718 0.0732424
R2297 VSS.n8718 VSS.n8716 2.21488
R2298 VSS.n8720 VSS.n8721 0.0732424
R2299 VSS.n8721 VSS.n8716 2.21488
R2300 VSS.n8730 VSS.n8731 4.5005
R2301 VSS.n8733 VSS.n8732 0.0732424
R2302 VSS.n8731 VSS.n8733 2.21488
R2303 VSS.n8736 VSS.n8735 0.0732424
R2304 VSS.n8731 VSS.n8736 2.21488
R2305 VSS.n8745 VSS.n8746 4.5005
R2306 VSS.n8748 VSS.n8747 0.0732424
R2307 VSS.n8746 VSS.n8748 2.21488
R2308 VSS.n8751 VSS.n8750 0.0732424
R2309 VSS.n8746 VSS.n8751 2.21488
R2310 VSS.n8760 VSS.n8761 4.5005
R2311 VSS.n8763 VSS.n8762 0.0732424
R2312 VSS.n8761 VSS.n8763 2.21488
R2313 VSS.n8766 VSS.n8765 0.0732424
R2314 VSS.n8761 VSS.n8766 2.21488
R2315 VSS.n8775 VSS.n8776 4.5005
R2316 VSS.n8777 VSS.n8778 0.0732424
R2317 VSS.n8778 VSS.n8776 2.21488
R2318 VSS.n8780 VSS.n8781 0.0732424
R2319 VSS.n8781 VSS.n8776 2.21488
R2320 VSS.n8790 VSS.n8791 4.5005
R2321 VSS.n8793 VSS.n8792 0.0732424
R2322 VSS.n8791 VSS.n8793 2.21488
R2323 VSS.n8796 VSS.n8795 0.0732424
R2324 VSS.n8791 VSS.n8796 2.21488
R2325 VSS.n8805 VSS.n8806 4.5005
R2326 VSS.n8808 VSS.n8807 0.0732424
R2327 VSS.n8806 VSS.n8808 2.21488
R2328 VSS.n8811 VSS.n8810 0.0732424
R2329 VSS.n8806 VSS.n8811 2.21488
R2330 VSS.n8820 VSS.n8821 4.5005
R2331 VSS.n8823 VSS.n8822 0.0732424
R2332 VSS.n8821 VSS.n8823 2.21488
R2333 VSS.n8826 VSS.n8825 0.0732424
R2334 VSS.n8821 VSS.n8826 2.21488
R2335 VSS.n8835 VSS.n8836 4.5005
R2336 VSS.n8838 VSS.n8837 0.0732424
R2337 VSS.n8836 VSS.n8838 2.21488
R2338 VSS.n8841 VSS.n8840 0.0732424
R2339 VSS.n8836 VSS.n8841 2.21488
R2340 VSS.n8850 VSS.n8851 4.5005
R2341 VSS.n8853 VSS.n8852 0.0732424
R2342 VSS.n8851 VSS.n8853 2.21488
R2343 VSS.n8856 VSS.n8855 0.0732424
R2344 VSS.n8851 VSS.n8856 2.21488
R2345 VSS.n8865 VSS.n8866 4.5005
R2346 VSS.n8868 VSS.n8867 0.0732424
R2347 VSS.n8866 VSS.n8868 2.21488
R2348 VSS.n8871 VSS.n8870 0.0732424
R2349 VSS.n8866 VSS.n8871 2.21488
R2350 VSS.n8880 VSS.n8881 4.5005
R2351 VSS.n8882 VSS.n8883 0.0732424
R2352 VSS.n8883 VSS.n8881 2.21488
R2353 VSS.n8885 VSS.n8886 0.0732424
R2354 VSS.n8886 VSS.n8881 2.21488
R2355 VSS.n8895 VSS.n8896 4.5005
R2356 VSS.n8898 VSS.n8897 0.0732424
R2357 VSS.n8896 VSS.n8898 2.21488
R2358 VSS.n8901 VSS.n8900 0.0732424
R2359 VSS.n8896 VSS.n8901 2.21488
R2360 VSS.n8910 VSS.n8911 4.5005
R2361 VSS.n8913 VSS.n8912 0.0732424
R2362 VSS.n8911 VSS.n8913 2.21488
R2363 VSS.n8916 VSS.n8915 0.0732424
R2364 VSS.n8911 VSS.n8916 2.21488
R2365 VSS.n8925 VSS.n8926 4.5005
R2366 VSS.n8928 VSS.n8927 0.0732424
R2367 VSS.n8926 VSS.n8928 2.21488
R2368 VSS.n8931 VSS.n8930 0.0732424
R2369 VSS.n8926 VSS.n8931 2.21488
R2370 VSS.n8940 VSS.n8941 4.5005
R2371 VSS.n8942 VSS.n8943 0.0732424
R2372 VSS.n8943 VSS.n8941 2.21488
R2373 VSS.n8945 VSS.n8946 0.0732424
R2374 VSS.n8946 VSS.n8941 2.21488
R2375 VSS.n8955 VSS.n8956 4.5005
R2376 VSS.n8958 VSS.n8957 0.0732424
R2377 VSS.n8956 VSS.n8958 2.21488
R2378 VSS.n8961 VSS.n8960 0.0732424
R2379 VSS.n8956 VSS.n8961 2.21488
R2380 VSS.n8970 VSS.n8971 4.5005
R2381 VSS.n8973 VSS.n8972 0.0732424
R2382 VSS.n8971 VSS.n8973 2.21488
R2383 VSS.n8976 VSS.n8975 0.0732424
R2384 VSS.n8971 VSS.n8976 2.21488
R2385 VSS.n8985 VSS.n8986 4.5005
R2386 VSS.n8988 VSS.n8987 0.0732424
R2387 VSS.n8986 VSS.n8988 2.21488
R2388 VSS.n8991 VSS.n8990 0.0732424
R2389 VSS.n8986 VSS.n8991 2.21488
R2390 VSS.n9000 VSS.n9001 4.5005
R2391 VSS.n9003 VSS.n9002 0.0732424
R2392 VSS.n9001 VSS.n9003 2.21488
R2393 VSS.n9006 VSS.n9005 0.0732424
R2394 VSS.n9001 VSS.n9006 2.21488
R2395 VSS.n9015 VSS.n9016 4.5005
R2396 VSS.n9017 VSS.n9018 0.0732424
R2397 VSS.n9018 VSS.n9016 2.21488
R2398 VSS.n9020 VSS.n9021 0.0732424
R2399 VSS.n9021 VSS.n9016 2.21488
R2400 VSS.n9030 VSS.n9031 4.5005
R2401 VSS.n9033 VSS.n9032 0.0732424
R2402 VSS.n9031 VSS.n9033 2.21488
R2403 VSS.n9036 VSS.n9035 0.0732424
R2404 VSS.n9031 VSS.n9036 2.21488
R2405 VSS.n9045 VSS.n9046 4.5005
R2406 VSS.n9048 VSS.n9047 0.0732424
R2407 VSS.n9046 VSS.n9048 2.21488
R2408 VSS.n9051 VSS.n9050 0.0732424
R2409 VSS.n9046 VSS.n9051 2.21488
R2410 VSS.n9060 VSS.n9061 4.5005
R2411 VSS.n9063 VSS.n9062 0.0732424
R2412 VSS.n9061 VSS.n9063 2.21488
R2413 VSS.n9066 VSS.n9065 0.0732424
R2414 VSS.n9061 VSS.n9066 2.21488
R2415 VSS.n9075 VSS.n9076 4.5005
R2416 VSS.n9077 VSS.n9078 0.0732424
R2417 VSS.n9078 VSS.n9076 2.21488
R2418 VSS.n9080 VSS.n9081 0.0732424
R2419 VSS.n9081 VSS.n9076 2.21488
R2420 VSS.n9090 VSS.n9091 4.5005
R2421 VSS.n9093 VSS.n9092 0.0732424
R2422 VSS.n9091 VSS.n9093 2.21488
R2423 VSS.n9096 VSS.n9095 0.0732424
R2424 VSS.n9091 VSS.n9096 2.21488
R2425 VSS.n9105 VSS.n9106 4.5005
R2426 VSS.n9108 VSS.n9107 0.0732424
R2427 VSS.n9106 VSS.n9108 2.21488
R2428 VSS.n9111 VSS.n9110 0.0732424
R2429 VSS.n9106 VSS.n9111 2.21488
R2430 VSS.n9120 VSS.n9121 4.5005
R2431 VSS.n9123 VSS.n9122 0.0732424
R2432 VSS.n9121 VSS.n9123 2.21488
R2433 VSS.n9126 VSS.n9125 0.0732424
R2434 VSS.n9121 VSS.n9126 2.21488
R2435 VSS.n9135 VSS.n9136 4.5005
R2436 VSS.n9138 VSS.n9137 0.0732424
R2437 VSS.n9136 VSS.n9138 2.21488
R2438 VSS.n9141 VSS.n9140 0.0732424
R2439 VSS.n9136 VSS.n9141 2.21488
R2440 VSS.n9150 VSS.n9151 4.5005
R2441 VSS.n9153 VSS.n9152 0.0732424
R2442 VSS.n9151 VSS.n9153 2.21488
R2443 VSS.n9156 VSS.n9155 0.0732424
R2444 VSS.n9151 VSS.n9156 2.21488
R2445 VSS.n9165 VSS.n9166 4.5005
R2446 VSS.n9168 VSS.n9167 0.0732424
R2447 VSS.n9166 VSS.n9168 2.21488
R2448 VSS.n9171 VSS.n9170 0.0732424
R2449 VSS.n9166 VSS.n9171 2.21488
R2450 VSS.n9180 VSS.n9181 4.5005
R2451 VSS.n9182 VSS.n9183 0.0732424
R2452 VSS.n9183 VSS.n9181 2.21488
R2453 VSS.n9185 VSS.n9186 0.0732424
R2454 VSS.n9186 VSS.n9181 2.21488
R2455 VSS.n9195 VSS.n9196 4.5005
R2456 VSS.n9198 VSS.n9197 0.0732424
R2457 VSS.n9196 VSS.n9198 2.21488
R2458 VSS.n9201 VSS.n9200 0.0732424
R2459 VSS.n9196 VSS.n9201 2.21488
R2460 VSS.n9210 VSS.n9211 4.5005
R2461 VSS.n9213 VSS.n9212 0.0732424
R2462 VSS.n9211 VSS.n9213 2.21488
R2463 VSS.n9216 VSS.n9215 0.0732424
R2464 VSS.n9211 VSS.n9216 2.21488
R2465 VSS.n9225 VSS.n9226 4.5005
R2466 VSS.n9228 VSS.n9227 0.0732424
R2467 VSS.n9226 VSS.n9228 2.21488
R2468 VSS.n9231 VSS.n9230 0.0732424
R2469 VSS.n9226 VSS.n9231 2.21488
R2470 VSS.n9240 VSS.n9241 4.5005
R2471 VSS.n9242 VSS.n9243 0.0732424
R2472 VSS.n9243 VSS.n9241 2.21488
R2473 VSS.n9245 VSS.n9246 0.0732424
R2474 VSS.n9246 VSS.n9241 2.21488
R2475 VSS.n9255 VSS.n9256 4.5005
R2476 VSS.n9258 VSS.n9257 0.0732424
R2477 VSS.n9256 VSS.n9258 2.21488
R2478 VSS.n9261 VSS.n9260 0.0732424
R2479 VSS.n9256 VSS.n9261 2.21488
R2480 VSS.n9270 VSS.n9271 4.5005
R2481 VSS.n9273 VSS.n9272 0.0732424
R2482 VSS.n9271 VSS.n9273 2.21488
R2483 VSS.n9276 VSS.n9275 0.0732424
R2484 VSS.n9271 VSS.n9276 2.21488
R2485 VSS.n9285 VSS.n9286 4.5005
R2486 VSS.n9288 VSS.n9287 0.0732424
R2487 VSS.n9286 VSS.n9288 2.21488
R2488 VSS.n9291 VSS.n9290 0.0732424
R2489 VSS.n9286 VSS.n9291 2.21488
R2490 VSS.n9300 VSS.n9301 4.5005
R2491 VSS.n9303 VSS.n9302 0.0732424
R2492 VSS.n9301 VSS.n9303 2.21488
R2493 VSS.n9306 VSS.n9305 0.0732424
R2494 VSS.n9301 VSS.n9306 2.21488
R2495 VSS.n9315 VSS.n9316 4.5005
R2496 VSS.n9317 VSS.n9318 0.0732424
R2497 VSS.n9318 VSS.n9316 2.21488
R2498 VSS.n9320 VSS.n9321 0.0732424
R2499 VSS.n9321 VSS.n9316 2.21488
R2500 VSS.n9330 VSS.n9331 4.5005
R2501 VSS.n9333 VSS.n9332 0.0732424
R2502 VSS.n9331 VSS.n9333 2.21488
R2503 VSS.n9336 VSS.n9335 0.0732424
R2504 VSS.n9331 VSS.n9336 2.21488
R2505 VSS.n9345 VSS.n9346 4.5005
R2506 VSS.n9348 VSS.n9347 0.0732424
R2507 VSS.n9346 VSS.n9348 2.21488
R2508 VSS.n9351 VSS.n9350 0.0732424
R2509 VSS.n9346 VSS.n9351 2.21488
R2510 VSS.n9360 VSS.n9361 4.5005
R2511 VSS.n9363 VSS.n9362 0.0732424
R2512 VSS.n9361 VSS.n9363 2.21488
R2513 VSS.n9366 VSS.n9365 0.0732424
R2514 VSS.n9361 VSS.n9366 2.21488
R2515 VSS.n9375 VSS.n9376 4.5005
R2516 VSS.n9377 VSS.n9378 0.0732424
R2517 VSS.n9378 VSS.n9376 2.21488
R2518 VSS.n9380 VSS.n9381 0.0732424
R2519 VSS.n9381 VSS.n9376 2.21488
R2520 VSS.n9390 VSS.n9391 4.5005
R2521 VSS.n9393 VSS.n9392 0.0732424
R2522 VSS.n9391 VSS.n9393 2.21488
R2523 VSS.n9396 VSS.n9395 0.0732424
R2524 VSS.n9391 VSS.n9396 2.21488
R2525 VSS.n9405 VSS.n9406 4.5005
R2526 VSS.n9408 VSS.n9407 0.0732424
R2527 VSS.n9406 VSS.n9408 2.21488
R2528 VSS.n9411 VSS.n9410 0.0732424
R2529 VSS.n9406 VSS.n9411 2.21488
R2530 VSS.n9420 VSS.n9421 4.5005
R2531 VSS.n9423 VSS.n9422 0.0732424
R2532 VSS.n9421 VSS.n9423 2.21488
R2533 VSS.n9426 VSS.n9425 0.0732424
R2534 VSS.n9421 VSS.n9426 2.21488
R2535 VSS.n9435 VSS.n9436 4.5005
R2536 VSS.n9438 VSS.n9437 0.0732424
R2537 VSS.n9436 VSS.n9438 2.21488
R2538 VSS.n9441 VSS.n9440 0.0732424
R2539 VSS.n9436 VSS.n9441 2.21488
R2540 VSS.n9450 VSS.n9451 4.5005
R2541 VSS.n9453 VSS.n9452 0.0732424
R2542 VSS.n9451 VSS.n9453 2.21488
R2543 VSS.n9456 VSS.n9455 0.0732424
R2544 VSS.n9451 VSS.n9456 2.21488
R2545 VSS.n9465 VSS.n9466 4.5005
R2546 VSS.n9468 VSS.n9467 0.0732424
R2547 VSS.n9466 VSS.n9468 2.21488
R2548 VSS.n9471 VSS.n9470 0.0732424
R2549 VSS.n9466 VSS.n9471 2.21488
R2550 VSS.n9480 VSS.n9481 4.5005
R2551 VSS.n9482 VSS.n9483 0.0732424
R2552 VSS.n9483 VSS.n9481 2.21488
R2553 VSS.n9485 VSS.n9486 0.0732424
R2554 VSS.n9486 VSS.n9481 2.21488
R2555 VSS.n9495 VSS.n9496 4.5005
R2556 VSS.n9498 VSS.n9497 0.0732424
R2557 VSS.n9496 VSS.n9498 2.21488
R2558 VSS.n9501 VSS.n9500 0.0732424
R2559 VSS.n9496 VSS.n9501 2.21488
R2560 VSS.n9510 VSS.n9511 4.5005
R2561 VSS.n9513 VSS.n9512 0.0732424
R2562 VSS.n9511 VSS.n9513 2.21488
R2563 VSS.n9516 VSS.n9515 0.0732424
R2564 VSS.n9511 VSS.n9516 2.21488
R2565 VSS.n9525 VSS.n9526 4.5005
R2566 VSS.n9528 VSS.n9527 0.0732424
R2567 VSS.n9526 VSS.n9528 2.21488
R2568 VSS.n9531 VSS.n9530 0.0732424
R2569 VSS.n9526 VSS.n9531 2.21488
R2570 VSS.n9540 VSS.n9541 4.5005
R2571 VSS.n9543 VSS.n9542 0.0732424
R2572 VSS.n9541 VSS.n9543 2.21488
R2573 VSS.n9546 VSS.n9545 0.0732424
R2574 VSS.n9541 VSS.n9546 2.21488
R2575 VSS.n9555 VSS.n9556 4.5005
R2576 VSS.n9558 VSS.n9557 0.0732424
R2577 VSS.n9556 VSS.n9558 2.21488
R2578 VSS.n9561 VSS.n9560 0.0732424
R2579 VSS.n9556 VSS.n9561 2.21488
R2580 VSS.n9541 VSS.n9556 0.0584021
R2581 VSS.n7184 VSS.n9541 0.0596608
R2582 VSS.n7184 VSS.n9526 0.0244161
R2583 VSS.n9526 VSS.n9511 0.0585594
R2584 VSS.n9511 VSS.n9496 0.0584021
R2585 VSS.n9481 VSS.n9496 0.0596608
R2586 VSS.n9481 VSS.n9466 0.0244161
R2587 VSS.n9466 VSS.n9451 0.0585594
R2588 VSS.n9451 VSS.n9436 0.0584021
R2589 VSS.n9436 VSS 0.16272
R2590 VSS VSS.n9421 0.143052
R2591 VSS.n9406 VSS.n9421 0.0584021
R2592 VSS.n9391 VSS.n9406 0.0584021
R2593 VSS.n9376 VSS.n9391 0.0244161
R2594 VSS.n9376 VSS.n9361 0.0598182
R2595 VSS.n9361 VSS.n9346 0.0584021
R2596 VSS.n9331 VSS.n9346 0.0584021
R2597 VSS.n9316 VSS.n9331 0.0244161
R2598 VSS.n9316 VSS.n9301 0.0598182
R2599 VSS.n9301 VSS.n9286 0.0584021
R2600 VSS.n9286 VSS.n9271 0.0231573
R2601 VSS.n9256 VSS.n9271 0.0584021
R2602 VSS.n9241 VSS.n9256 0.0596608
R2603 VSS.n9241 VSS.n9226 0.0244161
R2604 VSS.n9226 VSS.n9211 0.0585594
R2605 VSS.n9211 VSS.n9196 0.0584021
R2606 VSS.n9181 VSS.n9196 0.0596608
R2607 VSS.n9181 VSS.n9166 0.0244161
R2608 VSS.n9166 VSS.n9151 0.0585594
R2609 VSS.n9151 VSS.n9136 0.0584021
R2610 VSS.n9136 VSS 0.16272
R2611 VSS VSS.n9121 0.143052
R2612 VSS.n9106 VSS.n9121 0.0584021
R2613 VSS.n9091 VSS.n9106 0.0584021
R2614 VSS.n9076 VSS.n9091 0.0244161
R2615 VSS.n9076 VSS.n9061 0.0598182
R2616 VSS.n9061 VSS.n9046 0.0584021
R2617 VSS.n9031 VSS.n9046 0.0584021
R2618 VSS.n9016 VSS.n9031 0.0244161
R2619 VSS.n9016 VSS.n9001 0.0598182
R2620 VSS.n9001 VSS.n8986 0.0584021
R2621 VSS.n8986 VSS.n8971 0.0231573
R2622 VSS.n8956 VSS.n8971 0.0584021
R2623 VSS.n8941 VSS.n8956 0.0596608
R2624 VSS.n8941 VSS.n8926 0.0244161
R2625 VSS.n8926 VSS.n8911 0.0585594
R2626 VSS.n8911 VSS.n8896 0.0584021
R2627 VSS.n8881 VSS.n8896 0.0596608
R2628 VSS.n8881 VSS.n8866 0.0244161
R2629 VSS.n8866 VSS.n8851 0.0585594
R2630 VSS.n8851 VSS.n8836 0.0584021
R2631 VSS.n8836 VSS 0.16272
R2632 VSS VSS.n8821 0.143052
R2633 VSS.n8806 VSS.n8821 0.0584021
R2634 VSS.n8791 VSS.n8806 0.0584021
R2635 VSS.n8776 VSS.n8791 0.0244161
R2636 VSS.n8776 VSS.n8761 0.0598182
R2637 VSS.n8761 VSS.n8746 0.0584021
R2638 VSS.n8731 VSS.n8746 0.0584021
R2639 VSS.n8716 VSS.n8731 0.0244161
R2640 VSS.n8716 VSS.n8701 0.0598182
R2641 VSS.n8701 VSS.n8686 0.0584021
R2642 VSS.n8686 VSS.n8671 0.0231573
R2643 VSS.n8656 VSS.n8671 0.0584021
R2644 VSS.n8641 VSS.n8656 0.0596608
R2645 VSS.n8641 VSS.n8626 0.0244161
R2646 VSS.n8626 VSS.n8611 0.0585594
R2647 VSS.n8611 VSS.n8596 0.0584021
R2648 VSS.n8581 VSS.n8596 0.0596608
R2649 VSS.n8581 VSS.n8566 0.0244161
R2650 VSS.n8566 VSS.n8551 0.0585594
R2651 VSS.n8551 VSS.n8536 0.0584021
R2652 VSS.n8536 VSS 0.16272
R2653 VSS VSS.n8521 0.143052
R2654 VSS.n8506 VSS.n8521 0.0584021
R2655 VSS.n8491 VSS.n8506 0.0584021
R2656 VSS.n8476 VSS.n8491 0.0244161
R2657 VSS.n8476 VSS.n8461 0.0598182
R2658 VSS.n8461 VSS.n8446 0.0584021
R2659 VSS.n8431 VSS.n8446 0.0584021
R2660 VSS.n8416 VSS.n8431 0.0244161
R2661 VSS.n8416 VSS.n8401 0.0598182
R2662 VSS.n8401 VSS.n8386 0.0584021
R2663 VSS.n8386 VSS.n8371 0.0231573
R2664 VSS.n8356 VSS.n8371 0.0584021
R2665 VSS.n8341 VSS.n8356 0.0596608
R2666 VSS.n8341 VSS.n8326 0.0244161
R2667 VSS.n8326 VSS.n8311 0.0585594
R2668 VSS.n8311 VSS.n8296 0.0584021
R2669 VSS.n8281 VSS.n8296 0.0596608
R2670 VSS.n8281 VSS.n8266 0.0244161
R2671 VSS.n8266 VSS.n8251 0.0585594
R2672 VSS.n8251 VSS.n8236 0.0584021
R2673 VSS.n8236 VSS 0.16272
R2674 VSS VSS.n8221 0.143052
R2675 VSS.n8206 VSS.n8221 0.0584021
R2676 VSS.n8191 VSS.n8206 0.0584021
R2677 VSS.n8176 VSS.n8191 0.0244161
R2678 VSS.n8176 VSS.n8161 0.0598182
R2679 VSS.n8161 VSS.n8146 0.0584021
R2680 VSS.n8131 VSS.n8146 0.0584021
R2681 VSS.n8116 VSS.n8131 0.0244161
R2682 VSS.n8116 VSS.n8101 0.0598182
R2683 VSS.n8101 VSS.n8086 0.0584021
R2684 VSS.n8086 VSS.n8071 0.0231573
R2685 VSS.n8056 VSS.n8071 0.0584021
R2686 VSS.n8041 VSS.n8056 0.0596608
R2687 VSS.n8041 VSS.n8026 0.0244161
R2688 VSS.n8026 VSS.n8011 0.0585594
R2689 VSS.n8011 VSS.n7996 0.0584021
R2690 VSS.n7981 VSS.n7996 0.0596608
R2691 VSS.n7981 VSS.n7966 0.0244161
R2692 VSS.n7966 VSS.n7951 0.0585594
R2693 VSS.n7951 VSS.n7936 0.0584021
R2694 VSS.n7936 VSS 0.16272
R2695 VSS VSS.n7921 0.143052
R2696 VSS.n7906 VSS.n7921 0.0584021
R2697 VSS.n7891 VSS.n7906 0.0584021
R2698 VSS.n7876 VSS.n7891 0.0244161
R2699 VSS.n7876 VSS.n7861 0.0598182
R2700 VSS.n7861 VSS.n7846 0.0584021
R2701 VSS.n7831 VSS.n7846 0.0584021
R2702 VSS.n7816 VSS.n7831 0.0244161
R2703 VSS.n7816 VSS.n7801 0.0598182
R2704 VSS.n7801 VSS.n7786 0.0584021
R2705 VSS.n7786 VSS.n7771 0.0231573
R2706 VSS.n7756 VSS.n7771 0.0584021
R2707 VSS.n7741 VSS.n7756 0.0596608
R2708 VSS.n7741 VSS.n7726 0.0244161
R2709 VSS.n7726 VSS.n7711 0.0585594
R2710 VSS.n7711 VSS.n7696 0.0584021
R2711 VSS.n7681 VSS.n7696 0.0596608
R2712 VSS.n7681 VSS.n7666 0.0244161
R2713 VSS.n7666 VSS.n7651 0.0585594
R2714 VSS.n7651 VSS.n7636 0.0584021
R2715 VSS.n7636 VSS 0.16272
R2716 VSS VSS.n7621 0.143052
R2717 VSS.n7606 VSS.n7621 0.0584021
R2718 VSS.n7591 VSS.n7606 0.0584021
R2719 VSS.n7576 VSS.n7591 0.0244161
R2720 VSS.n7576 VSS.n7561 0.0598182
R2721 VSS.n7561 VSS.n7546 0.0584021
R2722 VSS.n7531 VSS.n7546 0.0584021
R2723 VSS.n7516 VSS.n7531 0.0244161
R2724 VSS.n7516 VSS.n7501 0.0598182
R2725 VSS.n7501 VSS.n7486 0.0584021
R2726 VSS.n7486 VSS.n7471 0.0231573
R2727 VSS.n7456 VSS.n7471 0.0584021
R2728 VSS.n7441 VSS.n7456 0.0596608
R2729 VSS.n7441 VSS.n7426 0.0244161
R2730 VSS.n7426 VSS.n7411 0.0585594
R2731 VSS.n7411 VSS.n7396 0.0584021
R2732 VSS.n7381 VSS.n7396 0.0596608
R2733 VSS.n7381 VSS.n7366 0.0244161
R2734 VSS.n7366 VSS.n7351 0.0585594
R2735 VSS.n7351 VSS.n7336 0.0584021
R2736 VSS.n7336 VSS 0.16272
R2737 VSS VSS.n7321 0.143052
R2738 VSS.n7306 VSS.n7321 0.0584021
R2739 VSS.n7291 VSS.n7306 0.0584021
R2740 VSS.n7276 VSS.n7291 0.0244161
R2741 VSS.n7276 VSS.n7261 0.0598182
R2742 VSS.n7261 VSS.n7246 0.0584021
R2743 VSS.n7231 VSS.n7246 0.0584021
R2744 VSS.n7216 VSS.n7231 0.0244161
R2745 VSS.n7216 VSS.n7201 0.0598182
R2746 VSS.n7201 VSS.n7186 0.0584021
R2747 VSS.n9557 VSS.n9562 4.5005
R2748 VSS.n9559 VSS.n9563 4.5005
R2749 VSS.n9560 VSS.n9564 4.5005
R2750 VSS.n9561 VSS.n9565 4.57324
R2751 VSS.n9557 VSS.n9555 0.147342
R2752 VSS.n9558 VSS.n9559 0.0732424
R2753 VSS.n9559 VSS.n9560 0.147342
R2754 VSS.n9562 VSS.n9566 0.0721009
R2755 VSS.n9567 VSS.n9563 4.5005
R2756 VSS.n9568 VSS.n9564 4.5005
R2757 VSS.n9569 VSS.n9565 4.5005
R2758 VSS.n9555 VSS.n9566 4.57442
R2759 VSS.n9562 VSS.n9563 0.147342
R2760 VSS.n9563 VSS.n9564 0.147342
R2761 VSS.n9564 VSS.n9565 0.147342
R2762 VSS.n9566 VSS.n9567 2.39784
R2763 VSS.n9567 VSS.n9568 0.147342
R2764 VSS.n9568 VSS.n9569 0.147342
R2765 VSS.n9569 VSS.t47 3.13212
R2766 VSS.n9542 VSS.n9547 4.5005
R2767 VSS.n9544 VSS.n9548 4.5005
R2768 VSS.n9545 VSS.n9549 4.5005
R2769 VSS.n9546 VSS.n9550 4.57324
R2770 VSS.n9542 VSS.n9540 0.147342
R2771 VSS.n9543 VSS.n9544 0.0732424
R2772 VSS.n9544 VSS.n9545 0.147342
R2773 VSS.n9547 VSS.n9551 0.0721009
R2774 VSS.n9552 VSS.n9548 4.5005
R2775 VSS.n9553 VSS.n9549 4.5005
R2776 VSS.n9554 VSS.n9550 4.5005
R2777 VSS.n9540 VSS.n9551 4.57442
R2778 VSS.n9547 VSS.n9548 0.147342
R2779 VSS.n9548 VSS.n9549 0.147342
R2780 VSS.n9549 VSS.n9550 0.147342
R2781 VSS.n9551 VSS.n9552 2.39784
R2782 VSS.n9552 VSS.n9553 0.147342
R2783 VSS.n9553 VSS.n9554 0.147342
R2784 VSS.n9554 VSS.t509 3.13212
R2785 VSS.n9527 VSS.n9532 4.5005
R2786 VSS.n9529 VSS.n9533 4.5005
R2787 VSS.n9530 VSS.n9534 4.5005
R2788 VSS.n9531 VSS.n9535 4.57324
R2789 VSS.n9527 VSS.n9525 0.147342
R2790 VSS.n9528 VSS.n9529 0.0732424
R2791 VSS.n9529 VSS.n9530 0.147342
R2792 VSS.n9532 VSS.n9536 0.0721009
R2793 VSS.n9537 VSS.n9533 4.5005
R2794 VSS.n9538 VSS.n9534 4.5005
R2795 VSS.n9539 VSS.n9535 4.5005
R2796 VSS.n9525 VSS.n9536 4.57442
R2797 VSS.n9532 VSS.n9533 0.147342
R2798 VSS.n9533 VSS.n9534 0.147342
R2799 VSS.n9534 VSS.n9535 0.147342
R2800 VSS.n9536 VSS.n9537 2.39784
R2801 VSS.n9537 VSS.n9538 0.147342
R2802 VSS.n9538 VSS.n9539 0.147342
R2803 VSS.n9539 VSS.t56 3.13212
R2804 VSS.n9512 VSS.n9517 4.5005
R2805 VSS.n9514 VSS.n9518 4.5005
R2806 VSS.n9515 VSS.n9519 4.5005
R2807 VSS.n9516 VSS.n9520 4.57324
R2808 VSS.n9512 VSS.n9510 0.147342
R2809 VSS.n9513 VSS.n9514 0.0732424
R2810 VSS.n9514 VSS.n9515 0.147342
R2811 VSS.n9517 VSS.n9521 0.0721009
R2812 VSS.n9522 VSS.n9518 4.5005
R2813 VSS.n9523 VSS.n9519 4.5005
R2814 VSS.n9524 VSS.n9520 4.5005
R2815 VSS.n9510 VSS.n9521 4.57442
R2816 VSS.n9517 VSS.n9518 0.147342
R2817 VSS.n9518 VSS.n9519 0.147342
R2818 VSS.n9519 VSS.n9520 0.147342
R2819 VSS.n9521 VSS.n9522 2.39784
R2820 VSS.n9522 VSS.n9523 0.147342
R2821 VSS.n9523 VSS.n9524 0.147342
R2822 VSS.n9524 VSS.t205 3.13212
R2823 VSS.n9497 VSS.n9502 4.5005
R2824 VSS.n9499 VSS.n9503 4.5005
R2825 VSS.n9500 VSS.n9504 4.5005
R2826 VSS.n9501 VSS.n9505 4.57324
R2827 VSS.n9497 VSS.n9495 0.147342
R2828 VSS.n9498 VSS.n9499 0.0732424
R2829 VSS.n9499 VSS.n9500 0.147342
R2830 VSS.n9502 VSS.n9506 0.0721009
R2831 VSS.n9507 VSS.n9503 4.5005
R2832 VSS.n9508 VSS.n9504 4.5005
R2833 VSS.n9509 VSS.n9505 4.5005
R2834 VSS.n9495 VSS.n9506 4.57442
R2835 VSS.n9502 VSS.n9503 0.147342
R2836 VSS.n9503 VSS.n9504 0.147342
R2837 VSS.n9504 VSS.n9505 0.147342
R2838 VSS.n9506 VSS.n9507 2.39784
R2839 VSS.n9507 VSS.n9508 0.147342
R2840 VSS.n9508 VSS.n9509 0.147342
R2841 VSS.n9509 VSS.t423 3.13212
R2842 VSS.n9487 VSS.n9482 4.5005
R2843 VSS.n9488 VSS.n9484 4.5005
R2844 VSS.n9489 VSS.n9485 4.5005
R2845 VSS.n9490 VSS.n9486 4.57324
R2846 VSS.n9480 VSS.n9482 0.147342
R2847 VSS.n9483 VSS.n9484 0.0732424
R2848 VSS.n9484 VSS.n9485 0.147342
R2849 VSS.n9491 VSS.n9487 0.0722544
R2850 VSS.n9492 VSS.n9488 4.5005
R2851 VSS.n9493 VSS.n9489 4.5005
R2852 VSS.n9494 VSS.n9490 4.5005
R2853 VSS.n9491 VSS.n9480 4.57426
R2854 VSS.n9487 VSS.n9488 0.147342
R2855 VSS.n9488 VSS.n9489 0.147342
R2856 VSS.n9489 VSS.n9490 0.147342
R2857 VSS.n9492 VSS.n9491 2.37296
R2858 VSS.n9493 VSS.n9492 0.127318
R2859 VSS.n9494 VSS.n9493 0.127318
R2860 VSS.t41 VSS.n9494 2.73618
R2861 VSS.n9467 VSS.n9472 4.5005
R2862 VSS.n9469 VSS.n9473 4.5005
R2863 VSS.n9470 VSS.n9474 4.5005
R2864 VSS.n9471 VSS.n9475 4.57324
R2865 VSS.n9467 VSS.n9465 0.147342
R2866 VSS.n9468 VSS.n9469 0.0732424
R2867 VSS.n9469 VSS.n9470 0.147342
R2868 VSS.n9472 VSS.n9476 0.0721009
R2869 VSS.n9477 VSS.n9473 4.5005
R2870 VSS.n9478 VSS.n9474 4.5005
R2871 VSS.n9479 VSS.n9475 4.5005
R2872 VSS.n9465 VSS.n9476 4.57442
R2873 VSS.n9472 VSS.n9473 0.147342
R2874 VSS.n9473 VSS.n9474 0.147342
R2875 VSS.n9474 VSS.n9475 0.147342
R2876 VSS.n9476 VSS.n9477 2.39784
R2877 VSS.n9477 VSS.n9478 0.147342
R2878 VSS.n9478 VSS.n9479 0.147342
R2879 VSS.n9479 VSS.t552 3.13212
R2880 VSS.n9452 VSS.n9457 4.5005
R2881 VSS.n9454 VSS.n9458 4.5005
R2882 VSS.n9455 VSS.n9459 4.5005
R2883 VSS.n9456 VSS.n9460 4.57324
R2884 VSS.n9452 VSS.n9450 0.147342
R2885 VSS.n9453 VSS.n9454 0.0732424
R2886 VSS.n9454 VSS.n9455 0.147342
R2887 VSS.n9457 VSS.n9461 0.0721009
R2888 VSS.n9462 VSS.n9458 4.5005
R2889 VSS.n9463 VSS.n9459 4.5005
R2890 VSS.n9464 VSS.n9460 4.5005
R2891 VSS.n9450 VSS.n9461 4.57442
R2892 VSS.n9457 VSS.n9458 0.147342
R2893 VSS.n9458 VSS.n9459 0.147342
R2894 VSS.n9459 VSS.n9460 0.147342
R2895 VSS.n9461 VSS.n9462 2.39784
R2896 VSS.n9462 VSS.n9463 0.147342
R2897 VSS.n9463 VSS.n9464 0.147342
R2898 VSS.n9464 VSS.t454 3.13212
R2899 VSS.n9437 VSS.n9442 4.5005
R2900 VSS.n9439 VSS.n9443 4.5005
R2901 VSS.n9440 VSS.n9444 4.5005
R2902 VSS.n9441 VSS.n9445 4.57324
R2903 VSS.n9437 VSS.n9435 0.147342
R2904 VSS.n9438 VSS.n9439 0.0732424
R2905 VSS.n9439 VSS.n9440 0.147342
R2906 VSS.n9442 VSS.n9446 0.0721009
R2907 VSS.n9447 VSS.n9443 4.5005
R2908 VSS.n9448 VSS.n9444 4.5005
R2909 VSS.n9449 VSS.n9445 4.5005
R2910 VSS.n9435 VSS.n9446 4.57442
R2911 VSS.n9442 VSS.n9443 0.147342
R2912 VSS.n9443 VSS.n9444 0.147342
R2913 VSS.n9444 VSS.n9445 0.147342
R2914 VSS.n9446 VSS.n9447 2.39784
R2915 VSS.n9447 VSS.n9448 0.147342
R2916 VSS.n9448 VSS.n9449 0.147342
R2917 VSS.n9449 VSS.t588 3.13212
R2918 VSS.n9422 VSS.n9427 4.5005
R2919 VSS.n9424 VSS.n9428 4.5005
R2920 VSS.n9425 VSS.n9429 4.5005
R2921 VSS.n9426 VSS.n9430 4.57324
R2922 VSS.n9422 VSS.n9420 0.147342
R2923 VSS.n9423 VSS.n9424 0.0732424
R2924 VSS.n9424 VSS.n9425 0.147342
R2925 VSS.n9427 VSS.n9431 0.0721009
R2926 VSS.n9432 VSS.n9428 4.5005
R2927 VSS.n9433 VSS.n9429 4.5005
R2928 VSS.n9434 VSS.n9430 4.5005
R2929 VSS.n9420 VSS.n9431 4.57442
R2930 VSS.n9427 VSS.n9428 0.147342
R2931 VSS.n9428 VSS.n9429 0.147342
R2932 VSS.n9429 VSS.n9430 0.147342
R2933 VSS.n9431 VSS.n9432 2.39784
R2934 VSS.n9432 VSS.n9433 0.147342
R2935 VSS.n9433 VSS.n9434 0.147342
R2936 VSS.n9434 VSS.t486 3.13212
R2937 VSS.n9407 VSS.n9412 4.5005
R2938 VSS.n9409 VSS.n9413 4.5005
R2939 VSS.n9410 VSS.n9414 4.5005
R2940 VSS.n9411 VSS.n9415 4.57324
R2941 VSS.n9407 VSS.n9405 0.147342
R2942 VSS.n9408 VSS.n9409 0.0732424
R2943 VSS.n9409 VSS.n9410 0.147342
R2944 VSS.n9412 VSS.n9416 0.0721009
R2945 VSS.n9417 VSS.n9413 4.5005
R2946 VSS.n9418 VSS.n9414 4.5005
R2947 VSS.n9419 VSS.n9415 4.5005
R2948 VSS.n9405 VSS.n9416 4.57442
R2949 VSS.n9412 VSS.n9413 0.147342
R2950 VSS.n9413 VSS.n9414 0.147342
R2951 VSS.n9414 VSS.n9415 0.147342
R2952 VSS.n9416 VSS.n9417 2.39784
R2953 VSS.n9417 VSS.n9418 0.147342
R2954 VSS.n9418 VSS.n9419 0.147342
R2955 VSS.n9419 VSS.t114 3.13212
R2956 VSS.n9392 VSS.n9397 4.5005
R2957 VSS.n9394 VSS.n9398 4.5005
R2958 VSS.n9395 VSS.n9399 4.5005
R2959 VSS.n9396 VSS.n9400 4.57324
R2960 VSS.n9392 VSS.n9390 0.147342
R2961 VSS.n9393 VSS.n9394 0.0732424
R2962 VSS.n9394 VSS.n9395 0.147342
R2963 VSS.n9397 VSS.n9401 0.0721009
R2964 VSS.n9402 VSS.n9398 4.5005
R2965 VSS.n9403 VSS.n9399 4.5005
R2966 VSS.n9404 VSS.n9400 4.5005
R2967 VSS.n9390 VSS.n9401 4.57442
R2968 VSS.n9397 VSS.n9398 0.147342
R2969 VSS.n9398 VSS.n9399 0.147342
R2970 VSS.n9399 VSS.n9400 0.147342
R2971 VSS.n9401 VSS.n9402 2.39784
R2972 VSS.n9402 VSS.n9403 0.147342
R2973 VSS.n9403 VSS.n9404 0.147342
R2974 VSS.n9404 VSS.t445 3.13212
R2975 VSS.n9382 VSS.n9377 4.5005
R2976 VSS.n9383 VSS.n9379 4.5005
R2977 VSS.n9384 VSS.n9380 4.5005
R2978 VSS.n9385 VSS.n9381 4.57324
R2979 VSS.n9375 VSS.n9377 0.147342
R2980 VSS.n9378 VSS.n9379 0.0732424
R2981 VSS.n9379 VSS.n9380 0.147342
R2982 VSS.n9386 VSS.n9382 0.0722544
R2983 VSS.n9387 VSS.n9383 4.5005
R2984 VSS.n9388 VSS.n9384 4.5005
R2985 VSS.n9389 VSS.n9385 4.5005
R2986 VSS.n9386 VSS.n9375 4.57426
R2987 VSS.n9382 VSS.n9383 0.147342
R2988 VSS.n9383 VSS.n9384 0.147342
R2989 VSS.n9384 VSS.n9385 0.147342
R2990 VSS.n9387 VSS.n9386 2.37296
R2991 VSS.n9388 VSS.n9387 0.127318
R2992 VSS.n9389 VSS.n9388 0.127318
R2993 VSS.t41 VSS.n9389 2.73618
R2994 VSS.n9362 VSS.n9367 4.5005
R2995 VSS.n9364 VSS.n9368 4.5005
R2996 VSS.n9365 VSS.n9369 4.5005
R2997 VSS.n9366 VSS.n9370 4.57324
R2998 VSS.n9362 VSS.n9360 0.147342
R2999 VSS.n9363 VSS.n9364 0.0732424
R3000 VSS.n9364 VSS.n9365 0.147342
R3001 VSS.n9367 VSS.n9371 0.0721009
R3002 VSS.n9372 VSS.n9368 4.5005
R3003 VSS.n9373 VSS.n9369 4.5005
R3004 VSS.n9374 VSS.n9370 4.5005
R3005 VSS.n9360 VSS.n9371 4.57442
R3006 VSS.n9367 VSS.n9368 0.147342
R3007 VSS.n9368 VSS.n9369 0.147342
R3008 VSS.n9369 VSS.n9370 0.147342
R3009 VSS.n9371 VSS.n9372 2.39784
R3010 VSS.n9372 VSS.n9373 0.147342
R3011 VSS.n9373 VSS.n9374 0.147342
R3012 VSS.n9374 VSS.t617 3.13212
R3013 VSS.n9347 VSS.n9352 4.5005
R3014 VSS.n9349 VSS.n9353 4.5005
R3015 VSS.n9350 VSS.n9354 4.5005
R3016 VSS.n9351 VSS.n9355 4.57324
R3017 VSS.n9347 VSS.n9345 0.147342
R3018 VSS.n9348 VSS.n9349 0.0732424
R3019 VSS.n9349 VSS.n9350 0.147342
R3020 VSS.n9352 VSS.n9356 0.0721009
R3021 VSS.n9357 VSS.n9353 4.5005
R3022 VSS.n9358 VSS.n9354 4.5005
R3023 VSS.n9359 VSS.n9355 4.5005
R3024 VSS.n9345 VSS.n9356 4.57442
R3025 VSS.n9352 VSS.n9353 0.147342
R3026 VSS.n9353 VSS.n9354 0.147342
R3027 VSS.n9354 VSS.n9355 0.147342
R3028 VSS.n9356 VSS.n9357 2.39784
R3029 VSS.n9357 VSS.n9358 0.147342
R3030 VSS.n9358 VSS.n9359 0.147342
R3031 VSS.n9359 VSS.t521 3.13212
R3032 VSS.n9332 VSS.n9337 4.5005
R3033 VSS.n9334 VSS.n9338 4.5005
R3034 VSS.n9335 VSS.n9339 4.5005
R3035 VSS.n9336 VSS.n9340 4.57324
R3036 VSS.n9332 VSS.n9330 0.147342
R3037 VSS.n9333 VSS.n9334 0.0732424
R3038 VSS.n9334 VSS.n9335 0.147342
R3039 VSS.n9337 VSS.n9341 0.0721009
R3040 VSS.n9342 VSS.n9338 4.5005
R3041 VSS.n9343 VSS.n9339 4.5005
R3042 VSS.n9344 VSS.n9340 4.5005
R3043 VSS.n9330 VSS.n9341 4.57442
R3044 VSS.n9337 VSS.n9338 0.147342
R3045 VSS.n9338 VSS.n9339 0.147342
R3046 VSS.n9339 VSS.n9340 0.147342
R3047 VSS.n9341 VSS.n9342 2.39784
R3048 VSS.n9342 VSS.n9343 0.147342
R3049 VSS.n9343 VSS.n9344 0.147342
R3050 VSS.n9344 VSS.t526 3.13212
R3051 VSS.n9322 VSS.n9317 4.5005
R3052 VSS.n9323 VSS.n9319 4.5005
R3053 VSS.n9324 VSS.n9320 4.5005
R3054 VSS.n9325 VSS.n9321 4.57324
R3055 VSS.n9315 VSS.n9317 0.147342
R3056 VSS.n9318 VSS.n9319 0.0732424
R3057 VSS.n9319 VSS.n9320 0.147342
R3058 VSS.n9326 VSS.n9322 0.0722544
R3059 VSS.n9327 VSS.n9323 4.5005
R3060 VSS.n9328 VSS.n9324 4.5005
R3061 VSS.n9329 VSS.n9325 4.5005
R3062 VSS.n9326 VSS.n9315 4.57426
R3063 VSS.n9322 VSS.n9323 0.147342
R3064 VSS.n9323 VSS.n9324 0.147342
R3065 VSS.n9324 VSS.n9325 0.147342
R3066 VSS.n9327 VSS.n9326 2.37296
R3067 VSS.n9328 VSS.n9327 0.127318
R3068 VSS.n9329 VSS.n9328 0.127318
R3069 VSS.t41 VSS.n9329 2.73618
R3070 VSS.n9302 VSS.n9307 4.5005
R3071 VSS.n9304 VSS.n9308 4.5005
R3072 VSS.n9305 VSS.n9309 4.5005
R3073 VSS.n9306 VSS.n9310 4.57324
R3074 VSS.n9302 VSS.n9300 0.147342
R3075 VSS.n9303 VSS.n9304 0.0732424
R3076 VSS.n9304 VSS.n9305 0.147342
R3077 VSS.n9307 VSS.n9311 0.0721009
R3078 VSS.n9312 VSS.n9308 4.5005
R3079 VSS.n9313 VSS.n9309 4.5005
R3080 VSS.n9314 VSS.n9310 4.5005
R3081 VSS.n9300 VSS.n9311 4.57442
R3082 VSS.n9307 VSS.n9308 0.147342
R3083 VSS.n9308 VSS.n9309 0.147342
R3084 VSS.n9309 VSS.n9310 0.147342
R3085 VSS.n9311 VSS.n9312 2.39784
R3086 VSS.n9312 VSS.n9313 0.147342
R3087 VSS.n9313 VSS.n9314 0.147342
R3088 VSS.n9314 VSS.t151 3.13212
R3089 VSS.n9287 VSS.n9292 4.5005
R3090 VSS.n9289 VSS.n9293 4.5005
R3091 VSS.n9290 VSS.n9294 4.5005
R3092 VSS.n9291 VSS.n9295 4.57324
R3093 VSS.n9287 VSS.n9285 0.147342
R3094 VSS.n9288 VSS.n9289 0.0732424
R3095 VSS.n9289 VSS.n9290 0.147342
R3096 VSS.n9292 VSS.n9296 0.0721009
R3097 VSS.n9297 VSS.n9293 4.5005
R3098 VSS.n9298 VSS.n9294 4.5005
R3099 VSS.n9299 VSS.n9295 4.5005
R3100 VSS.n9285 VSS.n9296 4.57442
R3101 VSS.n9292 VSS.n9293 0.147342
R3102 VSS.n9293 VSS.n9294 0.147342
R3103 VSS.n9294 VSS.n9295 0.147342
R3104 VSS.n9296 VSS.n9297 2.39784
R3105 VSS.n9297 VSS.n9298 0.147342
R3106 VSS.n9298 VSS.n9299 0.147342
R3107 VSS.n9299 VSS.t475 3.13212
R3108 VSS.n9272 VSS.n9277 4.5005
R3109 VSS.n9274 VSS.n9278 4.5005
R3110 VSS.n9275 VSS.n9279 4.5005
R3111 VSS.n9276 VSS.n9280 4.57324
R3112 VSS.n9272 VSS.n9270 0.147342
R3113 VSS.n9273 VSS.n9274 0.0732424
R3114 VSS.n9274 VSS.n9275 0.147342
R3115 VSS.n9277 VSS.n9281 0.0721009
R3116 VSS.n9282 VSS.n9278 4.5005
R3117 VSS.n9283 VSS.n9279 4.5005
R3118 VSS.n9284 VSS.n9280 4.5005
R3119 VSS.n9270 VSS.n9281 4.57442
R3120 VSS.n9277 VSS.n9278 0.147342
R3121 VSS.n9278 VSS.n9279 0.147342
R3122 VSS.n9279 VSS.n9280 0.147342
R3123 VSS.n9281 VSS.n9282 2.39784
R3124 VSS.n9282 VSS.n9283 0.147342
R3125 VSS.n9283 VSS.n9284 0.147342
R3126 VSS.n9284 VSS.t46 3.13212
R3127 VSS.n9257 VSS.n9262 4.5005
R3128 VSS.n9259 VSS.n9263 4.5005
R3129 VSS.n9260 VSS.n9264 4.5005
R3130 VSS.n9261 VSS.n9265 4.57324
R3131 VSS.n9257 VSS.n9255 0.147342
R3132 VSS.n9258 VSS.n9259 0.0732424
R3133 VSS.n9259 VSS.n9260 0.147342
R3134 VSS.n9262 VSS.n9266 0.0721009
R3135 VSS.n9267 VSS.n9263 4.5005
R3136 VSS.n9268 VSS.n9264 4.5005
R3137 VSS.n9269 VSS.n9265 4.5005
R3138 VSS.n9255 VSS.n9266 4.57442
R3139 VSS.n9262 VSS.n9263 0.147342
R3140 VSS.n9263 VSS.n9264 0.147342
R3141 VSS.n9264 VSS.n9265 0.147342
R3142 VSS.n9266 VSS.n9267 2.39784
R3143 VSS.n9267 VSS.n9268 0.147342
R3144 VSS.n9268 VSS.n9269 0.147342
R3145 VSS.n9269 VSS.t508 3.13212
R3146 VSS.n9247 VSS.n9242 4.5005
R3147 VSS.n9248 VSS.n9244 4.5005
R3148 VSS.n9249 VSS.n9245 4.5005
R3149 VSS.n9250 VSS.n9246 4.57324
R3150 VSS.n9240 VSS.n9242 0.147342
R3151 VSS.n9243 VSS.n9244 0.0732424
R3152 VSS.n9244 VSS.n9245 0.147342
R3153 VSS.n9251 VSS.n9247 0.0722544
R3154 VSS.n9252 VSS.n9248 4.5005
R3155 VSS.n9253 VSS.n9249 4.5005
R3156 VSS.n9254 VSS.n9250 4.5005
R3157 VSS.n9251 VSS.n9240 4.57426
R3158 VSS.n9247 VSS.n9248 0.147342
R3159 VSS.n9248 VSS.n9249 0.147342
R3160 VSS.n9249 VSS.n9250 0.147342
R3161 VSS.n9252 VSS.n9251 2.37296
R3162 VSS.n9253 VSS.n9252 0.127318
R3163 VSS.n9254 VSS.n9253 0.127318
R3164 VSS.t41 VSS.n9254 2.73618
R3165 VSS.n9227 VSS.n9232 4.5005
R3166 VSS.n9229 VSS.n9233 4.5005
R3167 VSS.n9230 VSS.n9234 4.5005
R3168 VSS.n9231 VSS.n9235 4.57324
R3169 VSS.n9227 VSS.n9225 0.147342
R3170 VSS.n9228 VSS.n9229 0.0732424
R3171 VSS.n9229 VSS.n9230 0.147342
R3172 VSS.n9232 VSS.n9236 0.0721009
R3173 VSS.n9237 VSS.n9233 4.5005
R3174 VSS.n9238 VSS.n9234 4.5005
R3175 VSS.n9239 VSS.n9235 4.5005
R3176 VSS.n9225 VSS.n9236 4.57442
R3177 VSS.n9232 VSS.n9233 0.147342
R3178 VSS.n9233 VSS.n9234 0.147342
R3179 VSS.n9234 VSS.n9235 0.147342
R3180 VSS.n9236 VSS.n9237 2.39784
R3181 VSS.n9237 VSS.n9238 0.147342
R3182 VSS.n9238 VSS.n9239 0.147342
R3183 VSS.n9239 VSS.t576 3.13212
R3184 VSS.n9212 VSS.n9217 4.5005
R3185 VSS.n9214 VSS.n9218 4.5005
R3186 VSS.n9215 VSS.n9219 4.5005
R3187 VSS.n9216 VSS.n9220 4.57324
R3188 VSS.n9212 VSS.n9210 0.147342
R3189 VSS.n9213 VSS.n9214 0.0732424
R3190 VSS.n9214 VSS.n9215 0.147342
R3191 VSS.n9217 VSS.n9221 0.0721009
R3192 VSS.n9222 VSS.n9218 4.5005
R3193 VSS.n9223 VSS.n9219 4.5005
R3194 VSS.n9224 VSS.n9220 4.5005
R3195 VSS.n9210 VSS.n9221 4.57442
R3196 VSS.n9217 VSS.n9218 0.147342
R3197 VSS.n9218 VSS.n9219 0.147342
R3198 VSS.n9219 VSS.n9220 0.147342
R3199 VSS.n9221 VSS.n9222 2.39784
R3200 VSS.n9222 VSS.n9223 0.147342
R3201 VSS.n9223 VSS.n9224 0.147342
R3202 VSS.n9224 VSS.t201 3.13212
R3203 VSS.n9197 VSS.n9202 4.5005
R3204 VSS.n9199 VSS.n9203 4.5005
R3205 VSS.n9200 VSS.n9204 4.5005
R3206 VSS.n9201 VSS.n9205 4.57324
R3207 VSS.n9197 VSS.n9195 0.147342
R3208 VSS.n9198 VSS.n9199 0.0732424
R3209 VSS.n9199 VSS.n9200 0.147342
R3210 VSS.n9202 VSS.n9206 0.0721009
R3211 VSS.n9207 VSS.n9203 4.5005
R3212 VSS.n9208 VSS.n9204 4.5005
R3213 VSS.n9209 VSS.n9205 4.5005
R3214 VSS.n9195 VSS.n9206 4.57442
R3215 VSS.n9202 VSS.n9203 0.147342
R3216 VSS.n9203 VSS.n9204 0.147342
R3217 VSS.n9204 VSS.n9205 0.147342
R3218 VSS.n9206 VSS.n9207 2.39784
R3219 VSS.n9207 VSS.n9208 0.147342
R3220 VSS.n9208 VSS.n9209 0.147342
R3221 VSS.n9209 VSS.t389 3.13212
R3222 VSS.n9187 VSS.n9182 4.5005
R3223 VSS.n9188 VSS.n9184 4.5005
R3224 VSS.n9189 VSS.n9185 4.5005
R3225 VSS.n9190 VSS.n9186 4.57324
R3226 VSS.n9180 VSS.n9182 0.147342
R3227 VSS.n9183 VSS.n9184 0.0732424
R3228 VSS.n9184 VSS.n9185 0.147342
R3229 VSS.n9191 VSS.n9187 0.0722544
R3230 VSS.n9192 VSS.n9188 4.5005
R3231 VSS.n9193 VSS.n9189 4.5005
R3232 VSS.n9194 VSS.n9190 4.5005
R3233 VSS.n9191 VSS.n9180 4.57426
R3234 VSS.n9187 VSS.n9188 0.147342
R3235 VSS.n9188 VSS.n9189 0.147342
R3236 VSS.n9189 VSS.n9190 0.147342
R3237 VSS.n9192 VSS.n9191 2.37296
R3238 VSS.n9193 VSS.n9192 0.127318
R3239 VSS.n9194 VSS.n9193 0.127318
R3240 VSS.t41 VSS.n9194 2.73618
R3241 VSS.n9167 VSS.n9172 4.5005
R3242 VSS.n9169 VSS.n9173 4.5005
R3243 VSS.n9170 VSS.n9174 4.5005
R3244 VSS.n9171 VSS.n9175 4.57324
R3245 VSS.n9167 VSS.n9165 0.147342
R3246 VSS.n9168 VSS.n9169 0.0732424
R3247 VSS.n9169 VSS.n9170 0.147342
R3248 VSS.n9172 VSS.n9176 0.0721009
R3249 VSS.n9177 VSS.n9173 4.5005
R3250 VSS.n9178 VSS.n9174 4.5005
R3251 VSS.n9179 VSS.n9175 4.5005
R3252 VSS.n9165 VSS.n9176 4.57442
R3253 VSS.n9172 VSS.n9173 0.147342
R3254 VSS.n9173 VSS.n9174 0.147342
R3255 VSS.n9174 VSS.n9175 0.147342
R3256 VSS.n9176 VSS.n9177 2.39784
R3257 VSS.n9177 VSS.n9178 0.147342
R3258 VSS.n9178 VSS.n9179 0.147342
R3259 VSS.n9179 VSS.t541 3.13212
R3260 VSS.n9152 VSS.n9157 4.5005
R3261 VSS.n9154 VSS.n9158 4.5005
R3262 VSS.n9155 VSS.n9159 4.5005
R3263 VSS.n9156 VSS.n9160 4.57324
R3264 VSS.n9152 VSS.n9150 0.147342
R3265 VSS.n9153 VSS.n9154 0.0732424
R3266 VSS.n9154 VSS.n9155 0.147342
R3267 VSS.n9157 VSS.n9161 0.0721009
R3268 VSS.n9162 VSS.n9158 4.5005
R3269 VSS.n9163 VSS.n9159 4.5005
R3270 VSS.n9164 VSS.n9160 4.5005
R3271 VSS.n9150 VSS.n9161 4.57442
R3272 VSS.n9157 VSS.n9158 0.147342
R3273 VSS.n9158 VSS.n9159 0.147342
R3274 VSS.n9159 VSS.n9160 0.147342
R3275 VSS.n9161 VSS.n9162 2.39784
R3276 VSS.n9162 VSS.n9163 0.147342
R3277 VSS.n9163 VSS.n9164 0.147342
R3278 VSS.n9164 VSS.t452 3.13212
R3279 VSS.n9137 VSS.n9142 4.5005
R3280 VSS.n9139 VSS.n9143 4.5005
R3281 VSS.n9140 VSS.n9144 4.5005
R3282 VSS.n9141 VSS.n9145 4.57324
R3283 VSS.n9137 VSS.n9135 0.147342
R3284 VSS.n9138 VSS.n9139 0.0732424
R3285 VSS.n9139 VSS.n9140 0.147342
R3286 VSS.n9142 VSS.n9146 0.0721009
R3287 VSS.n9147 VSS.n9143 4.5005
R3288 VSS.n9148 VSS.n9144 4.5005
R3289 VSS.n9149 VSS.n9145 4.5005
R3290 VSS.n9135 VSS.n9146 4.57442
R3291 VSS.n9142 VSS.n9143 0.147342
R3292 VSS.n9143 VSS.n9144 0.147342
R3293 VSS.n9144 VSS.n9145 0.147342
R3294 VSS.n9146 VSS.n9147 2.39784
R3295 VSS.n9147 VSS.n9148 0.147342
R3296 VSS.n9148 VSS.n9149 0.147342
R3297 VSS.n9149 VSS.t586 3.13212
R3298 VSS.n9122 VSS.n9127 4.5005
R3299 VSS.n9124 VSS.n9128 4.5005
R3300 VSS.n9125 VSS.n9129 4.5005
R3301 VSS.n9126 VSS.n9130 4.57324
R3302 VSS.n9122 VSS.n9120 0.147342
R3303 VSS.n9123 VSS.n9124 0.0732424
R3304 VSS.n9124 VSS.n9125 0.147342
R3305 VSS.n9127 VSS.n9131 0.0721009
R3306 VSS.n9132 VSS.n9128 4.5005
R3307 VSS.n9133 VSS.n9129 4.5005
R3308 VSS.n9134 VSS.n9130 4.5005
R3309 VSS.n9120 VSS.n9131 4.57442
R3310 VSS.n9127 VSS.n9128 0.147342
R3311 VSS.n9128 VSS.n9129 0.147342
R3312 VSS.n9129 VSS.n9130 0.147342
R3313 VSS.n9131 VSS.n9132 2.39784
R3314 VSS.n9132 VSS.n9133 0.147342
R3315 VSS.n9133 VSS.n9134 0.147342
R3316 VSS.n9134 VSS.t66 3.13212
R3317 VSS.n9107 VSS.n9112 4.5005
R3318 VSS.n9109 VSS.n9113 4.5005
R3319 VSS.n9110 VSS.n9114 4.5005
R3320 VSS.n9111 VSS.n9115 4.57324
R3321 VSS.n9107 VSS.n9105 0.147342
R3322 VSS.n9108 VSS.n9109 0.0732424
R3323 VSS.n9109 VSS.n9110 0.147342
R3324 VSS.n9112 VSS.n9116 0.0721009
R3325 VSS.n9117 VSS.n9113 4.5005
R3326 VSS.n9118 VSS.n9114 4.5005
R3327 VSS.n9119 VSS.n9115 4.5005
R3328 VSS.n9105 VSS.n9116 4.57442
R3329 VSS.n9112 VSS.n9113 0.147342
R3330 VSS.n9113 VSS.n9114 0.147342
R3331 VSS.n9114 VSS.n9115 0.147342
R3332 VSS.n9116 VSS.n9117 2.39784
R3333 VSS.n9117 VSS.n9118 0.147342
R3334 VSS.n9118 VSS.n9119 0.147342
R3335 VSS.n9119 VSS.t116 3.13212
R3336 VSS.n9092 VSS.n9097 4.5005
R3337 VSS.n9094 VSS.n9098 4.5005
R3338 VSS.n9095 VSS.n9099 4.5005
R3339 VSS.n9096 VSS.n9100 4.57324
R3340 VSS.n9092 VSS.n9090 0.147342
R3341 VSS.n9093 VSS.n9094 0.0732424
R3342 VSS.n9094 VSS.n9095 0.147342
R3343 VSS.n9097 VSS.n9101 0.0721009
R3344 VSS.n9102 VSS.n9098 4.5005
R3345 VSS.n9103 VSS.n9099 4.5005
R3346 VSS.n9104 VSS.n9100 4.5005
R3347 VSS.n9090 VSS.n9101 4.57442
R3348 VSS.n9097 VSS.n9098 0.147342
R3349 VSS.n9098 VSS.n9099 0.147342
R3350 VSS.n9099 VSS.n9100 0.147342
R3351 VSS.n9101 VSS.n9102 2.39784
R3352 VSS.n9102 VSS.n9103 0.147342
R3353 VSS.n9103 VSS.n9104 0.147342
R3354 VSS.n9104 VSS.t477 3.13212
R3355 VSS.n9082 VSS.n9077 4.5005
R3356 VSS.n9083 VSS.n9079 4.5005
R3357 VSS.n9084 VSS.n9080 4.5005
R3358 VSS.n9085 VSS.n9081 4.57324
R3359 VSS.n9075 VSS.n9077 0.147342
R3360 VSS.n9078 VSS.n9079 0.0732424
R3361 VSS.n9079 VSS.n9080 0.147342
R3362 VSS.n9086 VSS.n9082 0.0722544
R3363 VSS.n9087 VSS.n9083 4.5005
R3364 VSS.n9088 VSS.n9084 4.5005
R3365 VSS.n9089 VSS.n9085 4.5005
R3366 VSS.n9086 VSS.n9075 4.57426
R3367 VSS.n9082 VSS.n9083 0.147342
R3368 VSS.n9083 VSS.n9084 0.147342
R3369 VSS.n9084 VSS.n9085 0.147342
R3370 VSS.n9087 VSS.n9086 2.37296
R3371 VSS.n9088 VSS.n9087 0.127318
R3372 VSS.n9089 VSS.n9088 0.127318
R3373 VSS.t41 VSS.n9089 2.73618
R3374 VSS.n9062 VSS.n9067 4.5005
R3375 VSS.n9064 VSS.n9068 4.5005
R3376 VSS.n9065 VSS.n9069 4.5005
R3377 VSS.n9066 VSS.n9070 4.57324
R3378 VSS.n9062 VSS.n9060 0.147342
R3379 VSS.n9063 VSS.n9064 0.0732424
R3380 VSS.n9064 VSS.n9065 0.147342
R3381 VSS.n9067 VSS.n9071 0.0721009
R3382 VSS.n9072 VSS.n9068 4.5005
R3383 VSS.n9073 VSS.n9069 4.5005
R3384 VSS.n9074 VSS.n9070 4.5005
R3385 VSS.n9060 VSS.n9071 4.57442
R3386 VSS.n9067 VSS.n9068 0.147342
R3387 VSS.n9068 VSS.n9069 0.147342
R3388 VSS.n9069 VSS.n9070 0.147342
R3389 VSS.n9071 VSS.n9072 2.39784
R3390 VSS.n9072 VSS.n9073 0.147342
R3391 VSS.n9073 VSS.n9074 0.147342
R3392 VSS.n9074 VSS.t573 3.13212
R3393 VSS.n9047 VSS.n9052 4.5005
R3394 VSS.n9049 VSS.n9053 4.5005
R3395 VSS.n9050 VSS.n9054 4.5005
R3396 VSS.n9051 VSS.n9055 4.57324
R3397 VSS.n9047 VSS.n9045 0.147342
R3398 VSS.n9048 VSS.n9049 0.0732424
R3399 VSS.n9049 VSS.n9050 0.147342
R3400 VSS.n9052 VSS.n9056 0.0721009
R3401 VSS.n9057 VSS.n9053 4.5005
R3402 VSS.n9058 VSS.n9054 4.5005
R3403 VSS.n9059 VSS.n9055 4.5005
R3404 VSS.n9045 VSS.n9056 4.57442
R3405 VSS.n9052 VSS.n9053 0.147342
R3406 VSS.n9053 VSS.n9054 0.147342
R3407 VSS.n9054 VSS.n9055 0.147342
R3408 VSS.n9056 VSS.n9057 2.39784
R3409 VSS.n9057 VSS.n9058 0.147342
R3410 VSS.n9058 VSS.n9059 0.147342
R3411 VSS.n9059 VSS.t51 3.13212
R3412 VSS.n9032 VSS.n9037 4.5005
R3413 VSS.n9034 VSS.n9038 4.5005
R3414 VSS.n9035 VSS.n9039 4.5005
R3415 VSS.n9036 VSS.n9040 4.57324
R3416 VSS.n9032 VSS.n9030 0.147342
R3417 VSS.n9033 VSS.n9034 0.0732424
R3418 VSS.n9034 VSS.n9035 0.147342
R3419 VSS.n9037 VSS.n9041 0.0721009
R3420 VSS.n9042 VSS.n9038 4.5005
R3421 VSS.n9043 VSS.n9039 4.5005
R3422 VSS.n9044 VSS.n9040 4.5005
R3423 VSS.n9030 VSS.n9041 4.57442
R3424 VSS.n9037 VSS.n9038 0.147342
R3425 VSS.n9038 VSS.n9039 0.147342
R3426 VSS.n9039 VSS.n9040 0.147342
R3427 VSS.n9041 VSS.n9042 2.39784
R3428 VSS.n9042 VSS.n9043 0.147342
R3429 VSS.n9043 VSS.n9044 0.147342
R3430 VSS.n9044 VSS.t532 3.13212
R3431 VSS.n9022 VSS.n9017 4.5005
R3432 VSS.n9023 VSS.n9019 4.5005
R3433 VSS.n9024 VSS.n9020 4.5005
R3434 VSS.n9025 VSS.n9021 4.57324
R3435 VSS.n9015 VSS.n9017 0.147342
R3436 VSS.n9018 VSS.n9019 0.0732424
R3437 VSS.n9019 VSS.n9020 0.147342
R3438 VSS.n9026 VSS.n9022 0.0722544
R3439 VSS.n9027 VSS.n9023 4.5005
R3440 VSS.n9028 VSS.n9024 4.5005
R3441 VSS.n9029 VSS.n9025 4.5005
R3442 VSS.n9026 VSS.n9015 4.57426
R3443 VSS.n9022 VSS.n9023 0.147342
R3444 VSS.n9023 VSS.n9024 0.147342
R3445 VSS.n9024 VSS.n9025 0.147342
R3446 VSS.n9027 VSS.n9026 2.37296
R3447 VSS.n9028 VSS.n9027 0.127318
R3448 VSS.n9029 VSS.n9028 0.127318
R3449 VSS.t41 VSS.n9029 2.73618
R3450 VSS.n9002 VSS.n9007 4.5005
R3451 VSS.n9004 VSS.n9008 4.5005
R3452 VSS.n9005 VSS.n9009 4.5005
R3453 VSS.n9006 VSS.n9010 4.57324
R3454 VSS.n9002 VSS.n9000 0.147342
R3455 VSS.n9003 VSS.n9004 0.0732424
R3456 VSS.n9004 VSS.n9005 0.147342
R3457 VSS.n9007 VSS.n9011 0.0721009
R3458 VSS.n9012 VSS.n9008 4.5005
R3459 VSS.n9013 VSS.n9009 4.5005
R3460 VSS.n9014 VSS.n9010 4.5005
R3461 VSS.n9000 VSS.n9011 4.57442
R3462 VSS.n9007 VSS.n9008 0.147342
R3463 VSS.n9008 VSS.n9009 0.147342
R3464 VSS.n9009 VSS.n9010 0.147342
R3465 VSS.n9011 VSS.n9012 2.39784
R3466 VSS.n9012 VSS.n9013 0.147342
R3467 VSS.n9013 VSS.n9014 0.147342
R3468 VSS.n9014 VSS.t149 3.13212
R3469 VSS.n8987 VSS.n8992 4.5005
R3470 VSS.n8989 VSS.n8993 4.5005
R3471 VSS.n8990 VSS.n8994 4.5005
R3472 VSS.n8991 VSS.n8995 4.57324
R3473 VSS.n8987 VSS.n8985 0.147342
R3474 VSS.n8988 VSS.n8989 0.0732424
R3475 VSS.n8989 VSS.n8990 0.147342
R3476 VSS.n8992 VSS.n8996 0.0721009
R3477 VSS.n8997 VSS.n8993 4.5005
R3478 VSS.n8998 VSS.n8994 4.5005
R3479 VSS.n8999 VSS.n8995 4.5005
R3480 VSS.n8985 VSS.n8996 4.57442
R3481 VSS.n8992 VSS.n8993 0.147342
R3482 VSS.n8993 VSS.n8994 0.147342
R3483 VSS.n8994 VSS.n8995 0.147342
R3484 VSS.n8996 VSS.n8997 2.39784
R3485 VSS.n8997 VSS.n8998 0.147342
R3486 VSS.n8998 VSS.n8999 0.147342
R3487 VSS.n8999 VSS.t500 3.13212
R3488 VSS.n8972 VSS.n8977 4.5005
R3489 VSS.n8974 VSS.n8978 4.5005
R3490 VSS.n8975 VSS.n8979 4.5005
R3491 VSS.n8976 VSS.n8980 4.57324
R3492 VSS.n8972 VSS.n8970 0.147342
R3493 VSS.n8973 VSS.n8974 0.0732424
R3494 VSS.n8974 VSS.n8975 0.147342
R3495 VSS.n8977 VSS.n8981 0.0721009
R3496 VSS.n8982 VSS.n8978 4.5005
R3497 VSS.n8983 VSS.n8979 4.5005
R3498 VSS.n8984 VSS.n8980 4.5005
R3499 VSS.n8970 VSS.n8981 4.57442
R3500 VSS.n8977 VSS.n8978 0.147342
R3501 VSS.n8978 VSS.n8979 0.147342
R3502 VSS.n8979 VSS.n8980 0.147342
R3503 VSS.n8981 VSS.n8982 2.39784
R3504 VSS.n8982 VSS.n8983 0.147342
R3505 VSS.n8983 VSS.n8984 0.147342
R3506 VSS.n8984 VSS.t44 3.13212
R3507 VSS.n8957 VSS.n8962 4.5005
R3508 VSS.n8959 VSS.n8963 4.5005
R3509 VSS.n8960 VSS.n8964 4.5005
R3510 VSS.n8961 VSS.n8965 4.57324
R3511 VSS.n8957 VSS.n8955 0.147342
R3512 VSS.n8958 VSS.n8959 0.0732424
R3513 VSS.n8959 VSS.n8960 0.147342
R3514 VSS.n8962 VSS.n8966 0.0721009
R3515 VSS.n8967 VSS.n8963 4.5005
R3516 VSS.n8968 VSS.n8964 4.5005
R3517 VSS.n8969 VSS.n8965 4.5005
R3518 VSS.n8955 VSS.n8966 4.57442
R3519 VSS.n8962 VSS.n8963 0.147342
R3520 VSS.n8963 VSS.n8964 0.147342
R3521 VSS.n8964 VSS.n8965 0.147342
R3522 VSS.n8966 VSS.n8967 2.39784
R3523 VSS.n8967 VSS.n8968 0.147342
R3524 VSS.n8968 VSS.n8969 0.147342
R3525 VSS.n8969 VSS.t606 3.13212
R3526 VSS.n8947 VSS.n8942 4.5005
R3527 VSS.n8948 VSS.n8944 4.5005
R3528 VSS.n8949 VSS.n8945 4.5005
R3529 VSS.n8950 VSS.n8946 4.57324
R3530 VSS.n8940 VSS.n8942 0.147342
R3531 VSS.n8943 VSS.n8944 0.0732424
R3532 VSS.n8944 VSS.n8945 0.147342
R3533 VSS.n8951 VSS.n8947 0.0722544
R3534 VSS.n8952 VSS.n8948 4.5005
R3535 VSS.n8953 VSS.n8949 4.5005
R3536 VSS.n8954 VSS.n8950 4.5005
R3537 VSS.n8951 VSS.n8940 4.57426
R3538 VSS.n8947 VSS.n8948 0.147342
R3539 VSS.n8948 VSS.n8949 0.147342
R3540 VSS.n8949 VSS.n8950 0.147342
R3541 VSS.n8952 VSS.n8951 2.37296
R3542 VSS.n8953 VSS.n8952 0.127318
R3543 VSS.n8954 VSS.n8953 0.127318
R3544 VSS.t41 VSS.n8954 2.73618
R3545 VSS.n8927 VSS.n8932 4.5005
R3546 VSS.n8929 VSS.n8933 4.5005
R3547 VSS.n8930 VSS.n8934 4.5005
R3548 VSS.n8931 VSS.n8935 4.57324
R3549 VSS.n8927 VSS.n8925 0.147342
R3550 VSS.n8928 VSS.n8929 0.0732424
R3551 VSS.n8929 VSS.n8930 0.147342
R3552 VSS.n8932 VSS.n8936 0.0721009
R3553 VSS.n8937 VSS.n8933 4.5005
R3554 VSS.n8938 VSS.n8934 4.5005
R3555 VSS.n8939 VSS.n8935 4.5005
R3556 VSS.n8925 VSS.n8936 4.57442
R3557 VSS.n8932 VSS.n8933 0.147342
R3558 VSS.n8933 VSS.n8934 0.147342
R3559 VSS.n8934 VSS.n8935 0.147342
R3560 VSS.n8936 VSS.n8937 2.39784
R3561 VSS.n8937 VSS.n8938 0.147342
R3562 VSS.n8938 VSS.n8939 0.147342
R3563 VSS.n8939 VSS.t574 3.13212
R3564 VSS.n8912 VSS.n8917 4.5005
R3565 VSS.n8914 VSS.n8918 4.5005
R3566 VSS.n8915 VSS.n8919 4.5005
R3567 VSS.n8916 VSS.n8920 4.57324
R3568 VSS.n8912 VSS.n8910 0.147342
R3569 VSS.n8913 VSS.n8914 0.0732424
R3570 VSS.n8914 VSS.n8915 0.147342
R3571 VSS.n8917 VSS.n8921 0.0721009
R3572 VSS.n8922 VSS.n8918 4.5005
R3573 VSS.n8923 VSS.n8919 4.5005
R3574 VSS.n8924 VSS.n8920 4.5005
R3575 VSS.n8910 VSS.n8921 4.57442
R3576 VSS.n8917 VSS.n8918 0.147342
R3577 VSS.n8918 VSS.n8919 0.147342
R3578 VSS.n8919 VSS.n8920 0.147342
R3579 VSS.n8921 VSS.n8922 2.39784
R3580 VSS.n8922 VSS.n8923 0.147342
R3581 VSS.n8923 VSS.n8924 0.147342
R3582 VSS.n8924 VSS.t198 3.13212
R3583 VSS.n8897 VSS.n8902 4.5005
R3584 VSS.n8899 VSS.n8903 4.5005
R3585 VSS.n8900 VSS.n8904 4.5005
R3586 VSS.n8901 VSS.n8905 4.57324
R3587 VSS.n8897 VSS.n8895 0.147342
R3588 VSS.n8898 VSS.n8899 0.0732424
R3589 VSS.n8899 VSS.n8900 0.147342
R3590 VSS.n8902 VSS.n8906 0.0721009
R3591 VSS.n8907 VSS.n8903 4.5005
R3592 VSS.n8908 VSS.n8904 4.5005
R3593 VSS.n8909 VSS.n8905 4.5005
R3594 VSS.n8895 VSS.n8906 4.57442
R3595 VSS.n8902 VSS.n8903 0.147342
R3596 VSS.n8903 VSS.n8904 0.147342
R3597 VSS.n8904 VSS.n8905 0.147342
R3598 VSS.n8906 VSS.n8907 2.39784
R3599 VSS.n8907 VSS.n8908 0.147342
R3600 VSS.n8908 VSS.n8909 0.147342
R3601 VSS.n8909 VSS.t421 3.13212
R3602 VSS.n8887 VSS.n8882 4.5005
R3603 VSS.n8888 VSS.n8884 4.5005
R3604 VSS.n8889 VSS.n8885 4.5005
R3605 VSS.n8890 VSS.n8886 4.57324
R3606 VSS.n8880 VSS.n8882 0.147342
R3607 VSS.n8883 VSS.n8884 0.0732424
R3608 VSS.n8884 VSS.n8885 0.147342
R3609 VSS.n8891 VSS.n8887 0.0722544
R3610 VSS.n8892 VSS.n8888 4.5005
R3611 VSS.n8893 VSS.n8889 4.5005
R3612 VSS.n8894 VSS.n8890 4.5005
R3613 VSS.n8891 VSS.n8880 4.57426
R3614 VSS.n8887 VSS.n8888 0.147342
R3615 VSS.n8888 VSS.n8889 0.147342
R3616 VSS.n8889 VSS.n8890 0.147342
R3617 VSS.n8892 VSS.n8891 2.37296
R3618 VSS.n8893 VSS.n8892 0.127318
R3619 VSS.n8894 VSS.n8893 0.127318
R3620 VSS.t41 VSS.n8894 2.73618
R3621 VSS.n8867 VSS.n8872 4.5005
R3622 VSS.n8869 VSS.n8873 4.5005
R3623 VSS.n8870 VSS.n8874 4.5005
R3624 VSS.n8871 VSS.n8875 4.57324
R3625 VSS.n8867 VSS.n8865 0.147342
R3626 VSS.n8868 VSS.n8869 0.0732424
R3627 VSS.n8869 VSS.n8870 0.147342
R3628 VSS.n8872 VSS.n8876 0.0721009
R3629 VSS.n8877 VSS.n8873 4.5005
R3630 VSS.n8878 VSS.n8874 4.5005
R3631 VSS.n8879 VSS.n8875 4.5005
R3632 VSS.n8865 VSS.n8876 4.57442
R3633 VSS.n8872 VSS.n8873 0.147342
R3634 VSS.n8873 VSS.n8874 0.147342
R3635 VSS.n8874 VSS.n8875 0.147342
R3636 VSS.n8876 VSS.n8877 2.39784
R3637 VSS.n8877 VSS.n8878 0.147342
R3638 VSS.n8878 VSS.n8879 0.147342
R3639 VSS.n8879 VSS.t557 3.13212
R3640 VSS.n8852 VSS.n8857 4.5005
R3641 VSS.n8854 VSS.n8858 4.5005
R3642 VSS.n8855 VSS.n8859 4.5005
R3643 VSS.n8856 VSS.n8860 4.57324
R3644 VSS.n8852 VSS.n8850 0.147342
R3645 VSS.n8853 VSS.n8854 0.0732424
R3646 VSS.n8854 VSS.n8855 0.147342
R3647 VSS.n8857 VSS.n8861 0.0721009
R3648 VSS.n8862 VSS.n8858 4.5005
R3649 VSS.n8863 VSS.n8859 4.5005
R3650 VSS.n8864 VSS.n8860 4.5005
R3651 VSS.n8850 VSS.n8861 4.57442
R3652 VSS.n8857 VSS.n8858 0.147342
R3653 VSS.n8858 VSS.n8859 0.147342
R3654 VSS.n8859 VSS.n8860 0.147342
R3655 VSS.n8861 VSS.n8862 2.39784
R3656 VSS.n8862 VSS.n8863 0.147342
R3657 VSS.n8863 VSS.n8864 0.147342
R3658 VSS.n8864 VSS.t457 3.13212
R3659 VSS.n8837 VSS.n8842 4.5005
R3660 VSS.n8839 VSS.n8843 4.5005
R3661 VSS.n8840 VSS.n8844 4.5005
R3662 VSS.n8841 VSS.n8845 4.57324
R3663 VSS.n8837 VSS.n8835 0.147342
R3664 VSS.n8838 VSS.n8839 0.0732424
R3665 VSS.n8839 VSS.n8840 0.147342
R3666 VSS.n8842 VSS.n8846 0.0721009
R3667 VSS.n8847 VSS.n8843 4.5005
R3668 VSS.n8848 VSS.n8844 4.5005
R3669 VSS.n8849 VSS.n8845 4.5005
R3670 VSS.n8835 VSS.n8846 4.57442
R3671 VSS.n8842 VSS.n8843 0.147342
R3672 VSS.n8843 VSS.n8844 0.147342
R3673 VSS.n8844 VSS.n8845 0.147342
R3674 VSS.n8846 VSS.n8847 2.39784
R3675 VSS.n8847 VSS.n8848 0.147342
R3676 VSS.n8848 VSS.n8849 0.147342
R3677 VSS.n8849 VSS.t589 3.13212
R3678 VSS.n8822 VSS.n8827 4.5005
R3679 VSS.n8824 VSS.n8828 4.5005
R3680 VSS.n8825 VSS.n8829 4.5005
R3681 VSS.n8826 VSS.n8830 4.57324
R3682 VSS.n8822 VSS.n8820 0.147342
R3683 VSS.n8823 VSS.n8824 0.0732424
R3684 VSS.n8824 VSS.n8825 0.147342
R3685 VSS.n8827 VSS.n8831 0.0721009
R3686 VSS.n8832 VSS.n8828 4.5005
R3687 VSS.n8833 VSS.n8829 4.5005
R3688 VSS.n8834 VSS.n8830 4.5005
R3689 VSS.n8820 VSS.n8831 4.57442
R3690 VSS.n8827 VSS.n8828 0.147342
R3691 VSS.n8828 VSS.n8829 0.147342
R3692 VSS.n8829 VSS.n8830 0.147342
R3693 VSS.n8831 VSS.n8832 2.39784
R3694 VSS.n8832 VSS.n8833 0.147342
R3695 VSS.n8833 VSS.n8834 0.147342
R3696 VSS.n8834 VSS.t68 3.13212
R3697 VSS.n8807 VSS.n8812 4.5005
R3698 VSS.n8809 VSS.n8813 4.5005
R3699 VSS.n8810 VSS.n8814 4.5005
R3700 VSS.n8811 VSS.n8815 4.57324
R3701 VSS.n8807 VSS.n8805 0.147342
R3702 VSS.n8808 VSS.n8809 0.0732424
R3703 VSS.n8809 VSS.n8810 0.147342
R3704 VSS.n8812 VSS.n8816 0.0721009
R3705 VSS.n8817 VSS.n8813 4.5005
R3706 VSS.n8818 VSS.n8814 4.5005
R3707 VSS.n8819 VSS.n8815 4.5005
R3708 VSS.n8805 VSS.n8816 4.57442
R3709 VSS.n8812 VSS.n8813 0.147342
R3710 VSS.n8813 VSS.n8814 0.147342
R3711 VSS.n8814 VSS.n8815 0.147342
R3712 VSS.n8816 VSS.n8817 2.39784
R3713 VSS.n8817 VSS.n8818 0.147342
R3714 VSS.n8818 VSS.n8819 0.147342
R3715 VSS.n8819 VSS.t78 3.13212
R3716 VSS.n8792 VSS.n8797 4.5005
R3717 VSS.n8794 VSS.n8798 4.5005
R3718 VSS.n8795 VSS.n8799 4.5005
R3719 VSS.n8796 VSS.n8800 4.57324
R3720 VSS.n8792 VSS.n8790 0.147342
R3721 VSS.n8793 VSS.n8794 0.0732424
R3722 VSS.n8794 VSS.n8795 0.147342
R3723 VSS.n8797 VSS.n8801 0.0721009
R3724 VSS.n8802 VSS.n8798 4.5005
R3725 VSS.n8803 VSS.n8799 4.5005
R3726 VSS.n8804 VSS.n8800 4.5005
R3727 VSS.n8790 VSS.n8801 4.57442
R3728 VSS.n8797 VSS.n8798 0.147342
R3729 VSS.n8798 VSS.n8799 0.147342
R3730 VSS.n8799 VSS.n8800 0.147342
R3731 VSS.n8801 VSS.n8802 2.39784
R3732 VSS.n8802 VSS.n8803 0.147342
R3733 VSS.n8803 VSS.n8804 0.147342
R3734 VSS.n8804 VSS.t450 3.13212
R3735 VSS.n8782 VSS.n8777 4.5005
R3736 VSS.n8783 VSS.n8779 4.5005
R3737 VSS.n8784 VSS.n8780 4.5005
R3738 VSS.n8785 VSS.n8781 4.57324
R3739 VSS.n8775 VSS.n8777 0.147342
R3740 VSS.n8778 VSS.n8779 0.0732424
R3741 VSS.n8779 VSS.n8780 0.147342
R3742 VSS.n8786 VSS.n8782 0.0722544
R3743 VSS.n8787 VSS.n8783 4.5005
R3744 VSS.n8788 VSS.n8784 4.5005
R3745 VSS.n8789 VSS.n8785 4.5005
R3746 VSS.n8786 VSS.n8775 4.57426
R3747 VSS.n8782 VSS.n8783 0.147342
R3748 VSS.n8783 VSS.n8784 0.147342
R3749 VSS.n8784 VSS.n8785 0.147342
R3750 VSS.n8787 VSS.n8786 2.37296
R3751 VSS.n8788 VSS.n8787 0.127318
R3752 VSS.n8789 VSS.n8788 0.127318
R3753 VSS.t41 VSS.n8789 2.73618
R3754 VSS.n8762 VSS.n8767 4.5005
R3755 VSS.n8764 VSS.n8768 4.5005
R3756 VSS.n8765 VSS.n8769 4.5005
R3757 VSS.n8766 VSS.n8770 4.57324
R3758 VSS.n8762 VSS.n8760 0.147342
R3759 VSS.n8763 VSS.n8764 0.0732424
R3760 VSS.n8764 VSS.n8765 0.147342
R3761 VSS.n8767 VSS.n8771 0.0721009
R3762 VSS.n8772 VSS.n8768 4.5005
R3763 VSS.n8773 VSS.n8769 4.5005
R3764 VSS.n8774 VSS.n8770 4.5005
R3765 VSS.n8760 VSS.n8771 4.57442
R3766 VSS.n8767 VSS.n8768 0.147342
R3767 VSS.n8768 VSS.n8769 0.147342
R3768 VSS.n8769 VSS.n8770 0.147342
R3769 VSS.n8771 VSS.n8772 2.39784
R3770 VSS.n8772 VSS.n8773 0.147342
R3771 VSS.n8773 VSS.n8774 0.147342
R3772 VSS.n8774 VSS.t613 3.13212
R3773 VSS.n8747 VSS.n8752 4.5005
R3774 VSS.n8749 VSS.n8753 4.5005
R3775 VSS.n8750 VSS.n8754 4.5005
R3776 VSS.n8751 VSS.n8755 4.57324
R3777 VSS.n8747 VSS.n8745 0.147342
R3778 VSS.n8748 VSS.n8749 0.0732424
R3779 VSS.n8749 VSS.n8750 0.147342
R3780 VSS.n8752 VSS.n8756 0.0721009
R3781 VSS.n8757 VSS.n8753 4.5005
R3782 VSS.n8758 VSS.n8754 4.5005
R3783 VSS.n8759 VSS.n8755 4.5005
R3784 VSS.n8745 VSS.n8756 4.57442
R3785 VSS.n8752 VSS.n8753 0.147342
R3786 VSS.n8753 VSS.n8754 0.147342
R3787 VSS.n8754 VSS.n8755 0.147342
R3788 VSS.n8756 VSS.n8757 2.39784
R3789 VSS.n8757 VSS.n8758 0.147342
R3790 VSS.n8758 VSS.n8759 0.147342
R3791 VSS.n8759 VSS.t53 3.13212
R3792 VSS.n8732 VSS.n8737 4.5005
R3793 VSS.n8734 VSS.n8738 4.5005
R3794 VSS.n8735 VSS.n8739 4.5005
R3795 VSS.n8736 VSS.n8740 4.57324
R3796 VSS.n8732 VSS.n8730 0.147342
R3797 VSS.n8733 VSS.n8734 0.0732424
R3798 VSS.n8734 VSS.n8735 0.147342
R3799 VSS.n8737 VSS.n8741 0.0721009
R3800 VSS.n8742 VSS.n8738 4.5005
R3801 VSS.n8743 VSS.n8739 4.5005
R3802 VSS.n8744 VSS.n8740 4.5005
R3803 VSS.n8730 VSS.n8741 4.57442
R3804 VSS.n8737 VSS.n8738 0.147342
R3805 VSS.n8738 VSS.n8739 0.147342
R3806 VSS.n8739 VSS.n8740 0.147342
R3807 VSS.n8741 VSS.n8742 2.39784
R3808 VSS.n8742 VSS.n8743 0.147342
R3809 VSS.n8743 VSS.n8744 0.147342
R3810 VSS.n8744 VSS.t534 3.13212
R3811 VSS.n8722 VSS.n8717 4.5005
R3812 VSS.n8723 VSS.n8719 4.5005
R3813 VSS.n8724 VSS.n8720 4.5005
R3814 VSS.n8725 VSS.n8721 4.57324
R3815 VSS.n8715 VSS.n8717 0.147342
R3816 VSS.n8718 VSS.n8719 0.0732424
R3817 VSS.n8719 VSS.n8720 0.147342
R3818 VSS.n8726 VSS.n8722 0.0722544
R3819 VSS.n8727 VSS.n8723 4.5005
R3820 VSS.n8728 VSS.n8724 4.5005
R3821 VSS.n8729 VSS.n8725 4.5005
R3822 VSS.n8726 VSS.n8715 4.57426
R3823 VSS.n8722 VSS.n8723 0.147342
R3824 VSS.n8723 VSS.n8724 0.147342
R3825 VSS.n8724 VSS.n8725 0.147342
R3826 VSS.n8727 VSS.n8726 2.37296
R3827 VSS.n8728 VSS.n8727 0.127318
R3828 VSS.n8729 VSS.n8728 0.127318
R3829 VSS.t41 VSS.n8729 2.73618
R3830 VSS.n8702 VSS.n8707 4.5005
R3831 VSS.n8704 VSS.n8708 4.5005
R3832 VSS.n8705 VSS.n8709 4.5005
R3833 VSS.n8706 VSS.n8710 4.57324
R3834 VSS.n8702 VSS.n8700 0.147342
R3835 VSS.n8703 VSS.n8704 0.0732424
R3836 VSS.n8704 VSS.n8705 0.147342
R3837 VSS.n8707 VSS.n8711 0.0721009
R3838 VSS.n8712 VSS.n8708 4.5005
R3839 VSS.n8713 VSS.n8709 4.5005
R3840 VSS.n8714 VSS.n8710 4.5005
R3841 VSS.n8700 VSS.n8711 4.57442
R3842 VSS.n8707 VSS.n8708 0.147342
R3843 VSS.n8708 VSS.n8709 0.147342
R3844 VSS.n8709 VSS.n8710 0.147342
R3845 VSS.n8711 VSS.n8712 2.39784
R3846 VSS.n8712 VSS.n8713 0.147342
R3847 VSS.n8713 VSS.n8714 0.147342
R3848 VSS.n8714 VSS.t150 3.13212
R3849 VSS.n8687 VSS.n8692 4.5005
R3850 VSS.n8689 VSS.n8693 4.5005
R3851 VSS.n8690 VSS.n8694 4.5005
R3852 VSS.n8691 VSS.n8695 4.57324
R3853 VSS.n8687 VSS.n8685 0.147342
R3854 VSS.n8688 VSS.n8689 0.0732424
R3855 VSS.n8689 VSS.n8690 0.147342
R3856 VSS.n8692 VSS.n8696 0.0721009
R3857 VSS.n8697 VSS.n8693 4.5005
R3858 VSS.n8698 VSS.n8694 4.5005
R3859 VSS.n8699 VSS.n8695 4.5005
R3860 VSS.n8685 VSS.n8696 4.57442
R3861 VSS.n8692 VSS.n8693 0.147342
R3862 VSS.n8693 VSS.n8694 0.147342
R3863 VSS.n8694 VSS.n8695 0.147342
R3864 VSS.n8696 VSS.n8697 2.39784
R3865 VSS.n8697 VSS.n8698 0.147342
R3866 VSS.n8698 VSS.n8699 0.147342
R3867 VSS.n8699 VSS.t472 3.13212
R3868 VSS.n8672 VSS.n8677 4.5005
R3869 VSS.n8674 VSS.n8678 4.5005
R3870 VSS.n8675 VSS.n8679 4.5005
R3871 VSS.n8676 VSS.n8680 4.57324
R3872 VSS.n8672 VSS.n8670 0.147342
R3873 VSS.n8673 VSS.n8674 0.0732424
R3874 VSS.n8674 VSS.n8675 0.147342
R3875 VSS.n8677 VSS.n8681 0.0721009
R3876 VSS.n8682 VSS.n8678 4.5005
R3877 VSS.n8683 VSS.n8679 4.5005
R3878 VSS.n8684 VSS.n8680 4.5005
R3879 VSS.n8670 VSS.n8681 4.57442
R3880 VSS.n8677 VSS.n8678 0.147342
R3881 VSS.n8678 VSS.n8679 0.147342
R3882 VSS.n8679 VSS.n8680 0.147342
R3883 VSS.n8681 VSS.n8682 2.39784
R3884 VSS.n8682 VSS.n8683 0.147342
R3885 VSS.n8683 VSS.n8684 0.147342
R3886 VSS.n8684 VSS.t42 3.13212
R3887 VSS.n8657 VSS.n8662 4.5005
R3888 VSS.n8659 VSS.n8663 4.5005
R3889 VSS.n8660 VSS.n8664 4.5005
R3890 VSS.n8661 VSS.n8665 4.57324
R3891 VSS.n8657 VSS.n8655 0.147342
R3892 VSS.n8658 VSS.n8659 0.0732424
R3893 VSS.n8659 VSS.n8660 0.147342
R3894 VSS.n8662 VSS.n8666 0.0721009
R3895 VSS.n8667 VSS.n8663 4.5005
R3896 VSS.n8668 VSS.n8664 4.5005
R3897 VSS.n8669 VSS.n8665 4.5005
R3898 VSS.n8655 VSS.n8666 4.57442
R3899 VSS.n8662 VSS.n8663 0.147342
R3900 VSS.n8663 VSS.n8664 0.147342
R3901 VSS.n8664 VSS.n8665 0.147342
R3902 VSS.n8666 VSS.n8667 2.39784
R3903 VSS.n8667 VSS.n8668 0.147342
R3904 VSS.n8668 VSS.n8669 0.147342
R3905 VSS.n8669 VSS.t608 3.13212
R3906 VSS.n8647 VSS.n8642 4.5005
R3907 VSS.n8648 VSS.n8644 4.5005
R3908 VSS.n8649 VSS.n8645 4.5005
R3909 VSS.n8650 VSS.n8646 4.57324
R3910 VSS.n8640 VSS.n8642 0.147342
R3911 VSS.n8643 VSS.n8644 0.0732424
R3912 VSS.n8644 VSS.n8645 0.147342
R3913 VSS.n8651 VSS.n8647 0.0722544
R3914 VSS.n8652 VSS.n8648 4.5005
R3915 VSS.n8653 VSS.n8649 4.5005
R3916 VSS.n8654 VSS.n8650 4.5005
R3917 VSS.n8651 VSS.n8640 4.57426
R3918 VSS.n8647 VSS.n8648 0.147342
R3919 VSS.n8648 VSS.n8649 0.147342
R3920 VSS.n8649 VSS.n8650 0.147342
R3921 VSS.n8652 VSS.n8651 2.37296
R3922 VSS.n8653 VSS.n8652 0.127318
R3923 VSS.n8654 VSS.n8653 0.127318
R3924 VSS.t41 VSS.n8654 2.73618
R3925 VSS.n8627 VSS.n8632 4.5005
R3926 VSS.n8629 VSS.n8633 4.5005
R3927 VSS.n8630 VSS.n8634 4.5005
R3928 VSS.n8631 VSS.n8635 4.57324
R3929 VSS.n8627 VSS.n8625 0.147342
R3930 VSS.n8628 VSS.n8629 0.0732424
R3931 VSS.n8629 VSS.n8630 0.147342
R3932 VSS.n8632 VSS.n8636 0.0721009
R3933 VSS.n8637 VSS.n8633 4.5005
R3934 VSS.n8638 VSS.n8634 4.5005
R3935 VSS.n8639 VSS.n8635 4.5005
R3936 VSS.n8625 VSS.n8636 4.57442
R3937 VSS.n8632 VSS.n8633 0.147342
R3938 VSS.n8633 VSS.n8634 0.147342
R3939 VSS.n8634 VSS.n8635 0.147342
R3940 VSS.n8636 VSS.n8637 2.39784
R3941 VSS.n8637 VSS.n8638 0.147342
R3942 VSS.n8638 VSS.n8639 0.147342
R3943 VSS.n8639 VSS.t577 3.13212
R3944 VSS.n8612 VSS.n8617 4.5005
R3945 VSS.n8614 VSS.n8618 4.5005
R3946 VSS.n8615 VSS.n8619 4.5005
R3947 VSS.n8616 VSS.n8620 4.57324
R3948 VSS.n8612 VSS.n8610 0.147342
R3949 VSS.n8613 VSS.n8614 0.0732424
R3950 VSS.n8614 VSS.n8615 0.147342
R3951 VSS.n8617 VSS.n8621 0.0721009
R3952 VSS.n8622 VSS.n8618 4.5005
R3953 VSS.n8623 VSS.n8619 4.5005
R3954 VSS.n8624 VSS.n8620 4.5005
R3955 VSS.n8610 VSS.n8621 4.57442
R3956 VSS.n8617 VSS.n8618 0.147342
R3957 VSS.n8618 VSS.n8619 0.147342
R3958 VSS.n8619 VSS.n8620 0.147342
R3959 VSS.n8621 VSS.n8622 2.39784
R3960 VSS.n8622 VSS.n8623 0.147342
R3961 VSS.n8623 VSS.n8624 0.147342
R3962 VSS.n8624 VSS.t200 3.13212
R3963 VSS.n8597 VSS.n8602 4.5005
R3964 VSS.n8599 VSS.n8603 4.5005
R3965 VSS.n8600 VSS.n8604 4.5005
R3966 VSS.n8601 VSS.n8605 4.57324
R3967 VSS.n8597 VSS.n8595 0.147342
R3968 VSS.n8598 VSS.n8599 0.0732424
R3969 VSS.n8599 VSS.n8600 0.147342
R3970 VSS.n8602 VSS.n8606 0.0721009
R3971 VSS.n8607 VSS.n8603 4.5005
R3972 VSS.n8608 VSS.n8604 4.5005
R3973 VSS.n8609 VSS.n8605 4.5005
R3974 VSS.n8595 VSS.n8606 4.57442
R3975 VSS.n8602 VSS.n8603 0.147342
R3976 VSS.n8603 VSS.n8604 0.147342
R3977 VSS.n8604 VSS.n8605 0.147342
R3978 VSS.n8606 VSS.n8607 2.39784
R3979 VSS.n8607 VSS.n8608 0.147342
R3980 VSS.n8608 VSS.n8609 0.147342
R3981 VSS.n8609 VSS.t410 3.13212
R3982 VSS.n8587 VSS.n8582 4.5005
R3983 VSS.n8588 VSS.n8584 4.5005
R3984 VSS.n8589 VSS.n8585 4.5005
R3985 VSS.n8590 VSS.n8586 4.57324
R3986 VSS.n8580 VSS.n8582 0.147342
R3987 VSS.n8583 VSS.n8584 0.0732424
R3988 VSS.n8584 VSS.n8585 0.147342
R3989 VSS.n8591 VSS.n8587 0.0722544
R3990 VSS.n8592 VSS.n8588 4.5005
R3991 VSS.n8593 VSS.n8589 4.5005
R3992 VSS.n8594 VSS.n8590 4.5005
R3993 VSS.n8591 VSS.n8580 4.57426
R3994 VSS.n8587 VSS.n8588 0.147342
R3995 VSS.n8588 VSS.n8589 0.147342
R3996 VSS.n8589 VSS.n8590 0.147342
R3997 VSS.n8592 VSS.n8591 2.37296
R3998 VSS.n8593 VSS.n8592 0.127318
R3999 VSS.n8594 VSS.n8593 0.127318
R4000 VSS.t41 VSS.n8594 2.73618
R4001 VSS.n8567 VSS.n8572 4.5005
R4002 VSS.n8569 VSS.n8573 4.5005
R4003 VSS.n8570 VSS.n8574 4.5005
R4004 VSS.n8571 VSS.n8575 4.57324
R4005 VSS.n8567 VSS.n8565 0.147342
R4006 VSS.n8568 VSS.n8569 0.0732424
R4007 VSS.n8569 VSS.n8570 0.147342
R4008 VSS.n8572 VSS.n8576 0.0721009
R4009 VSS.n8577 VSS.n8573 4.5005
R4010 VSS.n8578 VSS.n8574 4.5005
R4011 VSS.n8579 VSS.n8575 4.5005
R4012 VSS.n8565 VSS.n8576 4.57442
R4013 VSS.n8572 VSS.n8573 0.147342
R4014 VSS.n8573 VSS.n8574 0.147342
R4015 VSS.n8574 VSS.n8575 0.147342
R4016 VSS.n8576 VSS.n8577 2.39784
R4017 VSS.n8577 VSS.n8578 0.147342
R4018 VSS.n8578 VSS.n8579 0.147342
R4019 VSS.n8579 VSS.t554 3.13212
R4020 VSS.n8552 VSS.n8557 4.5005
R4021 VSS.n8554 VSS.n8558 4.5005
R4022 VSS.n8555 VSS.n8559 4.5005
R4023 VSS.n8556 VSS.n8560 4.57324
R4024 VSS.n8552 VSS.n8550 0.147342
R4025 VSS.n8553 VSS.n8554 0.0732424
R4026 VSS.n8554 VSS.n8555 0.147342
R4027 VSS.n8557 VSS.n8561 0.0721009
R4028 VSS.n8562 VSS.n8558 4.5005
R4029 VSS.n8563 VSS.n8559 4.5005
R4030 VSS.n8564 VSS.n8560 4.5005
R4031 VSS.n8550 VSS.n8561 4.57442
R4032 VSS.n8557 VSS.n8558 0.147342
R4033 VSS.n8558 VSS.n8559 0.147342
R4034 VSS.n8559 VSS.n8560 0.147342
R4035 VSS.n8561 VSS.n8562 2.39784
R4036 VSS.n8562 VSS.n8563 0.147342
R4037 VSS.n8563 VSS.n8564 0.147342
R4038 VSS.n8564 VSS.t601 3.13212
R4039 VSS.n8537 VSS.n8542 4.5005
R4040 VSS.n8539 VSS.n8543 4.5005
R4041 VSS.n8540 VSS.n8544 4.5005
R4042 VSS.n8541 VSS.n8545 4.57324
R4043 VSS.n8537 VSS.n8535 0.147342
R4044 VSS.n8538 VSS.n8539 0.0732424
R4045 VSS.n8539 VSS.n8540 0.147342
R4046 VSS.n8542 VSS.n8546 0.0721009
R4047 VSS.n8547 VSS.n8543 4.5005
R4048 VSS.n8548 VSS.n8544 4.5005
R4049 VSS.n8549 VSS.n8545 4.5005
R4050 VSS.n8535 VSS.n8546 4.57442
R4051 VSS.n8542 VSS.n8543 0.147342
R4052 VSS.n8543 VSS.n8544 0.147342
R4053 VSS.n8544 VSS.n8545 0.147342
R4054 VSS.n8546 VSS.n8547 2.39784
R4055 VSS.n8547 VSS.n8548 0.147342
R4056 VSS.n8548 VSS.n8549 0.147342
R4057 VSS.n8549 VSS.t590 3.13212
R4058 VSS.n8522 VSS.n8527 4.5005
R4059 VSS.n8524 VSS.n8528 4.5005
R4060 VSS.n8525 VSS.n8529 4.5005
R4061 VSS.n8526 VSS.n8530 4.57324
R4062 VSS.n8522 VSS.n8520 0.147342
R4063 VSS.n8523 VSS.n8524 0.0732424
R4064 VSS.n8524 VSS.n8525 0.147342
R4065 VSS.n8527 VSS.n8531 0.0721009
R4066 VSS.n8532 VSS.n8528 4.5005
R4067 VSS.n8533 VSS.n8529 4.5005
R4068 VSS.n8534 VSS.n8530 4.5005
R4069 VSS.n8520 VSS.n8531 4.57442
R4070 VSS.n8527 VSS.n8528 0.147342
R4071 VSS.n8528 VSS.n8529 0.147342
R4072 VSS.n8529 VSS.n8530 0.147342
R4073 VSS.n8531 VSS.n8532 2.39784
R4074 VSS.n8532 VSS.n8533 0.147342
R4075 VSS.n8533 VSS.n8534 0.147342
R4076 VSS.n8534 VSS.t488 3.13212
R4077 VSS.n8507 VSS.n8512 4.5005
R4078 VSS.n8509 VSS.n8513 4.5005
R4079 VSS.n8510 VSS.n8514 4.5005
R4080 VSS.n8511 VSS.n8515 4.57324
R4081 VSS.n8507 VSS.n8505 0.147342
R4082 VSS.n8508 VSS.n8509 0.0732424
R4083 VSS.n8509 VSS.n8510 0.147342
R4084 VSS.n8512 VSS.n8516 0.0721009
R4085 VSS.n8517 VSS.n8513 4.5005
R4086 VSS.n8518 VSS.n8514 4.5005
R4087 VSS.n8519 VSS.n8515 4.5005
R4088 VSS.n8505 VSS.n8516 4.57442
R4089 VSS.n8512 VSS.n8513 0.147342
R4090 VSS.n8513 VSS.n8514 0.147342
R4091 VSS.n8514 VSS.n8515 0.147342
R4092 VSS.n8516 VSS.n8517 2.39784
R4093 VSS.n8517 VSS.n8518 0.147342
R4094 VSS.n8518 VSS.n8519 0.147342
R4095 VSS.n8519 VSS.t115 3.13212
R4096 VSS.n8492 VSS.n8497 4.5005
R4097 VSS.n8494 VSS.n8498 4.5005
R4098 VSS.n8495 VSS.n8499 4.5005
R4099 VSS.n8496 VSS.n8500 4.57324
R4100 VSS.n8492 VSS.n8490 0.147342
R4101 VSS.n8493 VSS.n8494 0.0732424
R4102 VSS.n8494 VSS.n8495 0.147342
R4103 VSS.n8497 VSS.n8501 0.0721009
R4104 VSS.n8502 VSS.n8498 4.5005
R4105 VSS.n8503 VSS.n8499 4.5005
R4106 VSS.n8504 VSS.n8500 4.5005
R4107 VSS.n8490 VSS.n8501 4.57442
R4108 VSS.n8497 VSS.n8498 0.147342
R4109 VSS.n8498 VSS.n8499 0.147342
R4110 VSS.n8499 VSS.n8500 0.147342
R4111 VSS.n8501 VSS.n8502 2.39784
R4112 VSS.n8502 VSS.n8503 0.147342
R4113 VSS.n8503 VSS.n8504 0.147342
R4114 VSS.n8504 VSS.t446 3.13212
R4115 VSS.n8482 VSS.n8477 4.5005
R4116 VSS.n8483 VSS.n8479 4.5005
R4117 VSS.n8484 VSS.n8480 4.5005
R4118 VSS.n8485 VSS.n8481 4.57324
R4119 VSS.n8475 VSS.n8477 0.147342
R4120 VSS.n8478 VSS.n8479 0.0732424
R4121 VSS.n8479 VSS.n8480 0.147342
R4122 VSS.n8486 VSS.n8482 0.0722544
R4123 VSS.n8487 VSS.n8483 4.5005
R4124 VSS.n8488 VSS.n8484 4.5005
R4125 VSS.n8489 VSS.n8485 4.5005
R4126 VSS.n8486 VSS.n8475 4.57426
R4127 VSS.n8482 VSS.n8483 0.147342
R4128 VSS.n8483 VSS.n8484 0.147342
R4129 VSS.n8484 VSS.n8485 0.147342
R4130 VSS.n8487 VSS.n8486 2.37296
R4131 VSS.n8488 VSS.n8487 0.127318
R4132 VSS.n8489 VSS.n8488 0.127318
R4133 VSS.t41 VSS.n8489 2.73618
R4134 VSS.n8462 VSS.n8467 4.5005
R4135 VSS.n8464 VSS.n8468 4.5005
R4136 VSS.n8465 VSS.n8469 4.5005
R4137 VSS.n8466 VSS.n8470 4.57324
R4138 VSS.n8462 VSS.n8460 0.147342
R4139 VSS.n8463 VSS.n8464 0.0732424
R4140 VSS.n8464 VSS.n8465 0.147342
R4141 VSS.n8467 VSS.n8471 0.0721009
R4142 VSS.n8472 VSS.n8468 4.5005
R4143 VSS.n8473 VSS.n8469 4.5005
R4144 VSS.n8474 VSS.n8470 4.5005
R4145 VSS.n8460 VSS.n8471 4.57442
R4146 VSS.n8467 VSS.n8468 0.147342
R4147 VSS.n8468 VSS.n8469 0.147342
R4148 VSS.n8469 VSS.n8470 0.147342
R4149 VSS.n8471 VSS.n8472 2.39784
R4150 VSS.n8472 VSS.n8473 0.147342
R4151 VSS.n8473 VSS.n8474 0.147342
R4152 VSS.n8474 VSS.t618 3.13212
R4153 VSS.n8447 VSS.n8452 4.5005
R4154 VSS.n8449 VSS.n8453 4.5005
R4155 VSS.n8450 VSS.n8454 4.5005
R4156 VSS.n8451 VSS.n8455 4.57324
R4157 VSS.n8447 VSS.n8445 0.147342
R4158 VSS.n8448 VSS.n8449 0.0732424
R4159 VSS.n8449 VSS.n8450 0.147342
R4160 VSS.n8452 VSS.n8456 0.0721009
R4161 VSS.n8457 VSS.n8453 4.5005
R4162 VSS.n8458 VSS.n8454 4.5005
R4163 VSS.n8459 VSS.n8455 4.5005
R4164 VSS.n8445 VSS.n8456 4.57442
R4165 VSS.n8452 VSS.n8453 0.147342
R4166 VSS.n8453 VSS.n8454 0.147342
R4167 VSS.n8454 VSS.n8455 0.147342
R4168 VSS.n8456 VSS.n8457 2.39784
R4169 VSS.n8457 VSS.n8458 0.147342
R4170 VSS.n8458 VSS.n8459 0.147342
R4171 VSS.n8459 VSS.t520 3.13212
R4172 VSS.n8432 VSS.n8437 4.5005
R4173 VSS.n8434 VSS.n8438 4.5005
R4174 VSS.n8435 VSS.n8439 4.5005
R4175 VSS.n8436 VSS.n8440 4.57324
R4176 VSS.n8432 VSS.n8430 0.147342
R4177 VSS.n8433 VSS.n8434 0.0732424
R4178 VSS.n8434 VSS.n8435 0.147342
R4179 VSS.n8437 VSS.n8441 0.0721009
R4180 VSS.n8442 VSS.n8438 4.5005
R4181 VSS.n8443 VSS.n8439 4.5005
R4182 VSS.n8444 VSS.n8440 4.5005
R4183 VSS.n8430 VSS.n8441 4.57442
R4184 VSS.n8437 VSS.n8438 0.147342
R4185 VSS.n8438 VSS.n8439 0.147342
R4186 VSS.n8439 VSS.n8440 0.147342
R4187 VSS.n8441 VSS.n8442 2.39784
R4188 VSS.n8442 VSS.n8443 0.147342
R4189 VSS.n8443 VSS.n8444 0.147342
R4190 VSS.n8444 VSS.t525 3.13212
R4191 VSS.n8422 VSS.n8417 4.5005
R4192 VSS.n8423 VSS.n8419 4.5005
R4193 VSS.n8424 VSS.n8420 4.5005
R4194 VSS.n8425 VSS.n8421 4.57324
R4195 VSS.n8415 VSS.n8417 0.147342
R4196 VSS.n8418 VSS.n8419 0.0732424
R4197 VSS.n8419 VSS.n8420 0.147342
R4198 VSS.n8426 VSS.n8422 0.0722544
R4199 VSS.n8427 VSS.n8423 4.5005
R4200 VSS.n8428 VSS.n8424 4.5005
R4201 VSS.n8429 VSS.n8425 4.5005
R4202 VSS.n8426 VSS.n8415 4.57426
R4203 VSS.n8422 VSS.n8423 0.147342
R4204 VSS.n8423 VSS.n8424 0.147342
R4205 VSS.n8424 VSS.n8425 0.147342
R4206 VSS.n8427 VSS.n8426 2.37296
R4207 VSS.n8428 VSS.n8427 0.127318
R4208 VSS.n8429 VSS.n8428 0.127318
R4209 VSS.t41 VSS.n8429 2.73618
R4210 VSS.n8402 VSS.n8407 4.5005
R4211 VSS.n8404 VSS.n8408 4.5005
R4212 VSS.n8405 VSS.n8409 4.5005
R4213 VSS.n8406 VSS.n8410 4.57324
R4214 VSS.n8402 VSS.n8400 0.147342
R4215 VSS.n8403 VSS.n8404 0.0732424
R4216 VSS.n8404 VSS.n8405 0.147342
R4217 VSS.n8407 VSS.n8411 0.0721009
R4218 VSS.n8412 VSS.n8408 4.5005
R4219 VSS.n8413 VSS.n8409 4.5005
R4220 VSS.n8414 VSS.n8410 4.5005
R4221 VSS.n8400 VSS.n8411 4.57442
R4222 VSS.n8407 VSS.n8408 0.147342
R4223 VSS.n8408 VSS.n8409 0.147342
R4224 VSS.n8409 VSS.n8410 0.147342
R4225 VSS.n8411 VSS.n8412 2.39784
R4226 VSS.n8412 VSS.n8413 0.147342
R4227 VSS.n8413 VSS.n8414 0.147342
R4228 VSS.n8414 VSS.t112 3.13212
R4229 VSS.n8387 VSS.n8392 4.5005
R4230 VSS.n8389 VSS.n8393 4.5005
R4231 VSS.n8390 VSS.n8394 4.5005
R4232 VSS.n8391 VSS.n8395 4.57324
R4233 VSS.n8387 VSS.n8385 0.147342
R4234 VSS.n8388 VSS.n8389 0.0732424
R4235 VSS.n8389 VSS.n8390 0.147342
R4236 VSS.n8392 VSS.n8396 0.0721009
R4237 VSS.n8397 VSS.n8393 4.5005
R4238 VSS.n8398 VSS.n8394 4.5005
R4239 VSS.n8399 VSS.n8395 4.5005
R4240 VSS.n8385 VSS.n8396 4.57442
R4241 VSS.n8392 VSS.n8393 0.147342
R4242 VSS.n8393 VSS.n8394 0.147342
R4243 VSS.n8394 VSS.n8395 0.147342
R4244 VSS.n8396 VSS.n8397 2.39784
R4245 VSS.n8397 VSS.n8398 0.147342
R4246 VSS.n8398 VSS.n8399 0.147342
R4247 VSS.n8399 VSS.t474 3.13212
R4248 VSS.n8372 VSS.n8377 4.5005
R4249 VSS.n8374 VSS.n8378 4.5005
R4250 VSS.n8375 VSS.n8379 4.5005
R4251 VSS.n8376 VSS.n8380 4.57324
R4252 VSS.n8372 VSS.n8370 0.147342
R4253 VSS.n8373 VSS.n8374 0.0732424
R4254 VSS.n8374 VSS.n8375 0.147342
R4255 VSS.n8377 VSS.n8381 0.0721009
R4256 VSS.n8382 VSS.n8378 4.5005
R4257 VSS.n8383 VSS.n8379 4.5005
R4258 VSS.n8384 VSS.n8380 4.5005
R4259 VSS.n8370 VSS.n8381 4.57442
R4260 VSS.n8377 VSS.n8378 0.147342
R4261 VSS.n8378 VSS.n8379 0.147342
R4262 VSS.n8379 VSS.n8380 0.147342
R4263 VSS.n8381 VSS.n8382 2.39784
R4264 VSS.n8382 VSS.n8383 0.147342
R4265 VSS.n8383 VSS.n8384 0.147342
R4266 VSS.n8384 VSS.t45 3.13212
R4267 VSS.n8357 VSS.n8362 4.5005
R4268 VSS.n8359 VSS.n8363 4.5005
R4269 VSS.n8360 VSS.n8364 4.5005
R4270 VSS.n8361 VSS.n8365 4.57324
R4271 VSS.n8357 VSS.n8355 0.147342
R4272 VSS.n8358 VSS.n8359 0.0732424
R4273 VSS.n8359 VSS.n8360 0.147342
R4274 VSS.n8362 VSS.n8366 0.0721009
R4275 VSS.n8367 VSS.n8363 4.5005
R4276 VSS.n8368 VSS.n8364 4.5005
R4277 VSS.n8369 VSS.n8365 4.5005
R4278 VSS.n8355 VSS.n8366 4.57442
R4279 VSS.n8362 VSS.n8363 0.147342
R4280 VSS.n8363 VSS.n8364 0.147342
R4281 VSS.n8364 VSS.n8365 0.147342
R4282 VSS.n8366 VSS.n8367 2.39784
R4283 VSS.n8367 VSS.n8368 0.147342
R4284 VSS.n8368 VSS.n8369 0.147342
R4285 VSS.n8369 VSS.t507 3.13212
R4286 VSS.n8347 VSS.n8342 4.5005
R4287 VSS.n8348 VSS.n8344 4.5005
R4288 VSS.n8349 VSS.n8345 4.5005
R4289 VSS.n8350 VSS.n8346 4.57324
R4290 VSS.n8340 VSS.n8342 0.147342
R4291 VSS.n8343 VSS.n8344 0.0732424
R4292 VSS.n8344 VSS.n8345 0.147342
R4293 VSS.n8351 VSS.n8347 0.0722544
R4294 VSS.n8352 VSS.n8348 4.5005
R4295 VSS.n8353 VSS.n8349 4.5005
R4296 VSS.n8354 VSS.n8350 4.5005
R4297 VSS.n8351 VSS.n8340 4.57426
R4298 VSS.n8347 VSS.n8348 0.147342
R4299 VSS.n8348 VSS.n8349 0.147342
R4300 VSS.n8349 VSS.n8350 0.147342
R4301 VSS.n8352 VSS.n8351 2.37296
R4302 VSS.n8353 VSS.n8352 0.127318
R4303 VSS.n8354 VSS.n8353 0.127318
R4304 VSS.t41 VSS.n8354 2.73618
R4305 VSS.n8327 VSS.n8332 4.5005
R4306 VSS.n8329 VSS.n8333 4.5005
R4307 VSS.n8330 VSS.n8334 4.5005
R4308 VSS.n8331 VSS.n8335 4.57324
R4309 VSS.n8327 VSS.n8325 0.147342
R4310 VSS.n8328 VSS.n8329 0.0732424
R4311 VSS.n8329 VSS.n8330 0.147342
R4312 VSS.n8332 VSS.n8336 0.0721009
R4313 VSS.n8337 VSS.n8333 4.5005
R4314 VSS.n8338 VSS.n8334 4.5005
R4315 VSS.n8339 VSS.n8335 4.5005
R4316 VSS.n8325 VSS.n8336 4.57442
R4317 VSS.n8332 VSS.n8333 0.147342
R4318 VSS.n8333 VSS.n8334 0.147342
R4319 VSS.n8334 VSS.n8335 0.147342
R4320 VSS.n8336 VSS.n8337 2.39784
R4321 VSS.n8337 VSS.n8338 0.147342
R4322 VSS.n8338 VSS.n8339 0.147342
R4323 VSS.n8339 VSS.t55 3.13212
R4324 VSS.n8312 VSS.n8317 4.5005
R4325 VSS.n8314 VSS.n8318 4.5005
R4326 VSS.n8315 VSS.n8319 4.5005
R4327 VSS.n8316 VSS.n8320 4.57324
R4328 VSS.n8312 VSS.n8310 0.147342
R4329 VSS.n8313 VSS.n8314 0.0732424
R4330 VSS.n8314 VSS.n8315 0.147342
R4331 VSS.n8317 VSS.n8321 0.0721009
R4332 VSS.n8322 VSS.n8318 4.5005
R4333 VSS.n8323 VSS.n8319 4.5005
R4334 VSS.n8324 VSS.n8320 4.5005
R4335 VSS.n8310 VSS.n8321 4.57442
R4336 VSS.n8317 VSS.n8318 0.147342
R4337 VSS.n8318 VSS.n8319 0.147342
R4338 VSS.n8319 VSS.n8320 0.147342
R4339 VSS.n8321 VSS.n8322 2.39784
R4340 VSS.n8322 VSS.n8323 0.147342
R4341 VSS.n8323 VSS.n8324 0.147342
R4342 VSS.n8324 VSS.t206 3.13212
R4343 VSS.n8297 VSS.n8302 4.5005
R4344 VSS.n8299 VSS.n8303 4.5005
R4345 VSS.n8300 VSS.n8304 4.5005
R4346 VSS.n8301 VSS.n8305 4.57324
R4347 VSS.n8297 VSS.n8295 0.147342
R4348 VSS.n8298 VSS.n8299 0.0732424
R4349 VSS.n8299 VSS.n8300 0.147342
R4350 VSS.n8302 VSS.n8306 0.0721009
R4351 VSS.n8307 VSS.n8303 4.5005
R4352 VSS.n8308 VSS.n8304 4.5005
R4353 VSS.n8309 VSS.n8305 4.5005
R4354 VSS.n8295 VSS.n8306 4.57442
R4355 VSS.n8302 VSS.n8303 0.147342
R4356 VSS.n8303 VSS.n8304 0.147342
R4357 VSS.n8304 VSS.n8305 0.147342
R4358 VSS.n8306 VSS.n8307 2.39784
R4359 VSS.n8307 VSS.n8308 0.147342
R4360 VSS.n8308 VSS.n8309 0.147342
R4361 VSS.n8309 VSS.t390 3.13212
R4362 VSS.n8287 VSS.n8282 4.5005
R4363 VSS.n8288 VSS.n8284 4.5005
R4364 VSS.n8289 VSS.n8285 4.5005
R4365 VSS.n8290 VSS.n8286 4.57324
R4366 VSS.n8280 VSS.n8282 0.147342
R4367 VSS.n8283 VSS.n8284 0.0732424
R4368 VSS.n8284 VSS.n8285 0.147342
R4369 VSS.n8291 VSS.n8287 0.0722544
R4370 VSS.n8292 VSS.n8288 4.5005
R4371 VSS.n8293 VSS.n8289 4.5005
R4372 VSS.n8294 VSS.n8290 4.5005
R4373 VSS.n8291 VSS.n8280 4.57426
R4374 VSS.n8287 VSS.n8288 0.147342
R4375 VSS.n8288 VSS.n8289 0.147342
R4376 VSS.n8289 VSS.n8290 0.147342
R4377 VSS.n8292 VSS.n8291 2.37296
R4378 VSS.n8293 VSS.n8292 0.127318
R4379 VSS.n8294 VSS.n8293 0.127318
R4380 VSS.t41 VSS.n8294 2.73618
R4381 VSS.n8267 VSS.n8272 4.5005
R4382 VSS.n8269 VSS.n8273 4.5005
R4383 VSS.n8270 VSS.n8274 4.5005
R4384 VSS.n8271 VSS.n8275 4.57324
R4385 VSS.n8267 VSS.n8265 0.147342
R4386 VSS.n8268 VSS.n8269 0.0732424
R4387 VSS.n8269 VSS.n8270 0.147342
R4388 VSS.n8272 VSS.n8276 0.0721009
R4389 VSS.n8277 VSS.n8273 4.5005
R4390 VSS.n8278 VSS.n8274 4.5005
R4391 VSS.n8279 VSS.n8275 4.5005
R4392 VSS.n8265 VSS.n8276 4.57442
R4393 VSS.n8272 VSS.n8273 0.147342
R4394 VSS.n8273 VSS.n8274 0.147342
R4395 VSS.n8274 VSS.n8275 0.147342
R4396 VSS.n8276 VSS.n8277 2.39784
R4397 VSS.n8277 VSS.n8278 0.147342
R4398 VSS.n8278 VSS.n8279 0.147342
R4399 VSS.n8279 VSS.t556 3.13212
R4400 VSS.n8252 VSS.n8257 4.5005
R4401 VSS.n8254 VSS.n8258 4.5005
R4402 VSS.n8255 VSS.n8259 4.5005
R4403 VSS.n8256 VSS.n8260 4.57324
R4404 VSS.n8252 VSS.n8250 0.147342
R4405 VSS.n8253 VSS.n8254 0.0732424
R4406 VSS.n8254 VSS.n8255 0.147342
R4407 VSS.n8257 VSS.n8261 0.0721009
R4408 VSS.n8262 VSS.n8258 4.5005
R4409 VSS.n8263 VSS.n8259 4.5005
R4410 VSS.n8264 VSS.n8260 4.5005
R4411 VSS.n8250 VSS.n8261 4.57442
R4412 VSS.n8257 VSS.n8258 0.147342
R4413 VSS.n8258 VSS.n8259 0.147342
R4414 VSS.n8259 VSS.n8260 0.147342
R4415 VSS.n8261 VSS.n8262 2.39784
R4416 VSS.n8262 VSS.n8263 0.147342
R4417 VSS.n8263 VSS.n8264 0.147342
R4418 VSS.n8264 VSS.t451 3.13212
R4419 VSS.n8237 VSS.n8242 4.5005
R4420 VSS.n8239 VSS.n8243 4.5005
R4421 VSS.n8240 VSS.n8244 4.5005
R4422 VSS.n8241 VSS.n8245 4.57324
R4423 VSS.n8237 VSS.n8235 0.147342
R4424 VSS.n8238 VSS.n8239 0.0732424
R4425 VSS.n8239 VSS.n8240 0.147342
R4426 VSS.n8242 VSS.n8246 0.0721009
R4427 VSS.n8247 VSS.n8243 4.5005
R4428 VSS.n8248 VSS.n8244 4.5005
R4429 VSS.n8249 VSS.n8245 4.5005
R4430 VSS.n8235 VSS.n8246 4.57442
R4431 VSS.n8242 VSS.n8243 0.147342
R4432 VSS.n8243 VSS.n8244 0.147342
R4433 VSS.n8244 VSS.n8245 0.147342
R4434 VSS.n8246 VSS.n8247 2.39784
R4435 VSS.n8247 VSS.n8248 0.147342
R4436 VSS.n8248 VSS.n8249 0.147342
R4437 VSS.n8249 VSS.t585 3.13212
R4438 VSS.n8222 VSS.n8227 4.5005
R4439 VSS.n8224 VSS.n8228 4.5005
R4440 VSS.n8225 VSS.n8229 4.5005
R4441 VSS.n8226 VSS.n8230 4.57324
R4442 VSS.n8222 VSS.n8220 0.147342
R4443 VSS.n8223 VSS.n8224 0.0732424
R4444 VSS.n8224 VSS.n8225 0.147342
R4445 VSS.n8227 VSS.n8231 0.0721009
R4446 VSS.n8232 VSS.n8228 4.5005
R4447 VSS.n8233 VSS.n8229 4.5005
R4448 VSS.n8234 VSS.n8230 4.5005
R4449 VSS.n8220 VSS.n8231 4.57442
R4450 VSS.n8227 VSS.n8228 0.147342
R4451 VSS.n8228 VSS.n8229 0.147342
R4452 VSS.n8229 VSS.n8230 0.147342
R4453 VSS.n8231 VSS.n8232 2.39784
R4454 VSS.n8232 VSS.n8233 0.147342
R4455 VSS.n8233 VSS.n8234 0.147342
R4456 VSS.n8234 VSS.t489 3.13212
R4457 VSS.n8207 VSS.n8212 4.5005
R4458 VSS.n8209 VSS.n8213 4.5005
R4459 VSS.n8210 VSS.n8214 4.5005
R4460 VSS.n8211 VSS.n8215 4.57324
R4461 VSS.n8207 VSS.n8205 0.147342
R4462 VSS.n8208 VSS.n8209 0.0732424
R4463 VSS.n8209 VSS.n8210 0.147342
R4464 VSS.n8212 VSS.n8216 0.0721009
R4465 VSS.n8217 VSS.n8213 4.5005
R4466 VSS.n8218 VSS.n8214 4.5005
R4467 VSS.n8219 VSS.n8215 4.5005
R4468 VSS.n8205 VSS.n8216 4.57442
R4469 VSS.n8212 VSS.n8213 0.147342
R4470 VSS.n8213 VSS.n8214 0.147342
R4471 VSS.n8214 VSS.n8215 0.147342
R4472 VSS.n8216 VSS.n8217 2.39784
R4473 VSS.n8217 VSS.n8218 0.147342
R4474 VSS.n8218 VSS.n8219 0.147342
R4475 VSS.n8219 VSS.t273 3.13212
R4476 VSS.n8192 VSS.n8197 4.5005
R4477 VSS.n8194 VSS.n8198 4.5005
R4478 VSS.n8195 VSS.n8199 4.5005
R4479 VSS.n8196 VSS.n8200 4.57324
R4480 VSS.n8192 VSS.n8190 0.147342
R4481 VSS.n8193 VSS.n8194 0.0732424
R4482 VSS.n8194 VSS.n8195 0.147342
R4483 VSS.n8197 VSS.n8201 0.0721009
R4484 VSS.n8202 VSS.n8198 4.5005
R4485 VSS.n8203 VSS.n8199 4.5005
R4486 VSS.n8204 VSS.n8200 4.5005
R4487 VSS.n8190 VSS.n8201 4.57442
R4488 VSS.n8197 VSS.n8198 0.147342
R4489 VSS.n8198 VSS.n8199 0.147342
R4490 VSS.n8199 VSS.n8200 0.147342
R4491 VSS.n8201 VSS.n8202 2.39784
R4492 VSS.n8202 VSS.n8203 0.147342
R4493 VSS.n8203 VSS.n8204 0.147342
R4494 VSS.n8204 VSS.t448 3.13212
R4495 VSS.n8182 VSS.n8177 4.5005
R4496 VSS.n8183 VSS.n8179 4.5005
R4497 VSS.n8184 VSS.n8180 4.5005
R4498 VSS.n8185 VSS.n8181 4.57324
R4499 VSS.n8175 VSS.n8177 0.147342
R4500 VSS.n8178 VSS.n8179 0.0732424
R4501 VSS.n8179 VSS.n8180 0.147342
R4502 VSS.n8186 VSS.n8182 0.0722544
R4503 VSS.n8187 VSS.n8183 4.5005
R4504 VSS.n8188 VSS.n8184 4.5005
R4505 VSS.n8189 VSS.n8185 4.5005
R4506 VSS.n8186 VSS.n8175 4.57426
R4507 VSS.n8182 VSS.n8183 0.147342
R4508 VSS.n8183 VSS.n8184 0.147342
R4509 VSS.n8184 VSS.n8185 0.147342
R4510 VSS.n8187 VSS.n8186 2.37296
R4511 VSS.n8188 VSS.n8187 0.127318
R4512 VSS.n8189 VSS.n8188 0.127318
R4513 VSS.t41 VSS.n8189 2.73618
R4514 VSS.n8162 VSS.n8167 4.5005
R4515 VSS.n8164 VSS.n8168 4.5005
R4516 VSS.n8165 VSS.n8169 4.5005
R4517 VSS.n8166 VSS.n8170 4.57324
R4518 VSS.n8162 VSS.n8160 0.147342
R4519 VSS.n8163 VSS.n8164 0.0732424
R4520 VSS.n8164 VSS.n8165 0.147342
R4521 VSS.n8167 VSS.n8171 0.0721009
R4522 VSS.n8172 VSS.n8168 4.5005
R4523 VSS.n8173 VSS.n8169 4.5005
R4524 VSS.n8174 VSS.n8170 4.5005
R4525 VSS.n8160 VSS.n8171 4.57442
R4526 VSS.n8167 VSS.n8168 0.147342
R4527 VSS.n8168 VSS.n8169 0.147342
R4528 VSS.n8169 VSS.n8170 0.147342
R4529 VSS.n8171 VSS.n8172 2.39784
R4530 VSS.n8172 VSS.n8173 0.147342
R4531 VSS.n8173 VSS.n8174 0.147342
R4532 VSS.n8174 VSS.t616 3.13212
R4533 VSS.n8147 VSS.n8152 4.5005
R4534 VSS.n8149 VSS.n8153 4.5005
R4535 VSS.n8150 VSS.n8154 4.5005
R4536 VSS.n8151 VSS.n8155 4.57324
R4537 VSS.n8147 VSS.n8145 0.147342
R4538 VSS.n8148 VSS.n8149 0.0732424
R4539 VSS.n8149 VSS.n8150 0.147342
R4540 VSS.n8152 VSS.n8156 0.0721009
R4541 VSS.n8157 VSS.n8153 4.5005
R4542 VSS.n8158 VSS.n8154 4.5005
R4543 VSS.n8159 VSS.n8155 4.5005
R4544 VSS.n8145 VSS.n8156 4.57442
R4545 VSS.n8152 VSS.n8153 0.147342
R4546 VSS.n8153 VSS.n8154 0.147342
R4547 VSS.n8154 VSS.n8155 0.147342
R4548 VSS.n8156 VSS.n8157 2.39784
R4549 VSS.n8157 VSS.n8158 0.147342
R4550 VSS.n8158 VSS.n8159 0.147342
R4551 VSS.n8159 VSS.t522 3.13212
R4552 VSS.n8132 VSS.n8137 4.5005
R4553 VSS.n8134 VSS.n8138 4.5005
R4554 VSS.n8135 VSS.n8139 4.5005
R4555 VSS.n8136 VSS.n8140 4.57324
R4556 VSS.n8132 VSS.n8130 0.147342
R4557 VSS.n8133 VSS.n8134 0.0732424
R4558 VSS.n8134 VSS.n8135 0.147342
R4559 VSS.n8137 VSS.n8141 0.0721009
R4560 VSS.n8142 VSS.n8138 4.5005
R4561 VSS.n8143 VSS.n8139 4.5005
R4562 VSS.n8144 VSS.n8140 4.5005
R4563 VSS.n8130 VSS.n8141 4.57442
R4564 VSS.n8137 VSS.n8138 0.147342
R4565 VSS.n8138 VSS.n8139 0.147342
R4566 VSS.n8139 VSS.n8140 0.147342
R4567 VSS.n8141 VSS.n8142 2.39784
R4568 VSS.n8142 VSS.n8143 0.147342
R4569 VSS.n8143 VSS.n8144 0.147342
R4570 VSS.n8144 VSS.t527 3.13212
R4571 VSS.n8122 VSS.n8117 4.5005
R4572 VSS.n8123 VSS.n8119 4.5005
R4573 VSS.n8124 VSS.n8120 4.5005
R4574 VSS.n8125 VSS.n8121 4.57324
R4575 VSS.n8115 VSS.n8117 0.147342
R4576 VSS.n8118 VSS.n8119 0.0732424
R4577 VSS.n8119 VSS.n8120 0.147342
R4578 VSS.n8126 VSS.n8122 0.0722544
R4579 VSS.n8127 VSS.n8123 4.5005
R4580 VSS.n8128 VSS.n8124 4.5005
R4581 VSS.n8129 VSS.n8125 4.5005
R4582 VSS.n8126 VSS.n8115 4.57426
R4583 VSS.n8122 VSS.n8123 0.147342
R4584 VSS.n8123 VSS.n8124 0.147342
R4585 VSS.n8124 VSS.n8125 0.147342
R4586 VSS.n8127 VSS.n8126 2.37296
R4587 VSS.n8128 VSS.n8127 0.127318
R4588 VSS.n8129 VSS.n8128 0.127318
R4589 VSS.t41 VSS.n8129 2.73618
R4590 VSS.n8102 VSS.n8107 4.5005
R4591 VSS.n8104 VSS.n8108 4.5005
R4592 VSS.n8105 VSS.n8109 4.5005
R4593 VSS.n8106 VSS.n8110 4.57324
R4594 VSS.n8102 VSS.n8100 0.147342
R4595 VSS.n8103 VSS.n8104 0.0732424
R4596 VSS.n8104 VSS.n8105 0.147342
R4597 VSS.n8107 VSS.n8111 0.0721009
R4598 VSS.n8112 VSS.n8108 4.5005
R4599 VSS.n8113 VSS.n8109 4.5005
R4600 VSS.n8114 VSS.n8110 4.5005
R4601 VSS.n8100 VSS.n8111 4.57442
R4602 VSS.n8107 VSS.n8108 0.147342
R4603 VSS.n8108 VSS.n8109 0.147342
R4604 VSS.n8109 VSS.n8110 0.147342
R4605 VSS.n8111 VSS.n8112 2.39784
R4606 VSS.n8112 VSS.n8113 0.147342
R4607 VSS.n8113 VSS.n8114 0.147342
R4608 VSS.n8114 VSS.t110 3.13212
R4609 VSS.n8087 VSS.n8092 4.5005
R4610 VSS.n8089 VSS.n8093 4.5005
R4611 VSS.n8090 VSS.n8094 4.5005
R4612 VSS.n8091 VSS.n8095 4.57324
R4613 VSS.n8087 VSS.n8085 0.147342
R4614 VSS.n8088 VSS.n8089 0.0732424
R4615 VSS.n8089 VSS.n8090 0.147342
R4616 VSS.n8092 VSS.n8096 0.0721009
R4617 VSS.n8097 VSS.n8093 4.5005
R4618 VSS.n8098 VSS.n8094 4.5005
R4619 VSS.n8099 VSS.n8095 4.5005
R4620 VSS.n8085 VSS.n8096 4.57442
R4621 VSS.n8092 VSS.n8093 0.147342
R4622 VSS.n8093 VSS.n8094 0.147342
R4623 VSS.n8094 VSS.n8095 0.147342
R4624 VSS.n8096 VSS.n8097 2.39784
R4625 VSS.n8097 VSS.n8098 0.147342
R4626 VSS.n8098 VSS.n8099 0.147342
R4627 VSS.n8099 VSS.t499 3.13212
R4628 VSS.n8072 VSS.n8077 4.5005
R4629 VSS.n8074 VSS.n8078 4.5005
R4630 VSS.n8075 VSS.n8079 4.5005
R4631 VSS.n8076 VSS.n8080 4.57324
R4632 VSS.n8072 VSS.n8070 0.147342
R4633 VSS.n8073 VSS.n8074 0.0732424
R4634 VSS.n8074 VSS.n8075 0.147342
R4635 VSS.n8077 VSS.n8081 0.0721009
R4636 VSS.n8082 VSS.n8078 4.5005
R4637 VSS.n8083 VSS.n8079 4.5005
R4638 VSS.n8084 VSS.n8080 4.5005
R4639 VSS.n8070 VSS.n8081 4.57442
R4640 VSS.n8077 VSS.n8078 0.147342
R4641 VSS.n8078 VSS.n8079 0.147342
R4642 VSS.n8079 VSS.n8080 0.147342
R4643 VSS.n8081 VSS.n8082 2.39784
R4644 VSS.n8082 VSS.n8083 0.147342
R4645 VSS.n8083 VSS.n8084 0.147342
R4646 VSS.n8084 VSS.t614 3.13212
R4647 VSS.n8057 VSS.n8062 4.5005
R4648 VSS.n8059 VSS.n8063 4.5005
R4649 VSS.n8060 VSS.n8064 4.5005
R4650 VSS.n8061 VSS.n8065 4.57324
R4651 VSS.n8057 VSS.n8055 0.147342
R4652 VSS.n8058 VSS.n8059 0.0732424
R4653 VSS.n8059 VSS.n8060 0.147342
R4654 VSS.n8062 VSS.n8066 0.0721009
R4655 VSS.n8067 VSS.n8063 4.5005
R4656 VSS.n8068 VSS.n8064 4.5005
R4657 VSS.n8069 VSS.n8065 4.5005
R4658 VSS.n8055 VSS.n8066 4.57442
R4659 VSS.n8062 VSS.n8063 0.147342
R4660 VSS.n8063 VSS.n8064 0.147342
R4661 VSS.n8064 VSS.n8065 0.147342
R4662 VSS.n8066 VSS.n8067 2.39784
R4663 VSS.n8067 VSS.n8068 0.147342
R4664 VSS.n8068 VSS.n8069 0.147342
R4665 VSS.n8069 VSS.t604 3.13212
R4666 VSS.n8047 VSS.n8042 4.5005
R4667 VSS.n8048 VSS.n8044 4.5005
R4668 VSS.n8049 VSS.n8045 4.5005
R4669 VSS.n8050 VSS.n8046 4.57324
R4670 VSS.n8040 VSS.n8042 0.147342
R4671 VSS.n8043 VSS.n8044 0.0732424
R4672 VSS.n8044 VSS.n8045 0.147342
R4673 VSS.n8051 VSS.n8047 0.0722544
R4674 VSS.n8052 VSS.n8048 4.5005
R4675 VSS.n8053 VSS.n8049 4.5005
R4676 VSS.n8054 VSS.n8050 4.5005
R4677 VSS.n8051 VSS.n8040 4.57426
R4678 VSS.n8047 VSS.n8048 0.147342
R4679 VSS.n8048 VSS.n8049 0.147342
R4680 VSS.n8049 VSS.n8050 0.147342
R4681 VSS.n8052 VSS.n8051 2.37296
R4682 VSS.n8053 VSS.n8052 0.127318
R4683 VSS.n8054 VSS.n8053 0.127318
R4684 VSS.t41 VSS.n8054 2.73618
R4685 VSS.n8027 VSS.n8032 4.5005
R4686 VSS.n8029 VSS.n8033 4.5005
R4687 VSS.n8030 VSS.n8034 4.5005
R4688 VSS.n8031 VSS.n8035 4.57324
R4689 VSS.n8027 VSS.n8025 0.147342
R4690 VSS.n8028 VSS.n8029 0.0732424
R4691 VSS.n8029 VSS.n8030 0.147342
R4692 VSS.n8032 VSS.n8036 0.0721009
R4693 VSS.n8037 VSS.n8033 4.5005
R4694 VSS.n8038 VSS.n8034 4.5005
R4695 VSS.n8039 VSS.n8035 4.5005
R4696 VSS.n8025 VSS.n8036 4.57442
R4697 VSS.n8032 VSS.n8033 0.147342
R4698 VSS.n8033 VSS.n8034 0.147342
R4699 VSS.n8034 VSS.n8035 0.147342
R4700 VSS.n8036 VSS.n8037 2.39784
R4701 VSS.n8037 VSS.n8038 0.147342
R4702 VSS.n8038 VSS.n8039 0.147342
R4703 VSS.n8039 VSS.t578 3.13212
R4704 VSS.n8012 VSS.n8017 4.5005
R4705 VSS.n8014 VSS.n8018 4.5005
R4706 VSS.n8015 VSS.n8019 4.5005
R4707 VSS.n8016 VSS.n8020 4.57324
R4708 VSS.n8012 VSS.n8010 0.147342
R4709 VSS.n8013 VSS.n8014 0.0732424
R4710 VSS.n8014 VSS.n8015 0.147342
R4711 VSS.n8017 VSS.n8021 0.0721009
R4712 VSS.n8022 VSS.n8018 4.5005
R4713 VSS.n8023 VSS.n8019 4.5005
R4714 VSS.n8024 VSS.n8020 4.5005
R4715 VSS.n8010 VSS.n8021 4.57442
R4716 VSS.n8017 VSS.n8018 0.147342
R4717 VSS.n8018 VSS.n8019 0.147342
R4718 VSS.n8019 VSS.n8020 0.147342
R4719 VSS.n8021 VSS.n8022 2.39784
R4720 VSS.n8022 VSS.n8023 0.147342
R4721 VSS.n8023 VSS.n8024 0.147342
R4722 VSS.n8024 VSS.t202 3.13212
R4723 VSS.n7997 VSS.n8002 4.5005
R4724 VSS.n7999 VSS.n8003 4.5005
R4725 VSS.n8000 VSS.n8004 4.5005
R4726 VSS.n8001 VSS.n8005 4.57324
R4727 VSS.n7997 VSS.n7995 0.147342
R4728 VSS.n7998 VSS.n7999 0.0732424
R4729 VSS.n7999 VSS.n8000 0.147342
R4730 VSS.n8002 VSS.n8006 0.0721009
R4731 VSS.n8007 VSS.n8003 4.5005
R4732 VSS.n8008 VSS.n8004 4.5005
R4733 VSS.n8009 VSS.n8005 4.5005
R4734 VSS.n7995 VSS.n8006 4.57442
R4735 VSS.n8002 VSS.n8003 0.147342
R4736 VSS.n8003 VSS.n8004 0.147342
R4737 VSS.n8004 VSS.n8005 0.147342
R4738 VSS.n8006 VSS.n8007 2.39784
R4739 VSS.n8007 VSS.n8008 0.147342
R4740 VSS.n8008 VSS.n8009 0.147342
R4741 VSS.n8009 VSS.t409 3.13212
R4742 VSS.n7987 VSS.n7982 4.5005
R4743 VSS.n7988 VSS.n7984 4.5005
R4744 VSS.n7989 VSS.n7985 4.5005
R4745 VSS.n7990 VSS.n7986 4.57324
R4746 VSS.n7980 VSS.n7982 0.147342
R4747 VSS.n7983 VSS.n7984 0.0732424
R4748 VSS.n7984 VSS.n7985 0.147342
R4749 VSS.n7991 VSS.n7987 0.0722544
R4750 VSS.n7992 VSS.n7988 4.5005
R4751 VSS.n7993 VSS.n7989 4.5005
R4752 VSS.n7994 VSS.n7990 4.5005
R4753 VSS.n7991 VSS.n7980 4.57426
R4754 VSS.n7987 VSS.n7988 0.147342
R4755 VSS.n7988 VSS.n7989 0.147342
R4756 VSS.n7989 VSS.n7990 0.147342
R4757 VSS.n7992 VSS.n7991 2.37296
R4758 VSS.n7993 VSS.n7992 0.127318
R4759 VSS.n7994 VSS.n7993 0.127318
R4760 VSS.t41 VSS.n7994 2.73618
R4761 VSS.n7967 VSS.n7972 4.5005
R4762 VSS.n7969 VSS.n7973 4.5005
R4763 VSS.n7970 VSS.n7974 4.5005
R4764 VSS.n7971 VSS.n7975 4.57324
R4765 VSS.n7967 VSS.n7965 0.147342
R4766 VSS.n7968 VSS.n7969 0.0732424
R4767 VSS.n7969 VSS.n7970 0.147342
R4768 VSS.n7972 VSS.n7976 0.0721009
R4769 VSS.n7977 VSS.n7973 4.5005
R4770 VSS.n7978 VSS.n7974 4.5005
R4771 VSS.n7979 VSS.n7975 4.5005
R4772 VSS.n7965 VSS.n7976 4.57442
R4773 VSS.n7972 VSS.n7973 0.147342
R4774 VSS.n7973 VSS.n7974 0.147342
R4775 VSS.n7974 VSS.n7975 0.147342
R4776 VSS.n7976 VSS.n7977 2.39784
R4777 VSS.n7977 VSS.n7978 0.147342
R4778 VSS.n7978 VSS.n7979 0.147342
R4779 VSS.n7979 VSS.t540 3.13212
R4780 VSS.n7952 VSS.n7957 4.5005
R4781 VSS.n7954 VSS.n7958 4.5005
R4782 VSS.n7955 VSS.n7959 4.5005
R4783 VSS.n7956 VSS.n7960 4.57324
R4784 VSS.n7952 VSS.n7950 0.147342
R4785 VSS.n7953 VSS.n7954 0.0732424
R4786 VSS.n7954 VSS.n7955 0.147342
R4787 VSS.n7957 VSS.n7961 0.0721009
R4788 VSS.n7962 VSS.n7958 4.5005
R4789 VSS.n7963 VSS.n7959 4.5005
R4790 VSS.n7964 VSS.n7960 4.5005
R4791 VSS.n7950 VSS.n7961 4.57442
R4792 VSS.n7957 VSS.n7958 0.147342
R4793 VSS.n7958 VSS.n7959 0.147342
R4794 VSS.n7959 VSS.n7960 0.147342
R4795 VSS.n7961 VSS.n7962 2.39784
R4796 VSS.n7962 VSS.n7963 0.147342
R4797 VSS.n7963 VSS.n7964 0.147342
R4798 VSS.n7964 VSS.t453 3.13212
R4799 VSS.n7937 VSS.n7942 4.5005
R4800 VSS.n7939 VSS.n7943 4.5005
R4801 VSS.n7940 VSS.n7944 4.5005
R4802 VSS.n7941 VSS.n7945 4.57324
R4803 VSS.n7937 VSS.n7935 0.147342
R4804 VSS.n7938 VSS.n7939 0.0732424
R4805 VSS.n7939 VSS.n7940 0.147342
R4806 VSS.n7942 VSS.n7946 0.0721009
R4807 VSS.n7947 VSS.n7943 4.5005
R4808 VSS.n7948 VSS.n7944 4.5005
R4809 VSS.n7949 VSS.n7945 4.5005
R4810 VSS.n7935 VSS.n7946 4.57442
R4811 VSS.n7942 VSS.n7943 0.147342
R4812 VSS.n7943 VSS.n7944 0.147342
R4813 VSS.n7944 VSS.n7945 0.147342
R4814 VSS.n7946 VSS.n7947 2.39784
R4815 VSS.n7947 VSS.n7948 0.147342
R4816 VSS.n7948 VSS.n7949 0.147342
R4817 VSS.n7949 VSS.t591 3.13212
R4818 VSS.n7922 VSS.n7927 4.5005
R4819 VSS.n7924 VSS.n7928 4.5005
R4820 VSS.n7925 VSS.n7929 4.5005
R4821 VSS.n7926 VSS.n7930 4.57324
R4822 VSS.n7922 VSS.n7920 0.147342
R4823 VSS.n7923 VSS.n7924 0.0732424
R4824 VSS.n7924 VSS.n7925 0.147342
R4825 VSS.n7927 VSS.n7931 0.0721009
R4826 VSS.n7932 VSS.n7928 4.5005
R4827 VSS.n7933 VSS.n7929 4.5005
R4828 VSS.n7934 VSS.n7930 4.5005
R4829 VSS.n7920 VSS.n7931 4.57442
R4830 VSS.n7927 VSS.n7928 0.147342
R4831 VSS.n7928 VSS.n7929 0.147342
R4832 VSS.n7929 VSS.n7930 0.147342
R4833 VSS.n7931 VSS.n7932 2.39784
R4834 VSS.n7932 VSS.n7933 0.147342
R4835 VSS.n7933 VSS.n7934 0.147342
R4836 VSS.n7934 VSS.t67 3.13212
R4837 VSS.n7907 VSS.n7912 4.5005
R4838 VSS.n7909 VSS.n7913 4.5005
R4839 VSS.n7910 VSS.n7914 4.5005
R4840 VSS.n7911 VSS.n7915 4.57324
R4841 VSS.n7907 VSS.n7905 0.147342
R4842 VSS.n7908 VSS.n7909 0.0732424
R4843 VSS.n7909 VSS.n7910 0.147342
R4844 VSS.n7912 VSS.n7916 0.0721009
R4845 VSS.n7917 VSS.n7913 4.5005
R4846 VSS.n7918 VSS.n7914 4.5005
R4847 VSS.n7919 VSS.n7915 4.5005
R4848 VSS.n7905 VSS.n7916 4.57442
R4849 VSS.n7912 VSS.n7913 0.147342
R4850 VSS.n7913 VSS.n7914 0.147342
R4851 VSS.n7914 VSS.n7915 0.147342
R4852 VSS.n7916 VSS.n7917 2.39784
R4853 VSS.n7917 VSS.n7918 0.147342
R4854 VSS.n7918 VSS.n7919 0.147342
R4855 VSS.n7919 VSS.t274 3.13212
R4856 VSS.n7892 VSS.n7897 4.5005
R4857 VSS.n7894 VSS.n7898 4.5005
R4858 VSS.n7895 VSS.n7899 4.5005
R4859 VSS.n7896 VSS.n7900 4.57324
R4860 VSS.n7892 VSS.n7890 0.147342
R4861 VSS.n7893 VSS.n7894 0.0732424
R4862 VSS.n7894 VSS.n7895 0.147342
R4863 VSS.n7897 VSS.n7901 0.0721009
R4864 VSS.n7902 VSS.n7898 4.5005
R4865 VSS.n7903 VSS.n7899 4.5005
R4866 VSS.n7904 VSS.n7900 4.5005
R4867 VSS.n7890 VSS.n7901 4.57442
R4868 VSS.n7897 VSS.n7898 0.147342
R4869 VSS.n7898 VSS.n7899 0.147342
R4870 VSS.n7899 VSS.n7900 0.147342
R4871 VSS.n7901 VSS.n7902 2.39784
R4872 VSS.n7902 VSS.n7903 0.147342
R4873 VSS.n7903 VSS.n7904 0.147342
R4874 VSS.n7904 VSS.t447 3.13212
R4875 VSS.n7882 VSS.n7877 4.5005
R4876 VSS.n7883 VSS.n7879 4.5005
R4877 VSS.n7884 VSS.n7880 4.5005
R4878 VSS.n7885 VSS.n7881 4.57324
R4879 VSS.n7875 VSS.n7877 0.147342
R4880 VSS.n7878 VSS.n7879 0.0732424
R4881 VSS.n7879 VSS.n7880 0.147342
R4882 VSS.n7886 VSS.n7882 0.0722544
R4883 VSS.n7887 VSS.n7883 4.5005
R4884 VSS.n7888 VSS.n7884 4.5005
R4885 VSS.n7889 VSS.n7885 4.5005
R4886 VSS.n7886 VSS.n7875 4.57426
R4887 VSS.n7882 VSS.n7883 0.147342
R4888 VSS.n7883 VSS.n7884 0.147342
R4889 VSS.n7884 VSS.n7885 0.147342
R4890 VSS.n7887 VSS.n7886 2.37296
R4891 VSS.n7888 VSS.n7887 0.127318
R4892 VSS.n7889 VSS.n7888 0.127318
R4893 VSS.t41 VSS.n7889 2.73618
R4894 VSS.n7862 VSS.n7867 4.5005
R4895 VSS.n7864 VSS.n7868 4.5005
R4896 VSS.n7865 VSS.n7869 4.5005
R4897 VSS.n7866 VSS.n7870 4.57324
R4898 VSS.n7862 VSS.n7860 0.147342
R4899 VSS.n7863 VSS.n7864 0.0732424
R4900 VSS.n7864 VSS.n7865 0.147342
R4901 VSS.n7867 VSS.n7871 0.0721009
R4902 VSS.n7872 VSS.n7868 4.5005
R4903 VSS.n7873 VSS.n7869 4.5005
R4904 VSS.n7874 VSS.n7870 4.5005
R4905 VSS.n7860 VSS.n7871 4.57442
R4906 VSS.n7867 VSS.n7868 0.147342
R4907 VSS.n7868 VSS.n7869 0.147342
R4908 VSS.n7869 VSS.n7870 0.147342
R4909 VSS.n7871 VSS.n7872 2.39784
R4910 VSS.n7872 VSS.n7873 0.147342
R4911 VSS.n7873 VSS.n7874 0.147342
R4912 VSS.n7874 VSS.t612 3.13212
R4913 VSS.n7847 VSS.n7852 4.5005
R4914 VSS.n7849 VSS.n7853 4.5005
R4915 VSS.n7850 VSS.n7854 4.5005
R4916 VSS.n7851 VSS.n7855 4.57324
R4917 VSS.n7847 VSS.n7845 0.147342
R4918 VSS.n7848 VSS.n7849 0.0732424
R4919 VSS.n7849 VSS.n7850 0.147342
R4920 VSS.n7852 VSS.n7856 0.0721009
R4921 VSS.n7857 VSS.n7853 4.5005
R4922 VSS.n7858 VSS.n7854 4.5005
R4923 VSS.n7859 VSS.n7855 4.5005
R4924 VSS.n7845 VSS.n7856 4.57442
R4925 VSS.n7852 VSS.n7853 0.147342
R4926 VSS.n7853 VSS.n7854 0.147342
R4927 VSS.n7854 VSS.n7855 0.147342
R4928 VSS.n7856 VSS.n7857 2.39784
R4929 VSS.n7857 VSS.n7858 0.147342
R4930 VSS.n7858 VSS.n7859 0.147342
R4931 VSS.n7859 VSS.t49 3.13212
R4932 VSS.n7832 VSS.n7837 4.5005
R4933 VSS.n7834 VSS.n7838 4.5005
R4934 VSS.n7835 VSS.n7839 4.5005
R4935 VSS.n7836 VSS.n7840 4.57324
R4936 VSS.n7832 VSS.n7830 0.147342
R4937 VSS.n7833 VSS.n7834 0.0732424
R4938 VSS.n7834 VSS.n7835 0.147342
R4939 VSS.n7837 VSS.n7841 0.0721009
R4940 VSS.n7842 VSS.n7838 4.5005
R4941 VSS.n7843 VSS.n7839 4.5005
R4942 VSS.n7844 VSS.n7840 4.5005
R4943 VSS.n7830 VSS.n7841 4.57442
R4944 VSS.n7837 VSS.n7838 0.147342
R4945 VSS.n7838 VSS.n7839 0.147342
R4946 VSS.n7839 VSS.n7840 0.147342
R4947 VSS.n7841 VSS.n7842 2.39784
R4948 VSS.n7842 VSS.n7843 0.147342
R4949 VSS.n7843 VSS.n7844 0.147342
R4950 VSS.n7844 VSS.t533 3.13212
R4951 VSS.n7822 VSS.n7817 4.5005
R4952 VSS.n7823 VSS.n7819 4.5005
R4953 VSS.n7824 VSS.n7820 4.5005
R4954 VSS.n7825 VSS.n7821 4.57324
R4955 VSS.n7815 VSS.n7817 0.147342
R4956 VSS.n7818 VSS.n7819 0.0732424
R4957 VSS.n7819 VSS.n7820 0.147342
R4958 VSS.n7826 VSS.n7822 0.0722544
R4959 VSS.n7827 VSS.n7823 4.5005
R4960 VSS.n7828 VSS.n7824 4.5005
R4961 VSS.n7829 VSS.n7825 4.5005
R4962 VSS.n7826 VSS.n7815 4.57426
R4963 VSS.n7822 VSS.n7823 0.147342
R4964 VSS.n7823 VSS.n7824 0.147342
R4965 VSS.n7824 VSS.n7825 0.147342
R4966 VSS.n7827 VSS.n7826 2.37296
R4967 VSS.n7828 VSS.n7827 0.127318
R4968 VSS.n7829 VSS.n7828 0.127318
R4969 VSS.t41 VSS.n7829 2.73618
R4970 VSS.n7802 VSS.n7807 4.5005
R4971 VSS.n7804 VSS.n7808 4.5005
R4972 VSS.n7805 VSS.n7809 4.5005
R4973 VSS.n7806 VSS.n7810 4.57324
R4974 VSS.n7802 VSS.n7800 0.147342
R4975 VSS.n7803 VSS.n7804 0.0732424
R4976 VSS.n7804 VSS.n7805 0.147342
R4977 VSS.n7807 VSS.n7811 0.0721009
R4978 VSS.n7812 VSS.n7808 4.5005
R4979 VSS.n7813 VSS.n7809 4.5005
R4980 VSS.n7814 VSS.n7810 4.5005
R4981 VSS.n7800 VSS.n7811 4.57442
R4982 VSS.n7807 VSS.n7808 0.147342
R4983 VSS.n7808 VSS.n7809 0.147342
R4984 VSS.n7809 VSS.n7810 0.147342
R4985 VSS.n7811 VSS.n7812 2.39784
R4986 VSS.n7812 VSS.n7813 0.147342
R4987 VSS.n7813 VSS.n7814 0.147342
R4988 VSS.n7814 VSS.t113 3.13212
R4989 VSS.n7787 VSS.n7792 4.5005
R4990 VSS.n7789 VSS.n7793 4.5005
R4991 VSS.n7790 VSS.n7794 4.5005
R4992 VSS.n7791 VSS.n7795 4.57324
R4993 VSS.n7787 VSS.n7785 0.147342
R4994 VSS.n7788 VSS.n7789 0.0732424
R4995 VSS.n7789 VSS.n7790 0.147342
R4996 VSS.n7792 VSS.n7796 0.0721009
R4997 VSS.n7797 VSS.n7793 4.5005
R4998 VSS.n7798 VSS.n7794 4.5005
R4999 VSS.n7799 VSS.n7795 4.5005
R5000 VSS.n7785 VSS.n7796 4.57442
R5001 VSS.n7792 VSS.n7793 0.147342
R5002 VSS.n7793 VSS.n7794 0.147342
R5003 VSS.n7794 VSS.n7795 0.147342
R5004 VSS.n7796 VSS.n7797 2.39784
R5005 VSS.n7797 VSS.n7798 0.147342
R5006 VSS.n7798 VSS.n7799 0.147342
R5007 VSS.n7799 VSS.t501 3.13212
R5008 VSS.n7772 VSS.n7777 4.5005
R5009 VSS.n7774 VSS.n7778 4.5005
R5010 VSS.n7775 VSS.n7779 4.5005
R5011 VSS.n7776 VSS.n7780 4.57324
R5012 VSS.n7772 VSS.n7770 0.147342
R5013 VSS.n7773 VSS.n7774 0.0732424
R5014 VSS.n7774 VSS.n7775 0.147342
R5015 VSS.n7777 VSS.n7781 0.0721009
R5016 VSS.n7782 VSS.n7778 4.5005
R5017 VSS.n7783 VSS.n7779 4.5005
R5018 VSS.n7784 VSS.n7780 4.5005
R5019 VSS.n7770 VSS.n7781 4.57442
R5020 VSS.n7777 VSS.n7778 0.147342
R5021 VSS.n7778 VSS.n7779 0.147342
R5022 VSS.n7779 VSS.n7780 0.147342
R5023 VSS.n7781 VSS.n7782 2.39784
R5024 VSS.n7782 VSS.n7783 0.147342
R5025 VSS.n7783 VSS.n7784 0.147342
R5026 VSS.n7784 VSS.t615 3.13212
R5027 VSS.n7757 VSS.n7762 4.5005
R5028 VSS.n7759 VSS.n7763 4.5005
R5029 VSS.n7760 VSS.n7764 4.5005
R5030 VSS.n7761 VSS.n7765 4.57324
R5031 VSS.n7757 VSS.n7755 0.147342
R5032 VSS.n7758 VSS.n7759 0.0732424
R5033 VSS.n7759 VSS.n7760 0.147342
R5034 VSS.n7762 VSS.n7766 0.0721009
R5035 VSS.n7767 VSS.n7763 4.5005
R5036 VSS.n7768 VSS.n7764 4.5005
R5037 VSS.n7769 VSS.n7765 4.5005
R5038 VSS.n7755 VSS.n7766 4.57442
R5039 VSS.n7762 VSS.n7763 0.147342
R5040 VSS.n7763 VSS.n7764 0.147342
R5041 VSS.n7764 VSS.n7765 0.147342
R5042 VSS.n7766 VSS.n7767 2.39784
R5043 VSS.n7767 VSS.n7768 0.147342
R5044 VSS.n7768 VSS.n7769 0.147342
R5045 VSS.n7769 VSS.t605 3.13212
R5046 VSS.n7747 VSS.n7742 4.5005
R5047 VSS.n7748 VSS.n7744 4.5005
R5048 VSS.n7749 VSS.n7745 4.5005
R5049 VSS.n7750 VSS.n7746 4.57324
R5050 VSS.n7740 VSS.n7742 0.147342
R5051 VSS.n7743 VSS.n7744 0.0732424
R5052 VSS.n7744 VSS.n7745 0.147342
R5053 VSS.n7751 VSS.n7747 0.0722544
R5054 VSS.n7752 VSS.n7748 4.5005
R5055 VSS.n7753 VSS.n7749 4.5005
R5056 VSS.n7754 VSS.n7750 4.5005
R5057 VSS.n7751 VSS.n7740 4.57426
R5058 VSS.n7747 VSS.n7748 0.147342
R5059 VSS.n7748 VSS.n7749 0.147342
R5060 VSS.n7749 VSS.n7750 0.147342
R5061 VSS.n7752 VSS.n7751 2.37296
R5062 VSS.n7753 VSS.n7752 0.127318
R5063 VSS.n7754 VSS.n7753 0.127318
R5064 VSS.t41 VSS.n7754 2.73618
R5065 VSS.n7727 VSS.n7732 4.5005
R5066 VSS.n7729 VSS.n7733 4.5005
R5067 VSS.n7730 VSS.n7734 4.5005
R5068 VSS.n7731 VSS.n7735 4.57324
R5069 VSS.n7727 VSS.n7725 0.147342
R5070 VSS.n7728 VSS.n7729 0.0732424
R5071 VSS.n7729 VSS.n7730 0.147342
R5072 VSS.n7732 VSS.n7736 0.0721009
R5073 VSS.n7737 VSS.n7733 4.5005
R5074 VSS.n7738 VSS.n7734 4.5005
R5075 VSS.n7739 VSS.n7735 4.5005
R5076 VSS.n7725 VSS.n7736 4.57442
R5077 VSS.n7732 VSS.n7733 0.147342
R5078 VSS.n7733 VSS.n7734 0.147342
R5079 VSS.n7734 VSS.n7735 0.147342
R5080 VSS.n7736 VSS.n7737 2.39784
R5081 VSS.n7737 VSS.n7738 0.147342
R5082 VSS.n7738 VSS.n7739 0.147342
R5083 VSS.n7739 VSS.t575 3.13212
R5084 VSS.n7712 VSS.n7717 4.5005
R5085 VSS.n7714 VSS.n7718 4.5005
R5086 VSS.n7715 VSS.n7719 4.5005
R5087 VSS.n7716 VSS.n7720 4.57324
R5088 VSS.n7712 VSS.n7710 0.147342
R5089 VSS.n7713 VSS.n7714 0.0732424
R5090 VSS.n7714 VSS.n7715 0.147342
R5091 VSS.n7717 VSS.n7721 0.0721009
R5092 VSS.n7722 VSS.n7718 4.5005
R5093 VSS.n7723 VSS.n7719 4.5005
R5094 VSS.n7724 VSS.n7720 4.5005
R5095 VSS.n7710 VSS.n7721 4.57442
R5096 VSS.n7717 VSS.n7718 0.147342
R5097 VSS.n7718 VSS.n7719 0.147342
R5098 VSS.n7719 VSS.n7720 0.147342
R5099 VSS.n7721 VSS.n7722 2.39784
R5100 VSS.n7722 VSS.n7723 0.147342
R5101 VSS.n7723 VSS.n7724 0.147342
R5102 VSS.n7724 VSS.t207 3.13212
R5103 VSS.n7697 VSS.n7702 4.5005
R5104 VSS.n7699 VSS.n7703 4.5005
R5105 VSS.n7700 VSS.n7704 4.5005
R5106 VSS.n7701 VSS.n7705 4.57324
R5107 VSS.n7697 VSS.n7695 0.147342
R5108 VSS.n7698 VSS.n7699 0.0732424
R5109 VSS.n7699 VSS.n7700 0.147342
R5110 VSS.n7702 VSS.n7706 0.0721009
R5111 VSS.n7707 VSS.n7703 4.5005
R5112 VSS.n7708 VSS.n7704 4.5005
R5113 VSS.n7709 VSS.n7705 4.5005
R5114 VSS.n7695 VSS.n7706 4.57442
R5115 VSS.n7702 VSS.n7703 0.147342
R5116 VSS.n7703 VSS.n7704 0.147342
R5117 VSS.n7704 VSS.n7705 0.147342
R5118 VSS.n7706 VSS.n7707 2.39784
R5119 VSS.n7707 VSS.n7708 0.147342
R5120 VSS.n7708 VSS.n7709 0.147342
R5121 VSS.n7709 VSS.t411 3.13212
R5122 VSS.n7687 VSS.n7682 4.5005
R5123 VSS.n7688 VSS.n7684 4.5005
R5124 VSS.n7689 VSS.n7685 4.5005
R5125 VSS.n7690 VSS.n7686 4.57324
R5126 VSS.n7680 VSS.n7682 0.147342
R5127 VSS.n7683 VSS.n7684 0.0732424
R5128 VSS.n7684 VSS.n7685 0.147342
R5129 VSS.n7691 VSS.n7687 0.0722544
R5130 VSS.n7692 VSS.n7688 4.5005
R5131 VSS.n7693 VSS.n7689 4.5005
R5132 VSS.n7694 VSS.n7690 4.5005
R5133 VSS.n7691 VSS.n7680 4.57426
R5134 VSS.n7687 VSS.n7688 0.147342
R5135 VSS.n7688 VSS.n7689 0.147342
R5136 VSS.n7689 VSS.n7690 0.147342
R5137 VSS.n7692 VSS.n7691 2.37296
R5138 VSS.n7693 VSS.n7692 0.127318
R5139 VSS.n7694 VSS.n7693 0.127318
R5140 VSS.t41 VSS.n7694 2.73618
R5141 VSS.n7667 VSS.n7672 4.5005
R5142 VSS.n7669 VSS.n7673 4.5005
R5143 VSS.n7670 VSS.n7674 4.5005
R5144 VSS.n7671 VSS.n7675 4.57324
R5145 VSS.n7667 VSS.n7665 0.147342
R5146 VSS.n7668 VSS.n7669 0.0732424
R5147 VSS.n7669 VSS.n7670 0.147342
R5148 VSS.n7672 VSS.n7676 0.0721009
R5149 VSS.n7677 VSS.n7673 4.5005
R5150 VSS.n7678 VSS.n7674 4.5005
R5151 VSS.n7679 VSS.n7675 4.5005
R5152 VSS.n7665 VSS.n7676 4.57442
R5153 VSS.n7672 VSS.n7673 0.147342
R5154 VSS.n7673 VSS.n7674 0.147342
R5155 VSS.n7674 VSS.n7675 0.147342
R5156 VSS.n7676 VSS.n7677 2.39784
R5157 VSS.n7677 VSS.n7678 0.147342
R5158 VSS.n7678 VSS.n7679 0.147342
R5159 VSS.n7679 VSS.t553 3.13212
R5160 VSS.n7652 VSS.n7657 4.5005
R5161 VSS.n7654 VSS.n7658 4.5005
R5162 VSS.n7655 VSS.n7659 4.5005
R5163 VSS.n7656 VSS.n7660 4.57324
R5164 VSS.n7652 VSS.n7650 0.147342
R5165 VSS.n7653 VSS.n7654 0.0732424
R5166 VSS.n7654 VSS.n7655 0.147342
R5167 VSS.n7657 VSS.n7661 0.0721009
R5168 VSS.n7662 VSS.n7658 4.5005
R5169 VSS.n7663 VSS.n7659 4.5005
R5170 VSS.n7664 VSS.n7660 4.5005
R5171 VSS.n7650 VSS.n7661 4.57442
R5172 VSS.n7657 VSS.n7658 0.147342
R5173 VSS.n7658 VSS.n7659 0.147342
R5174 VSS.n7659 VSS.n7660 0.147342
R5175 VSS.n7661 VSS.n7662 2.39784
R5176 VSS.n7662 VSS.n7663 0.147342
R5177 VSS.n7663 VSS.n7664 0.147342
R5178 VSS.n7664 VSS.t455 3.13212
R5179 VSS.n7637 VSS.n7642 4.5005
R5180 VSS.n7639 VSS.n7643 4.5005
R5181 VSS.n7640 VSS.n7644 4.5005
R5182 VSS.n7641 VSS.n7645 4.57324
R5183 VSS.n7637 VSS.n7635 0.147342
R5184 VSS.n7638 VSS.n7639 0.0732424
R5185 VSS.n7639 VSS.n7640 0.147342
R5186 VSS.n7642 VSS.n7646 0.0721009
R5187 VSS.n7647 VSS.n7643 4.5005
R5188 VSS.n7648 VSS.n7644 4.5005
R5189 VSS.n7649 VSS.n7645 4.5005
R5190 VSS.n7635 VSS.n7646 4.57442
R5191 VSS.n7642 VSS.n7643 0.147342
R5192 VSS.n7643 VSS.n7644 0.147342
R5193 VSS.n7644 VSS.n7645 0.147342
R5194 VSS.n7646 VSS.n7647 2.39784
R5195 VSS.n7647 VSS.n7648 0.147342
R5196 VSS.n7648 VSS.n7649 0.147342
R5197 VSS.n7649 VSS.t587 3.13212
R5198 VSS.n7622 VSS.n7627 4.5005
R5199 VSS.n7624 VSS.n7628 4.5005
R5200 VSS.n7625 VSS.n7629 4.5005
R5201 VSS.n7626 VSS.n7630 4.57324
R5202 VSS.n7622 VSS.n7620 0.147342
R5203 VSS.n7623 VSS.n7624 0.0732424
R5204 VSS.n7624 VSS.n7625 0.147342
R5205 VSS.n7627 VSS.n7631 0.0721009
R5206 VSS.n7632 VSS.n7628 4.5005
R5207 VSS.n7633 VSS.n7629 4.5005
R5208 VSS.n7634 VSS.n7630 4.5005
R5209 VSS.n7620 VSS.n7631 4.57442
R5210 VSS.n7627 VSS.n7628 0.147342
R5211 VSS.n7628 VSS.n7629 0.147342
R5212 VSS.n7629 VSS.n7630 0.147342
R5213 VSS.n7631 VSS.n7632 2.39784
R5214 VSS.n7632 VSS.n7633 0.147342
R5215 VSS.n7633 VSS.n7634 0.147342
R5216 VSS.n7634 VSS.t65 3.13212
R5217 VSS.n7607 VSS.n7612 4.5005
R5218 VSS.n7609 VSS.n7613 4.5005
R5219 VSS.n7610 VSS.n7614 4.5005
R5220 VSS.n7611 VSS.n7615 4.57324
R5221 VSS.n7607 VSS.n7605 0.147342
R5222 VSS.n7608 VSS.n7609 0.0732424
R5223 VSS.n7609 VSS.n7610 0.147342
R5224 VSS.n7612 VSS.n7616 0.0721009
R5225 VSS.n7617 VSS.n7613 4.5005
R5226 VSS.n7618 VSS.n7614 4.5005
R5227 VSS.n7619 VSS.n7615 4.5005
R5228 VSS.n7605 VSS.n7616 4.57442
R5229 VSS.n7612 VSS.n7613 0.147342
R5230 VSS.n7613 VSS.n7614 0.147342
R5231 VSS.n7614 VSS.n7615 0.147342
R5232 VSS.n7616 VSS.n7617 2.39784
R5233 VSS.n7617 VSS.n7618 0.147342
R5234 VSS.n7618 VSS.n7619 0.147342
R5235 VSS.n7619 VSS.t79 3.13212
R5236 VSS.n7592 VSS.n7597 4.5005
R5237 VSS.n7594 VSS.n7598 4.5005
R5238 VSS.n7595 VSS.n7599 4.5005
R5239 VSS.n7596 VSS.n7600 4.57324
R5240 VSS.n7592 VSS.n7590 0.147342
R5241 VSS.n7593 VSS.n7594 0.0732424
R5242 VSS.n7594 VSS.n7595 0.147342
R5243 VSS.n7597 VSS.n7601 0.0721009
R5244 VSS.n7602 VSS.n7598 4.5005
R5245 VSS.n7603 VSS.n7599 4.5005
R5246 VSS.n7604 VSS.n7600 4.5005
R5247 VSS.n7590 VSS.n7601 4.57442
R5248 VSS.n7597 VSS.n7598 0.147342
R5249 VSS.n7598 VSS.n7599 0.147342
R5250 VSS.n7599 VSS.n7600 0.147342
R5251 VSS.n7601 VSS.n7602 2.39784
R5252 VSS.n7602 VSS.n7603 0.147342
R5253 VSS.n7603 VSS.n7604 0.147342
R5254 VSS.n7604 VSS.t449 3.13212
R5255 VSS.n7582 VSS.n7577 4.5005
R5256 VSS.n7583 VSS.n7579 4.5005
R5257 VSS.n7584 VSS.n7580 4.5005
R5258 VSS.n7585 VSS.n7581 4.57324
R5259 VSS.n7575 VSS.n7577 0.147342
R5260 VSS.n7578 VSS.n7579 0.0732424
R5261 VSS.n7579 VSS.n7580 0.147342
R5262 VSS.n7586 VSS.n7582 0.0722544
R5263 VSS.n7587 VSS.n7583 4.5005
R5264 VSS.n7588 VSS.n7584 4.5005
R5265 VSS.n7589 VSS.n7585 4.5005
R5266 VSS.n7586 VSS.n7575 4.57426
R5267 VSS.n7582 VSS.n7583 0.147342
R5268 VSS.n7583 VSS.n7584 0.147342
R5269 VSS.n7584 VSS.n7585 0.147342
R5270 VSS.n7587 VSS.n7586 2.37296
R5271 VSS.n7588 VSS.n7587 0.127318
R5272 VSS.n7589 VSS.n7588 0.127318
R5273 VSS.t41 VSS.n7589 2.73618
R5274 VSS.n7562 VSS.n7567 4.5005
R5275 VSS.n7564 VSS.n7568 4.5005
R5276 VSS.n7565 VSS.n7569 4.5005
R5277 VSS.n7566 VSS.n7570 4.57324
R5278 VSS.n7562 VSS.n7560 0.147342
R5279 VSS.n7563 VSS.n7564 0.0732424
R5280 VSS.n7564 VSS.n7565 0.147342
R5281 VSS.n7567 VSS.n7571 0.0721009
R5282 VSS.n7572 VSS.n7568 4.5005
R5283 VSS.n7573 VSS.n7569 4.5005
R5284 VSS.n7574 VSS.n7570 4.5005
R5285 VSS.n7560 VSS.n7571 4.57442
R5286 VSS.n7567 VSS.n7568 0.147342
R5287 VSS.n7568 VSS.n7569 0.147342
R5288 VSS.n7569 VSS.n7570 0.147342
R5289 VSS.n7571 VSS.n7572 2.39784
R5290 VSS.n7572 VSS.n7573 0.147342
R5291 VSS.n7573 VSS.n7574 0.147342
R5292 VSS.n7574 VSS.t610 3.13212
R5293 VSS.n7547 VSS.n7552 4.5005
R5294 VSS.n7549 VSS.n7553 4.5005
R5295 VSS.n7550 VSS.n7554 4.5005
R5296 VSS.n7551 VSS.n7555 4.57324
R5297 VSS.n7547 VSS.n7545 0.147342
R5298 VSS.n7548 VSS.n7549 0.0732424
R5299 VSS.n7549 VSS.n7550 0.147342
R5300 VSS.n7552 VSS.n7556 0.0721009
R5301 VSS.n7557 VSS.n7553 4.5005
R5302 VSS.n7558 VSS.n7554 4.5005
R5303 VSS.n7559 VSS.n7555 4.5005
R5304 VSS.n7545 VSS.n7556 4.57442
R5305 VSS.n7552 VSS.n7553 0.147342
R5306 VSS.n7553 VSS.n7554 0.147342
R5307 VSS.n7554 VSS.n7555 0.147342
R5308 VSS.n7556 VSS.n7557 2.39784
R5309 VSS.n7557 VSS.n7558 0.147342
R5310 VSS.n7558 VSS.n7559 0.147342
R5311 VSS.n7559 VSS.t52 3.13212
R5312 VSS.n7532 VSS.n7537 4.5005
R5313 VSS.n7534 VSS.n7538 4.5005
R5314 VSS.n7535 VSS.n7539 4.5005
R5315 VSS.n7536 VSS.n7540 4.57324
R5316 VSS.n7532 VSS.n7530 0.147342
R5317 VSS.n7533 VSS.n7534 0.0732424
R5318 VSS.n7534 VSS.n7535 0.147342
R5319 VSS.n7537 VSS.n7541 0.0721009
R5320 VSS.n7542 VSS.n7538 4.5005
R5321 VSS.n7543 VSS.n7539 4.5005
R5322 VSS.n7544 VSS.n7540 4.5005
R5323 VSS.n7530 VSS.n7541 4.57442
R5324 VSS.n7537 VSS.n7538 0.147342
R5325 VSS.n7538 VSS.n7539 0.147342
R5326 VSS.n7539 VSS.n7540 0.147342
R5327 VSS.n7541 VSS.n7542 2.39784
R5328 VSS.n7542 VSS.n7543 0.147342
R5329 VSS.n7543 VSS.n7544 0.147342
R5330 VSS.n7544 VSS.t535 3.13212
R5331 VSS.n7522 VSS.n7517 4.5005
R5332 VSS.n7523 VSS.n7519 4.5005
R5333 VSS.n7524 VSS.n7520 4.5005
R5334 VSS.n7525 VSS.n7521 4.57324
R5335 VSS.n7515 VSS.n7517 0.147342
R5336 VSS.n7518 VSS.n7519 0.0732424
R5337 VSS.n7519 VSS.n7520 0.147342
R5338 VSS.n7526 VSS.n7522 0.0722544
R5339 VSS.n7527 VSS.n7523 4.5005
R5340 VSS.n7528 VSS.n7524 4.5005
R5341 VSS.n7529 VSS.n7525 4.5005
R5342 VSS.n7526 VSS.n7515 4.57426
R5343 VSS.n7522 VSS.n7523 0.147342
R5344 VSS.n7523 VSS.n7524 0.147342
R5345 VSS.n7524 VSS.n7525 0.147342
R5346 VSS.n7527 VSS.n7526 2.37296
R5347 VSS.n7528 VSS.n7527 0.127318
R5348 VSS.n7529 VSS.n7528 0.127318
R5349 VSS.t41 VSS.n7529 2.73618
R5350 VSS.n7502 VSS.n7507 4.5005
R5351 VSS.n7504 VSS.n7508 4.5005
R5352 VSS.n7505 VSS.n7509 4.5005
R5353 VSS.n7506 VSS.n7510 4.57324
R5354 VSS.n7502 VSS.n7500 0.147342
R5355 VSS.n7503 VSS.n7504 0.0732424
R5356 VSS.n7504 VSS.n7505 0.147342
R5357 VSS.n7507 VSS.n7511 0.0721009
R5358 VSS.n7512 VSS.n7508 4.5005
R5359 VSS.n7513 VSS.n7509 4.5005
R5360 VSS.n7514 VSS.n7510 4.5005
R5361 VSS.n7500 VSS.n7511 4.57442
R5362 VSS.n7507 VSS.n7508 0.147342
R5363 VSS.n7508 VSS.n7509 0.147342
R5364 VSS.n7509 VSS.n7510 0.147342
R5365 VSS.n7511 VSS.n7512 2.39784
R5366 VSS.n7512 VSS.n7513 0.147342
R5367 VSS.n7513 VSS.n7514 0.147342
R5368 VSS.n7514 VSS.t111 3.13212
R5369 VSS.n7487 VSS.n7492 4.5005
R5370 VSS.n7489 VSS.n7493 4.5005
R5371 VSS.n7490 VSS.n7494 4.5005
R5372 VSS.n7491 VSS.n7495 4.57324
R5373 VSS.n7487 VSS.n7485 0.147342
R5374 VSS.n7488 VSS.n7489 0.0732424
R5375 VSS.n7489 VSS.n7490 0.147342
R5376 VSS.n7492 VSS.n7496 0.0721009
R5377 VSS.n7497 VSS.n7493 4.5005
R5378 VSS.n7498 VSS.n7494 4.5005
R5379 VSS.n7499 VSS.n7495 4.5005
R5380 VSS.n7485 VSS.n7496 4.57442
R5381 VSS.n7492 VSS.n7493 0.147342
R5382 VSS.n7493 VSS.n7494 0.147342
R5383 VSS.n7494 VSS.n7495 0.147342
R5384 VSS.n7496 VSS.n7497 2.39784
R5385 VSS.n7497 VSS.n7498 0.147342
R5386 VSS.n7498 VSS.n7499 0.147342
R5387 VSS.n7499 VSS.t498 3.13212
R5388 VSS.n7472 VSS.n7477 4.5005
R5389 VSS.n7474 VSS.n7478 4.5005
R5390 VSS.n7475 VSS.n7479 4.5005
R5391 VSS.n7476 VSS.n7480 4.57324
R5392 VSS.n7472 VSS.n7470 0.147342
R5393 VSS.n7473 VSS.n7474 0.0732424
R5394 VSS.n7474 VSS.n7475 0.147342
R5395 VSS.n7477 VSS.n7481 0.0721009
R5396 VSS.n7482 VSS.n7478 4.5005
R5397 VSS.n7483 VSS.n7479 4.5005
R5398 VSS.n7484 VSS.n7480 4.5005
R5399 VSS.n7470 VSS.n7481 4.57442
R5400 VSS.n7477 VSS.n7478 0.147342
R5401 VSS.n7478 VSS.n7479 0.147342
R5402 VSS.n7479 VSS.n7480 0.147342
R5403 VSS.n7481 VSS.n7482 2.39784
R5404 VSS.n7482 VSS.n7483 0.147342
R5405 VSS.n7483 VSS.n7484 0.147342
R5406 VSS.n7484 VSS.t43 3.13212
R5407 VSS.n7457 VSS.n7462 4.5005
R5408 VSS.n7459 VSS.n7463 4.5005
R5409 VSS.n7460 VSS.n7464 4.5005
R5410 VSS.n7461 VSS.n7465 4.57324
R5411 VSS.n7457 VSS.n7455 0.147342
R5412 VSS.n7458 VSS.n7459 0.0732424
R5413 VSS.n7459 VSS.n7460 0.147342
R5414 VSS.n7462 VSS.n7466 0.0721009
R5415 VSS.n7467 VSS.n7463 4.5005
R5416 VSS.n7468 VSS.n7464 4.5005
R5417 VSS.n7469 VSS.n7465 4.5005
R5418 VSS.n7455 VSS.n7466 4.57442
R5419 VSS.n7462 VSS.n7463 0.147342
R5420 VSS.n7463 VSS.n7464 0.147342
R5421 VSS.n7464 VSS.n7465 0.147342
R5422 VSS.n7466 VSS.n7467 2.39784
R5423 VSS.n7467 VSS.n7468 0.147342
R5424 VSS.n7468 VSS.n7469 0.147342
R5425 VSS.n7469 VSS.t607 3.13212
R5426 VSS.n7447 VSS.n7442 4.5005
R5427 VSS.n7448 VSS.n7444 4.5005
R5428 VSS.n7449 VSS.n7445 4.5005
R5429 VSS.n7450 VSS.n7446 4.57324
R5430 VSS.n7440 VSS.n7442 0.147342
R5431 VSS.n7443 VSS.n7444 0.0732424
R5432 VSS.n7444 VSS.n7445 0.147342
R5433 VSS.n7451 VSS.n7447 0.0722544
R5434 VSS.n7452 VSS.n7448 4.5005
R5435 VSS.n7453 VSS.n7449 4.5005
R5436 VSS.n7454 VSS.n7450 4.5005
R5437 VSS.n7451 VSS.n7440 4.57426
R5438 VSS.n7447 VSS.n7448 0.147342
R5439 VSS.n7448 VSS.n7449 0.147342
R5440 VSS.n7449 VSS.n7450 0.147342
R5441 VSS.n7452 VSS.n7451 2.37296
R5442 VSS.n7453 VSS.n7452 0.127318
R5443 VSS.n7454 VSS.n7453 0.127318
R5444 VSS.t41 VSS.n7454 2.73618
R5445 VSS.n7427 VSS.n7432 4.5005
R5446 VSS.n7429 VSS.n7433 4.5005
R5447 VSS.n7430 VSS.n7434 4.5005
R5448 VSS.n7431 VSS.n7435 4.57324
R5449 VSS.n7427 VSS.n7425 0.147342
R5450 VSS.n7428 VSS.n7429 0.0732424
R5451 VSS.n7429 VSS.n7430 0.147342
R5452 VSS.n7432 VSS.n7436 0.0721009
R5453 VSS.n7437 VSS.n7433 4.5005
R5454 VSS.n7438 VSS.n7434 4.5005
R5455 VSS.n7439 VSS.n7435 4.5005
R5456 VSS.n7425 VSS.n7436 4.57442
R5457 VSS.n7432 VSS.n7433 0.147342
R5458 VSS.n7433 VSS.n7434 0.147342
R5459 VSS.n7434 VSS.n7435 0.147342
R5460 VSS.n7436 VSS.n7437 2.39784
R5461 VSS.n7437 VSS.n7438 0.147342
R5462 VSS.n7438 VSS.n7439 0.147342
R5463 VSS.n7439 VSS.t54 3.13212
R5464 VSS.n7412 VSS.n7417 4.5005
R5465 VSS.n7414 VSS.n7418 4.5005
R5466 VSS.n7415 VSS.n7419 4.5005
R5467 VSS.n7416 VSS.n7420 4.57324
R5468 VSS.n7412 VSS.n7410 0.147342
R5469 VSS.n7413 VSS.n7414 0.0732424
R5470 VSS.n7414 VSS.n7415 0.147342
R5471 VSS.n7417 VSS.n7421 0.0721009
R5472 VSS.n7422 VSS.n7418 4.5005
R5473 VSS.n7423 VSS.n7419 4.5005
R5474 VSS.n7424 VSS.n7420 4.5005
R5475 VSS.n7410 VSS.n7421 4.57442
R5476 VSS.n7417 VSS.n7418 0.147342
R5477 VSS.n7418 VSS.n7419 0.147342
R5478 VSS.n7419 VSS.n7420 0.147342
R5479 VSS.n7421 VSS.n7422 2.39784
R5480 VSS.n7422 VSS.n7423 0.147342
R5481 VSS.n7423 VSS.n7424 0.147342
R5482 VSS.n7424 VSS.t199 3.13212
R5483 VSS.n7397 VSS.n7402 4.5005
R5484 VSS.n7399 VSS.n7403 4.5005
R5485 VSS.n7400 VSS.n7404 4.5005
R5486 VSS.n7401 VSS.n7405 4.57324
R5487 VSS.n7397 VSS.n7395 0.147342
R5488 VSS.n7398 VSS.n7399 0.0732424
R5489 VSS.n7399 VSS.n7400 0.147342
R5490 VSS.n7402 VSS.n7406 0.0721009
R5491 VSS.n7407 VSS.n7403 4.5005
R5492 VSS.n7408 VSS.n7404 4.5005
R5493 VSS.n7409 VSS.n7405 4.5005
R5494 VSS.n7395 VSS.n7406 4.57442
R5495 VSS.n7402 VSS.n7403 0.147342
R5496 VSS.n7403 VSS.n7404 0.147342
R5497 VSS.n7404 VSS.n7405 0.147342
R5498 VSS.n7406 VSS.n7407 2.39784
R5499 VSS.n7407 VSS.n7408 0.147342
R5500 VSS.n7408 VSS.n7409 0.147342
R5501 VSS.n7409 VSS.t422 3.13212
R5502 VSS.n7387 VSS.n7382 4.5005
R5503 VSS.n7388 VSS.n7384 4.5005
R5504 VSS.n7389 VSS.n7385 4.5005
R5505 VSS.n7390 VSS.n7386 4.57324
R5506 VSS.n7380 VSS.n7382 0.147342
R5507 VSS.n7383 VSS.n7384 0.0732424
R5508 VSS.n7384 VSS.n7385 0.147342
R5509 VSS.n7391 VSS.n7387 0.0722544
R5510 VSS.n7392 VSS.n7388 4.5005
R5511 VSS.n7393 VSS.n7389 4.5005
R5512 VSS.n7394 VSS.n7390 4.5005
R5513 VSS.n7391 VSS.n7380 4.57426
R5514 VSS.n7387 VSS.n7388 0.147342
R5515 VSS.n7388 VSS.n7389 0.147342
R5516 VSS.n7389 VSS.n7390 0.147342
R5517 VSS.n7392 VSS.n7391 2.37296
R5518 VSS.n7393 VSS.n7392 0.127318
R5519 VSS.n7394 VSS.n7393 0.127318
R5520 VSS.t41 VSS.n7394 2.73618
R5521 VSS.n7367 VSS.n7372 4.5005
R5522 VSS.n7369 VSS.n7373 4.5005
R5523 VSS.n7370 VSS.n7374 4.5005
R5524 VSS.n7371 VSS.n7375 4.57324
R5525 VSS.n7367 VSS.n7365 0.147342
R5526 VSS.n7368 VSS.n7369 0.0732424
R5527 VSS.n7369 VSS.n7370 0.147342
R5528 VSS.n7372 VSS.n7376 0.0721009
R5529 VSS.n7377 VSS.n7373 4.5005
R5530 VSS.n7378 VSS.n7374 4.5005
R5531 VSS.n7379 VSS.n7375 4.5005
R5532 VSS.n7365 VSS.n7376 4.57442
R5533 VSS.n7372 VSS.n7373 0.147342
R5534 VSS.n7373 VSS.n7374 0.147342
R5535 VSS.n7374 VSS.n7375 0.147342
R5536 VSS.n7376 VSS.n7377 2.39784
R5537 VSS.n7377 VSS.n7378 0.147342
R5538 VSS.n7378 VSS.n7379 0.147342
R5539 VSS.n7379 VSS.t555 3.13212
R5540 VSS.n7352 VSS.n7357 4.5005
R5541 VSS.n7354 VSS.n7358 4.5005
R5542 VSS.n7355 VSS.n7359 4.5005
R5543 VSS.n7356 VSS.n7360 4.57324
R5544 VSS.n7352 VSS.n7350 0.147342
R5545 VSS.n7353 VSS.n7354 0.0732424
R5546 VSS.n7354 VSS.n7355 0.147342
R5547 VSS.n7357 VSS.n7361 0.0721009
R5548 VSS.n7362 VSS.n7358 4.5005
R5549 VSS.n7363 VSS.n7359 4.5005
R5550 VSS.n7364 VSS.n7360 4.5005
R5551 VSS.n7350 VSS.n7361 4.57442
R5552 VSS.n7357 VSS.n7358 0.147342
R5553 VSS.n7358 VSS.n7359 0.147342
R5554 VSS.n7359 VSS.n7360 0.147342
R5555 VSS.n7361 VSS.n7362 2.39784
R5556 VSS.n7362 VSS.n7363 0.147342
R5557 VSS.n7363 VSS.n7364 0.147342
R5558 VSS.n7364 VSS.t456 3.13212
R5559 VSS.n7337 VSS.n7342 4.5005
R5560 VSS.n7339 VSS.n7343 4.5005
R5561 VSS.n7340 VSS.n7344 4.5005
R5562 VSS.n7341 VSS.n7345 4.57324
R5563 VSS.n7337 VSS.n7335 0.147342
R5564 VSS.n7338 VSS.n7339 0.0732424
R5565 VSS.n7339 VSS.n7340 0.147342
R5566 VSS.n7342 VSS.n7346 0.0721009
R5567 VSS.n7347 VSS.n7343 4.5005
R5568 VSS.n7348 VSS.n7344 4.5005
R5569 VSS.n7349 VSS.n7345 4.5005
R5570 VSS.n7335 VSS.n7346 4.57442
R5571 VSS.n7342 VSS.n7343 0.147342
R5572 VSS.n7343 VSS.n7344 0.147342
R5573 VSS.n7344 VSS.n7345 0.147342
R5574 VSS.n7346 VSS.n7347 2.39784
R5575 VSS.n7347 VSS.n7348 0.147342
R5576 VSS.n7348 VSS.n7349 0.147342
R5577 VSS.n7349 VSS.t592 3.13212
R5578 VSS.n7322 VSS.n7327 4.5005
R5579 VSS.n7324 VSS.n7328 4.5005
R5580 VSS.n7325 VSS.n7329 4.5005
R5581 VSS.n7326 VSS.n7330 4.57324
R5582 VSS.n7322 VSS.n7320 0.147342
R5583 VSS.n7323 VSS.n7324 0.0732424
R5584 VSS.n7324 VSS.n7325 0.147342
R5585 VSS.n7327 VSS.n7331 0.0721009
R5586 VSS.n7332 VSS.n7328 4.5005
R5587 VSS.n7333 VSS.n7329 4.5005
R5588 VSS.n7334 VSS.n7330 4.5005
R5589 VSS.n7320 VSS.n7331 4.57442
R5590 VSS.n7327 VSS.n7328 0.147342
R5591 VSS.n7328 VSS.n7329 0.147342
R5592 VSS.n7329 VSS.n7330 0.147342
R5593 VSS.n7331 VSS.n7332 2.39784
R5594 VSS.n7332 VSS.n7333 0.147342
R5595 VSS.n7333 VSS.n7334 0.147342
R5596 VSS.n7334 VSS.t487 3.13212
R5597 VSS.n7307 VSS.n7312 4.5005
R5598 VSS.n7309 VSS.n7313 4.5005
R5599 VSS.n7310 VSS.n7314 4.5005
R5600 VSS.n7311 VSS.n7315 4.57324
R5601 VSS.n7307 VSS.n7305 0.147342
R5602 VSS.n7308 VSS.n7309 0.0732424
R5603 VSS.n7309 VSS.n7310 0.147342
R5604 VSS.n7312 VSS.n7316 0.0721009
R5605 VSS.n7317 VSS.n7313 4.5005
R5606 VSS.n7318 VSS.n7314 4.5005
R5607 VSS.n7319 VSS.n7315 4.5005
R5608 VSS.n7305 VSS.n7316 4.57442
R5609 VSS.n7312 VSS.n7313 0.147342
R5610 VSS.n7313 VSS.n7314 0.147342
R5611 VSS.n7314 VSS.n7315 0.147342
R5612 VSS.n7316 VSS.n7317 2.39784
R5613 VSS.n7317 VSS.n7318 0.147342
R5614 VSS.n7318 VSS.n7319 0.147342
R5615 VSS.n7319 VSS.t117 3.13212
R5616 VSS.n7292 VSS.n7297 4.5005
R5617 VSS.n7294 VSS.n7298 4.5005
R5618 VSS.n7295 VSS.n7299 4.5005
R5619 VSS.n7296 VSS.n7300 4.57324
R5620 VSS.n7292 VSS.n7290 0.147342
R5621 VSS.n7293 VSS.n7294 0.0732424
R5622 VSS.n7294 VSS.n7295 0.147342
R5623 VSS.n7297 VSS.n7301 0.0721009
R5624 VSS.n7302 VSS.n7298 4.5005
R5625 VSS.n7303 VSS.n7299 4.5005
R5626 VSS.n7304 VSS.n7300 4.5005
R5627 VSS.n7290 VSS.n7301 4.57442
R5628 VSS.n7297 VSS.n7298 0.147342
R5629 VSS.n7298 VSS.n7299 0.147342
R5630 VSS.n7299 VSS.n7300 0.147342
R5631 VSS.n7301 VSS.n7302 2.39784
R5632 VSS.n7302 VSS.n7303 0.147342
R5633 VSS.n7303 VSS.n7304 0.147342
R5634 VSS.n7304 VSS.t476 3.13212
R5635 VSS.n7282 VSS.n7277 4.5005
R5636 VSS.n7283 VSS.n7279 4.5005
R5637 VSS.n7284 VSS.n7280 4.5005
R5638 VSS.n7285 VSS.n7281 4.57324
R5639 VSS.n7275 VSS.n7277 0.147342
R5640 VSS.n7278 VSS.n7279 0.0732424
R5641 VSS.n7279 VSS.n7280 0.147342
R5642 VSS.n7286 VSS.n7282 0.0722544
R5643 VSS.n7287 VSS.n7283 4.5005
R5644 VSS.n7288 VSS.n7284 4.5005
R5645 VSS.n7289 VSS.n7285 4.5005
R5646 VSS.n7286 VSS.n7275 4.57426
R5647 VSS.n7282 VSS.n7283 0.147342
R5648 VSS.n7283 VSS.n7284 0.147342
R5649 VSS.n7284 VSS.n7285 0.147342
R5650 VSS.n7287 VSS.n7286 2.37296
R5651 VSS.n7288 VSS.n7287 0.127318
R5652 VSS.n7289 VSS.n7288 0.127318
R5653 VSS.t41 VSS.n7289 2.73618
R5654 VSS.n7262 VSS.n7267 4.5005
R5655 VSS.n7264 VSS.n7268 4.5005
R5656 VSS.n7265 VSS.n7269 4.5005
R5657 VSS.n7266 VSS.n7270 4.57324
R5658 VSS.n7262 VSS.n7260 0.147342
R5659 VSS.n7263 VSS.n7264 0.0732424
R5660 VSS.n7264 VSS.n7265 0.147342
R5661 VSS.n7267 VSS.n7271 0.0721009
R5662 VSS.n7272 VSS.n7268 4.5005
R5663 VSS.n7273 VSS.n7269 4.5005
R5664 VSS.n7274 VSS.n7270 4.5005
R5665 VSS.n7260 VSS.n7271 4.57442
R5666 VSS.n7267 VSS.n7268 0.147342
R5667 VSS.n7268 VSS.n7269 0.147342
R5668 VSS.n7269 VSS.n7270 0.147342
R5669 VSS.n7271 VSS.n7272 2.39784
R5670 VSS.n7272 VSS.n7273 0.147342
R5671 VSS.n7273 VSS.n7274 0.147342
R5672 VSS.n7274 VSS.t611 3.13212
R5673 VSS.n7247 VSS.n7252 4.5005
R5674 VSS.n7249 VSS.n7253 4.5005
R5675 VSS.n7250 VSS.n7254 4.5005
R5676 VSS.n7251 VSS.n7255 4.57324
R5677 VSS.n7247 VSS.n7245 0.147342
R5678 VSS.n7248 VSS.n7249 0.0732424
R5679 VSS.n7249 VSS.n7250 0.147342
R5680 VSS.n7252 VSS.n7256 0.0721009
R5681 VSS.n7257 VSS.n7253 4.5005
R5682 VSS.n7258 VSS.n7254 4.5005
R5683 VSS.n7259 VSS.n7255 4.5005
R5684 VSS.n7245 VSS.n7256 4.57442
R5685 VSS.n7252 VSS.n7253 0.147342
R5686 VSS.n7253 VSS.n7254 0.147342
R5687 VSS.n7254 VSS.n7255 0.147342
R5688 VSS.n7256 VSS.n7257 2.39784
R5689 VSS.n7257 VSS.n7258 0.147342
R5690 VSS.n7258 VSS.n7259 0.147342
R5691 VSS.n7259 VSS.t50 3.13212
R5692 VSS.n7232 VSS.n7237 4.5005
R5693 VSS.n7234 VSS.n7238 4.5005
R5694 VSS.n7235 VSS.n7239 4.5005
R5695 VSS.n7236 VSS.n7240 4.57324
R5696 VSS.n7232 VSS.n7230 0.147342
R5697 VSS.n7233 VSS.n7234 0.0732424
R5698 VSS.n7234 VSS.n7235 0.147342
R5699 VSS.n7237 VSS.n7241 0.0721009
R5700 VSS.n7242 VSS.n7238 4.5005
R5701 VSS.n7243 VSS.n7239 4.5005
R5702 VSS.n7244 VSS.n7240 4.5005
R5703 VSS.n7230 VSS.n7241 4.57442
R5704 VSS.n7237 VSS.n7238 0.147342
R5705 VSS.n7238 VSS.n7239 0.147342
R5706 VSS.n7239 VSS.n7240 0.147342
R5707 VSS.n7241 VSS.n7242 2.39784
R5708 VSS.n7242 VSS.n7243 0.147342
R5709 VSS.n7243 VSS.n7244 0.147342
R5710 VSS.n7244 VSS.t536 3.13212
R5711 VSS.n7222 VSS.n7217 4.5005
R5712 VSS.n7223 VSS.n7219 4.5005
R5713 VSS.n7224 VSS.n7220 4.5005
R5714 VSS.n7225 VSS.n7221 4.57324
R5715 VSS.n7215 VSS.n7217 0.147342
R5716 VSS.n7218 VSS.n7219 0.0732424
R5717 VSS.n7219 VSS.n7220 0.147342
R5718 VSS.n7226 VSS.n7222 0.0722544
R5719 VSS.n7227 VSS.n7223 4.5005
R5720 VSS.n7228 VSS.n7224 4.5005
R5721 VSS.n7229 VSS.n7225 4.5005
R5722 VSS.n7226 VSS.n7215 4.57426
R5723 VSS.n7222 VSS.n7223 0.147342
R5724 VSS.n7223 VSS.n7224 0.147342
R5725 VSS.n7224 VSS.n7225 0.147342
R5726 VSS.n7227 VSS.n7226 2.37296
R5727 VSS.n7228 VSS.n7227 0.127318
R5728 VSS.n7229 VSS.n7228 0.127318
R5729 VSS.t41 VSS.n7229 2.73618
R5730 VSS.n7202 VSS.n7207 4.5005
R5731 VSS.n7204 VSS.n7208 4.5005
R5732 VSS.n7205 VSS.n7209 4.5005
R5733 VSS.n7206 VSS.n7210 4.57324
R5734 VSS.n7202 VSS.n7200 0.147342
R5735 VSS.n7203 VSS.n7204 0.0732424
R5736 VSS.n7204 VSS.n7205 0.147342
R5737 VSS.n7207 VSS.n7211 0.0721009
R5738 VSS.n7212 VSS.n7208 4.5005
R5739 VSS.n7213 VSS.n7209 4.5005
R5740 VSS.n7214 VSS.n7210 4.5005
R5741 VSS.n7200 VSS.n7211 4.57442
R5742 VSS.n7207 VSS.n7208 0.147342
R5743 VSS.n7208 VSS.n7209 0.147342
R5744 VSS.n7209 VSS.n7210 0.147342
R5745 VSS.n7211 VSS.n7212 2.39784
R5746 VSS.n7212 VSS.n7213 0.147342
R5747 VSS.n7213 VSS.n7214 0.147342
R5748 VSS.n7214 VSS.t148 3.13212
R5749 VSS.n7187 VSS.n7192 4.5005
R5750 VSS.n7189 VSS.n7193 4.5005
R5751 VSS.n7190 VSS.n7194 4.5005
R5752 VSS.n7191 VSS.n7195 4.57324
R5753 VSS.n7187 VSS.n7185 0.147342
R5754 VSS.n7188 VSS.n7189 0.0732424
R5755 VSS.n7189 VSS.n7190 0.147342
R5756 VSS.n7192 VSS.n7196 0.0721009
R5757 VSS.n7197 VSS.n7193 4.5005
R5758 VSS.n7198 VSS.n7194 4.5005
R5759 VSS.n7199 VSS.n7195 4.5005
R5760 VSS.n7185 VSS.n7196 4.57442
R5761 VSS.n7192 VSS.n7193 0.147342
R5762 VSS.n7193 VSS.n7194 0.147342
R5763 VSS.n7194 VSS.n7195 0.147342
R5764 VSS.n7196 VSS.n7197 2.39784
R5765 VSS.n7197 VSS.n7198 0.147342
R5766 VSS.n7198 VSS.n7199 0.147342
R5767 VSS.n7199 VSS.t473 3.13212
R5768 VSS.n4770 VSS.n4771 0.0722544
R5769 VSS.n4772 VSS.n4773 4.5005
R5770 VSS.n4774 VSS.n4775 4.5005
R5771 VSS.n4776 VSS.n4777 4.5005
R5772 VSS.n4772 VSS.n4770 2.37296
R5773 VSS.n4774 VSS.n4772 0.127318
R5774 VSS.n4776 VSS.n4774 0.127318
R5775 VSS.t0 VSS.n4776 2.73618
R5776 VSS.n4771 VSS.n4778 4.5005
R5777 VSS.n4773 VSS.n4779 4.5005
R5778 VSS.n4775 VSS.n4780 4.5005
R5779 VSS.n4777 VSS.n4781 4.5005
R5780 VSS.n4783 VSS.n4770 4.647
R5781 VSS.n4771 VSS.n4773 0.147342
R5782 VSS.n4773 VSS.n4775 0.147342
R5783 VSS.n4775 VSS.n4777 0.147342
R5784 VSS.n4783 VSS.n4784 2.21488
R5785 VSS.n4778 VSS.n4783 0.0732424
R5786 VSS.n4782 VSS.n4784 2.21488
R5787 VSS.n4782 VSS.n4780 0.0732424
R5788 VSS.n4781 VSS.n4784 4.5005
R5789 VSS.n4778 VSS.n4779 0.147342
R5790 VSS.n4779 VSS.n4782 0.0732424
R5791 VSS.n4780 VSS.n4781 0.147342
R5792 VSS.n4785 VSS.n4786 4.5005
R5793 VSS.n4788 VSS.n4787 0.0732424
R5794 VSS.n4786 VSS.n4788 2.21488
R5795 VSS.n4791 VSS.n4790 0.0732424
R5796 VSS.n4786 VSS.n4791 2.21488
R5797 VSS.n4800 VSS.n4801 4.5005
R5798 VSS.n4803 VSS.n4802 0.0732424
R5799 VSS.n4801 VSS.n4803 2.21488
R5800 VSS.n4806 VSS.n4805 0.0732424
R5801 VSS.n4801 VSS.n4806 2.21488
R5802 VSS.n4815 VSS.n4816 4.5005
R5803 VSS.n4817 VSS.n4818 0.0732424
R5804 VSS.n4818 VSS.n4816 2.21488
R5805 VSS.n4820 VSS.n4821 0.0732424
R5806 VSS.n4821 VSS.n4816 2.21488
R5807 VSS.n4830 VSS.n4831 4.5005
R5808 VSS.n4833 VSS.n4832 0.0732424
R5809 VSS.n4831 VSS.n4833 2.21488
R5810 VSS.n4836 VSS.n4835 0.0732424
R5811 VSS.n4831 VSS.n4836 2.21488
R5812 VSS.n4845 VSS.n4846 4.5005
R5813 VSS.n4848 VSS.n4847 0.0732424
R5814 VSS.n4846 VSS.n4848 2.21488
R5815 VSS.n4851 VSS.n4850 0.0732424
R5816 VSS.n4846 VSS.n4851 2.21488
R5817 VSS.n4860 VSS.n4861 4.5005
R5818 VSS.n4863 VSS.n4862 0.0732424
R5819 VSS.n4861 VSS.n4863 2.21488
R5820 VSS.n4866 VSS.n4865 0.0732424
R5821 VSS.n4861 VSS.n4866 2.21488
R5822 VSS.n4875 VSS.n4876 4.5005
R5823 VSS.n4877 VSS.n4878 0.0732424
R5824 VSS.n4878 VSS.n4876 2.21488
R5825 VSS.n4880 VSS.n4881 0.0732424
R5826 VSS.n4881 VSS.n4876 2.21488
R5827 VSS.n4890 VSS.n4891 4.5005
R5828 VSS.n4893 VSS.n4892 0.0732424
R5829 VSS.n4891 VSS.n4893 2.21488
R5830 VSS.n4896 VSS.n4895 0.0732424
R5831 VSS.n4891 VSS.n4896 2.21488
R5832 VSS.n4905 VSS.n4906 4.5005
R5833 VSS.n4908 VSS.n4907 0.0732424
R5834 VSS.n4906 VSS.n4908 2.21488
R5835 VSS.n4911 VSS.n4910 0.0732424
R5836 VSS.n4906 VSS.n4911 2.21488
R5837 VSS.n4920 VSS.n4921 4.5005
R5838 VSS.n4923 VSS.n4922 0.0732424
R5839 VSS.n4921 VSS.n4923 2.21488
R5840 VSS.n4926 VSS.n4925 0.0732424
R5841 VSS.n4921 VSS.n4926 2.21488
R5842 VSS.n4935 VSS.n4936 4.5005
R5843 VSS.n4938 VSS.n4937 0.0732424
R5844 VSS.n4936 VSS.n4938 2.21488
R5845 VSS.n4941 VSS.n4940 0.0732424
R5846 VSS.n4936 VSS.n4941 2.21488
R5847 VSS.n4950 VSS.n4951 4.5005
R5848 VSS.n4953 VSS.n4952 0.0732424
R5849 VSS.n4951 VSS.n4953 2.21488
R5850 VSS.n4956 VSS.n4955 0.0732424
R5851 VSS.n4951 VSS.n4956 2.21488
R5852 VSS.n4965 VSS.n4966 4.5005
R5853 VSS.n4968 VSS.n4967 0.0732424
R5854 VSS.n4966 VSS.n4968 2.21488
R5855 VSS.n4971 VSS.n4970 0.0732424
R5856 VSS.n4966 VSS.n4971 2.21488
R5857 VSS.n4980 VSS.n4981 4.5005
R5858 VSS.n4982 VSS.n4983 0.0732424
R5859 VSS.n4983 VSS.n4981 2.21488
R5860 VSS.n4985 VSS.n4986 0.0732424
R5861 VSS.n4986 VSS.n4981 2.21488
R5862 VSS.n4995 VSS.n4996 4.5005
R5863 VSS.n4998 VSS.n4997 0.0732424
R5864 VSS.n4996 VSS.n4998 2.21488
R5865 VSS.n5001 VSS.n5000 0.0732424
R5866 VSS.n4996 VSS.n5001 2.21488
R5867 VSS.n5010 VSS.n5011 4.5005
R5868 VSS.n5013 VSS.n5012 0.0732424
R5869 VSS.n5011 VSS.n5013 2.21488
R5870 VSS.n5016 VSS.n5015 0.0732424
R5871 VSS.n5011 VSS.n5016 2.21488
R5872 VSS.n5025 VSS.n5026 4.5005
R5873 VSS.n5028 VSS.n5027 0.0732424
R5874 VSS.n5026 VSS.n5028 2.21488
R5875 VSS.n5031 VSS.n5030 0.0732424
R5876 VSS.n5026 VSS.n5031 2.21488
R5877 VSS.n5040 VSS.n5041 4.5005
R5878 VSS.n5042 VSS.n5043 0.0732424
R5879 VSS.n5043 VSS.n5041 2.21488
R5880 VSS.n5045 VSS.n5046 0.0732424
R5881 VSS.n5046 VSS.n5041 2.21488
R5882 VSS.n5055 VSS.n5056 4.5005
R5883 VSS.n5058 VSS.n5057 0.0732424
R5884 VSS.n5056 VSS.n5058 2.21488
R5885 VSS.n5061 VSS.n5060 0.0732424
R5886 VSS.n5056 VSS.n5061 2.21488
R5887 VSS.n5070 VSS.n5071 4.5005
R5888 VSS.n5073 VSS.n5072 0.0732424
R5889 VSS.n5071 VSS.n5073 2.21488
R5890 VSS.n5076 VSS.n5075 0.0732424
R5891 VSS.n5071 VSS.n5076 2.21488
R5892 VSS.n5085 VSS.n5086 4.5005
R5893 VSS.n5088 VSS.n5087 0.0732424
R5894 VSS.n5086 VSS.n5088 2.21488
R5895 VSS.n5091 VSS.n5090 0.0732424
R5896 VSS.n5086 VSS.n5091 2.21488
R5897 VSS.n5100 VSS.n5101 4.5005
R5898 VSS.n5103 VSS.n5102 0.0732424
R5899 VSS.n5101 VSS.n5103 2.21488
R5900 VSS.n5106 VSS.n5105 0.0732424
R5901 VSS.n5101 VSS.n5106 2.21488
R5902 VSS.n5115 VSS.n5116 4.5005
R5903 VSS.n5117 VSS.n5118 0.0732424
R5904 VSS.n5118 VSS.n5116 2.21488
R5905 VSS.n5120 VSS.n5121 0.0732424
R5906 VSS.n5121 VSS.n5116 2.21488
R5907 VSS.n5130 VSS.n5131 4.5005
R5908 VSS.n5133 VSS.n5132 0.0732424
R5909 VSS.n5131 VSS.n5133 2.21488
R5910 VSS.n5136 VSS.n5135 0.0732424
R5911 VSS.n5131 VSS.n5136 2.21488
R5912 VSS.n5145 VSS.n5146 4.5005
R5913 VSS.n5148 VSS.n5147 0.0732424
R5914 VSS.n5146 VSS.n5148 2.21488
R5915 VSS.n5151 VSS.n5150 0.0732424
R5916 VSS.n5146 VSS.n5151 2.21488
R5917 VSS.n5160 VSS.n5161 4.5005
R5918 VSS.n5163 VSS.n5162 0.0732424
R5919 VSS.n5161 VSS.n5163 2.21488
R5920 VSS.n5166 VSS.n5165 0.0732424
R5921 VSS.n5161 VSS.n5166 2.21488
R5922 VSS.n5175 VSS.n5176 4.5005
R5923 VSS.n5177 VSS.n5178 0.0732424
R5924 VSS.n5178 VSS.n5176 2.21488
R5925 VSS.n5180 VSS.n5181 0.0732424
R5926 VSS.n5181 VSS.n5176 2.21488
R5927 VSS.n5190 VSS.n5191 4.5005
R5928 VSS.n5193 VSS.n5192 0.0732424
R5929 VSS.n5191 VSS.n5193 2.21488
R5930 VSS.n5196 VSS.n5195 0.0732424
R5931 VSS.n5191 VSS.n5196 2.21488
R5932 VSS.n5205 VSS.n5206 4.5005
R5933 VSS.n5208 VSS.n5207 0.0732424
R5934 VSS.n5206 VSS.n5208 2.21488
R5935 VSS.n5211 VSS.n5210 0.0732424
R5936 VSS.n5206 VSS.n5211 2.21488
R5937 VSS.n5220 VSS.n5221 4.5005
R5938 VSS.n5223 VSS.n5222 0.0732424
R5939 VSS.n5221 VSS.n5223 2.21488
R5940 VSS.n5226 VSS.n5225 0.0732424
R5941 VSS.n5221 VSS.n5226 2.21488
R5942 VSS.n5235 VSS.n5236 4.5005
R5943 VSS.n5238 VSS.n5237 0.0732424
R5944 VSS.n5236 VSS.n5238 2.21488
R5945 VSS.n5241 VSS.n5240 0.0732424
R5946 VSS.n5236 VSS.n5241 2.21488
R5947 VSS.n5250 VSS.n5251 4.5005
R5948 VSS.n5253 VSS.n5252 0.0732424
R5949 VSS.n5251 VSS.n5253 2.21488
R5950 VSS.n5256 VSS.n5255 0.0732424
R5951 VSS.n5251 VSS.n5256 2.21488
R5952 VSS.n5265 VSS.n5266 4.5005
R5953 VSS.n5268 VSS.n5267 0.0732424
R5954 VSS.n5266 VSS.n5268 2.21488
R5955 VSS.n5271 VSS.n5270 0.0732424
R5956 VSS.n5266 VSS.n5271 2.21488
R5957 VSS.n5280 VSS.n5281 4.5005
R5958 VSS.n5282 VSS.n5283 0.0732424
R5959 VSS.n5283 VSS.n5281 2.21488
R5960 VSS.n5285 VSS.n5286 0.0732424
R5961 VSS.n5286 VSS.n5281 2.21488
R5962 VSS.n5295 VSS.n5296 4.5005
R5963 VSS.n5298 VSS.n5297 0.0732424
R5964 VSS.n5296 VSS.n5298 2.21488
R5965 VSS.n5301 VSS.n5300 0.0732424
R5966 VSS.n5296 VSS.n5301 2.21488
R5967 VSS.n5310 VSS.n5311 4.5005
R5968 VSS.n5313 VSS.n5312 0.0732424
R5969 VSS.n5311 VSS.n5313 2.21488
R5970 VSS.n5316 VSS.n5315 0.0732424
R5971 VSS.n5311 VSS.n5316 2.21488
R5972 VSS.n5325 VSS.n5326 4.5005
R5973 VSS.n5328 VSS.n5327 0.0732424
R5974 VSS.n5326 VSS.n5328 2.21488
R5975 VSS.n5331 VSS.n5330 0.0732424
R5976 VSS.n5326 VSS.n5331 2.21488
R5977 VSS.n5340 VSS.n5341 4.5005
R5978 VSS.n5342 VSS.n5343 0.0732424
R5979 VSS.n5343 VSS.n5341 2.21488
R5980 VSS.n5345 VSS.n5346 0.0732424
R5981 VSS.n5346 VSS.n5341 2.21488
R5982 VSS.n5355 VSS.n5356 4.5005
R5983 VSS.n5358 VSS.n5357 0.0732424
R5984 VSS.n5356 VSS.n5358 2.21488
R5985 VSS.n5361 VSS.n5360 0.0732424
R5986 VSS.n5356 VSS.n5361 2.21488
R5987 VSS.n5370 VSS.n5371 4.5005
R5988 VSS.n5373 VSS.n5372 0.0732424
R5989 VSS.n5371 VSS.n5373 2.21488
R5990 VSS.n5376 VSS.n5375 0.0732424
R5991 VSS.n5371 VSS.n5376 2.21488
R5992 VSS.n5385 VSS.n5386 4.5005
R5993 VSS.n5388 VSS.n5387 0.0732424
R5994 VSS.n5386 VSS.n5388 2.21488
R5995 VSS.n5391 VSS.n5390 0.0732424
R5996 VSS.n5386 VSS.n5391 2.21488
R5997 VSS.n5400 VSS.n5401 4.5005
R5998 VSS.n5403 VSS.n5402 0.0732424
R5999 VSS.n5401 VSS.n5403 2.21488
R6000 VSS.n5406 VSS.n5405 0.0732424
R6001 VSS.n5401 VSS.n5406 2.21488
R6002 VSS.n5415 VSS.n5416 4.5005
R6003 VSS.n5417 VSS.n5418 0.0732424
R6004 VSS.n5418 VSS.n5416 2.21488
R6005 VSS.n5420 VSS.n5421 0.0732424
R6006 VSS.n5421 VSS.n5416 2.21488
R6007 VSS.n5430 VSS.n5431 4.5005
R6008 VSS.n5433 VSS.n5432 0.0732424
R6009 VSS.n5431 VSS.n5433 2.21488
R6010 VSS.n5436 VSS.n5435 0.0732424
R6011 VSS.n5431 VSS.n5436 2.21488
R6012 VSS.n5445 VSS.n5446 4.5005
R6013 VSS.n5448 VSS.n5447 0.0732424
R6014 VSS.n5446 VSS.n5448 2.21488
R6015 VSS.n5451 VSS.n5450 0.0732424
R6016 VSS.n5446 VSS.n5451 2.21488
R6017 VSS.n5460 VSS.n5461 4.5005
R6018 VSS.n5463 VSS.n5462 0.0732424
R6019 VSS.n5461 VSS.n5463 2.21488
R6020 VSS.n5466 VSS.n5465 0.0732424
R6021 VSS.n5461 VSS.n5466 2.21488
R6022 VSS.n5475 VSS.n5476 4.5005
R6023 VSS.n5477 VSS.n5478 0.0732424
R6024 VSS.n5478 VSS.n5476 2.21488
R6025 VSS.n5480 VSS.n5481 0.0732424
R6026 VSS.n5481 VSS.n5476 2.21488
R6027 VSS.n5490 VSS.n5491 4.5005
R6028 VSS.n5493 VSS.n5492 0.0732424
R6029 VSS.n5491 VSS.n5493 2.21488
R6030 VSS.n5496 VSS.n5495 0.0732424
R6031 VSS.n5491 VSS.n5496 2.21488
R6032 VSS.n5505 VSS.n5506 4.5005
R6033 VSS.n5508 VSS.n5507 0.0732424
R6034 VSS.n5506 VSS.n5508 2.21488
R6035 VSS.n5511 VSS.n5510 0.0732424
R6036 VSS.n5506 VSS.n5511 2.21488
R6037 VSS.n5520 VSS.n5521 4.5005
R6038 VSS.n5523 VSS.n5522 0.0732424
R6039 VSS.n5521 VSS.n5523 2.21488
R6040 VSS.n5526 VSS.n5525 0.0732424
R6041 VSS.n5521 VSS.n5526 2.21488
R6042 VSS.n5535 VSS.n5536 4.5005
R6043 VSS.n5538 VSS.n5537 0.0732424
R6044 VSS.n5536 VSS.n5538 2.21488
R6045 VSS.n5541 VSS.n5540 0.0732424
R6046 VSS.n5536 VSS.n5541 2.21488
R6047 VSS.n5550 VSS.n5551 4.5005
R6048 VSS.n5553 VSS.n5552 0.0732424
R6049 VSS.n5551 VSS.n5553 2.21488
R6050 VSS.n5556 VSS.n5555 0.0732424
R6051 VSS.n5551 VSS.n5556 2.21488
R6052 VSS.n5565 VSS.n5566 4.5005
R6053 VSS.n5568 VSS.n5567 0.0732424
R6054 VSS.n5566 VSS.n5568 2.21488
R6055 VSS.n5571 VSS.n5570 0.0732424
R6056 VSS.n5566 VSS.n5571 2.21488
R6057 VSS.n5580 VSS.n5581 4.5005
R6058 VSS.n5582 VSS.n5583 0.0732424
R6059 VSS.n5583 VSS.n5581 2.21488
R6060 VSS.n5585 VSS.n5586 0.0732424
R6061 VSS.n5586 VSS.n5581 2.21488
R6062 VSS.n5595 VSS.n5596 4.5005
R6063 VSS.n5598 VSS.n5597 0.0732424
R6064 VSS.n5596 VSS.n5598 2.21488
R6065 VSS.n5601 VSS.n5600 0.0732424
R6066 VSS.n5596 VSS.n5601 2.21488
R6067 VSS.n5610 VSS.n5611 4.5005
R6068 VSS.n5613 VSS.n5612 0.0732424
R6069 VSS.n5611 VSS.n5613 2.21488
R6070 VSS.n5616 VSS.n5615 0.0732424
R6071 VSS.n5611 VSS.n5616 2.21488
R6072 VSS.n5625 VSS.n5626 4.5005
R6073 VSS.n5628 VSS.n5627 0.0732424
R6074 VSS.n5626 VSS.n5628 2.21488
R6075 VSS.n5631 VSS.n5630 0.0732424
R6076 VSS.n5626 VSS.n5631 2.21488
R6077 VSS.n5640 VSS.n5641 4.5005
R6078 VSS.n5642 VSS.n5643 0.0732424
R6079 VSS.n5643 VSS.n5641 2.21488
R6080 VSS.n5645 VSS.n5646 0.0732424
R6081 VSS.n5646 VSS.n5641 2.21488
R6082 VSS.n5655 VSS.n5656 4.5005
R6083 VSS.n5658 VSS.n5657 0.0732424
R6084 VSS.n5656 VSS.n5658 2.21488
R6085 VSS.n5661 VSS.n5660 0.0732424
R6086 VSS.n5656 VSS.n5661 2.21488
R6087 VSS.n5670 VSS.n5671 4.5005
R6088 VSS.n5673 VSS.n5672 0.0732424
R6089 VSS.n5671 VSS.n5673 2.21488
R6090 VSS.n5676 VSS.n5675 0.0732424
R6091 VSS.n5671 VSS.n5676 2.21488
R6092 VSS.n5685 VSS.n5686 4.5005
R6093 VSS.n5688 VSS.n5687 0.0732424
R6094 VSS.n5686 VSS.n5688 2.21488
R6095 VSS.n5691 VSS.n5690 0.0732424
R6096 VSS.n5686 VSS.n5691 2.21488
R6097 VSS.n5700 VSS.n5701 4.5005
R6098 VSS.n5703 VSS.n5702 0.0732424
R6099 VSS.n5701 VSS.n5703 2.21488
R6100 VSS.n5706 VSS.n5705 0.0732424
R6101 VSS.n5701 VSS.n5706 2.21488
R6102 VSS.n5715 VSS.n5716 4.5005
R6103 VSS.n5717 VSS.n5718 0.0732424
R6104 VSS.n5718 VSS.n5716 2.21488
R6105 VSS.n5720 VSS.n5721 0.0732424
R6106 VSS.n5721 VSS.n5716 2.21488
R6107 VSS.n5730 VSS.n5731 4.5005
R6108 VSS.n5733 VSS.n5732 0.0732424
R6109 VSS.n5731 VSS.n5733 2.21488
R6110 VSS.n5736 VSS.n5735 0.0732424
R6111 VSS.n5731 VSS.n5736 2.21488
R6112 VSS.n5745 VSS.n5746 4.5005
R6113 VSS.n5748 VSS.n5747 0.0732424
R6114 VSS.n5746 VSS.n5748 2.21488
R6115 VSS.n5751 VSS.n5750 0.0732424
R6116 VSS.n5746 VSS.n5751 2.21488
R6117 VSS.n5760 VSS.n5761 4.5005
R6118 VSS.n5763 VSS.n5762 0.0732424
R6119 VSS.n5761 VSS.n5763 2.21488
R6120 VSS.n5766 VSS.n5765 0.0732424
R6121 VSS.n5761 VSS.n5766 2.21488
R6122 VSS.n5775 VSS.n5776 4.5005
R6123 VSS.n5777 VSS.n5778 0.0732424
R6124 VSS.n5778 VSS.n5776 2.21488
R6125 VSS.n5780 VSS.n5781 0.0732424
R6126 VSS.n5781 VSS.n5776 2.21488
R6127 VSS.n5790 VSS.n5791 4.5005
R6128 VSS.n5793 VSS.n5792 0.0732424
R6129 VSS.n5791 VSS.n5793 2.21488
R6130 VSS.n5796 VSS.n5795 0.0732424
R6131 VSS.n5791 VSS.n5796 2.21488
R6132 VSS.n5805 VSS.n5806 4.5005
R6133 VSS.n5808 VSS.n5807 0.0732424
R6134 VSS.n5806 VSS.n5808 2.21488
R6135 VSS.n5811 VSS.n5810 0.0732424
R6136 VSS.n5806 VSS.n5811 2.21488
R6137 VSS.n5820 VSS.n5821 4.5005
R6138 VSS.n5823 VSS.n5822 0.0732424
R6139 VSS.n5821 VSS.n5823 2.21488
R6140 VSS.n5826 VSS.n5825 0.0732424
R6141 VSS.n5821 VSS.n5826 2.21488
R6142 VSS.n5835 VSS.n5836 4.5005
R6143 VSS.n5838 VSS.n5837 0.0732424
R6144 VSS.n5836 VSS.n5838 2.21488
R6145 VSS.n5841 VSS.n5840 0.0732424
R6146 VSS.n5836 VSS.n5841 2.21488
R6147 VSS.n5850 VSS.n5851 4.5005
R6148 VSS.n5853 VSS.n5852 0.0732424
R6149 VSS.n5851 VSS.n5853 2.21488
R6150 VSS.n5856 VSS.n5855 0.0732424
R6151 VSS.n5851 VSS.n5856 2.21488
R6152 VSS.n5865 VSS.n5866 4.5005
R6153 VSS.n5868 VSS.n5867 0.0732424
R6154 VSS.n5866 VSS.n5868 2.21488
R6155 VSS.n5871 VSS.n5870 0.0732424
R6156 VSS.n5866 VSS.n5871 2.21488
R6157 VSS.n5880 VSS.n5881 4.5005
R6158 VSS.n5882 VSS.n5883 0.0732424
R6159 VSS.n5883 VSS.n5881 2.21488
R6160 VSS.n5885 VSS.n5886 0.0732424
R6161 VSS.n5886 VSS.n5881 2.21488
R6162 VSS.n5895 VSS.n5896 4.5005
R6163 VSS.n5898 VSS.n5897 0.0732424
R6164 VSS.n5896 VSS.n5898 2.21488
R6165 VSS.n5901 VSS.n5900 0.0732424
R6166 VSS.n5896 VSS.n5901 2.21488
R6167 VSS.n5910 VSS.n5911 4.5005
R6168 VSS.n5913 VSS.n5912 0.0732424
R6169 VSS.n5911 VSS.n5913 2.21488
R6170 VSS.n5916 VSS.n5915 0.0732424
R6171 VSS.n5911 VSS.n5916 2.21488
R6172 VSS.n5925 VSS.n5926 4.5005
R6173 VSS.n5928 VSS.n5927 0.0732424
R6174 VSS.n5926 VSS.n5928 2.21488
R6175 VSS.n5931 VSS.n5930 0.0732424
R6176 VSS.n5926 VSS.n5931 2.21488
R6177 VSS.n5940 VSS.n5941 4.5005
R6178 VSS.n5942 VSS.n5943 0.0732424
R6179 VSS.n5943 VSS.n5941 2.21488
R6180 VSS.n5945 VSS.n5946 0.0732424
R6181 VSS.n5946 VSS.n5941 2.21488
R6182 VSS.n5955 VSS.n5956 4.5005
R6183 VSS.n5958 VSS.n5957 0.0732424
R6184 VSS.n5956 VSS.n5958 2.21488
R6185 VSS.n5961 VSS.n5960 0.0732424
R6186 VSS.n5956 VSS.n5961 2.21488
R6187 VSS.n5970 VSS.n5971 4.5005
R6188 VSS.n5973 VSS.n5972 0.0732424
R6189 VSS.n5971 VSS.n5973 2.21488
R6190 VSS.n5976 VSS.n5975 0.0732424
R6191 VSS.n5971 VSS.n5976 2.21488
R6192 VSS.n5985 VSS.n5986 4.5005
R6193 VSS.n5988 VSS.n5987 0.0732424
R6194 VSS.n5986 VSS.n5988 2.21488
R6195 VSS.n5991 VSS.n5990 0.0732424
R6196 VSS.n5986 VSS.n5991 2.21488
R6197 VSS.n6000 VSS.n6001 4.5005
R6198 VSS.n6003 VSS.n6002 0.0732424
R6199 VSS.n6001 VSS.n6003 2.21488
R6200 VSS.n6006 VSS.n6005 0.0732424
R6201 VSS.n6001 VSS.n6006 2.21488
R6202 VSS.n6015 VSS.n6016 4.5005
R6203 VSS.n6017 VSS.n6018 0.0732424
R6204 VSS.n6018 VSS.n6016 2.21488
R6205 VSS.n6020 VSS.n6021 0.0732424
R6206 VSS.n6021 VSS.n6016 2.21488
R6207 VSS.n6030 VSS.n6031 4.5005
R6208 VSS.n6033 VSS.n6032 0.0732424
R6209 VSS.n6031 VSS.n6033 2.21488
R6210 VSS.n6036 VSS.n6035 0.0732424
R6211 VSS.n6031 VSS.n6036 2.21488
R6212 VSS.n6045 VSS.n6046 4.5005
R6213 VSS.n6048 VSS.n6047 0.0732424
R6214 VSS.n6046 VSS.n6048 2.21488
R6215 VSS.n6051 VSS.n6050 0.0732424
R6216 VSS.n6046 VSS.n6051 2.21488
R6217 VSS.n6060 VSS.n6061 4.5005
R6218 VSS.n6063 VSS.n6062 0.0732424
R6219 VSS.n6061 VSS.n6063 2.21488
R6220 VSS.n6066 VSS.n6065 0.0732424
R6221 VSS.n6061 VSS.n6066 2.21488
R6222 VSS.n6075 VSS.n6076 4.5005
R6223 VSS.n6077 VSS.n6078 0.0732424
R6224 VSS.n6078 VSS.n6076 2.21488
R6225 VSS.n6080 VSS.n6081 0.0732424
R6226 VSS.n6081 VSS.n6076 2.21488
R6227 VSS.n6090 VSS.n6091 4.5005
R6228 VSS.n6093 VSS.n6092 0.0732424
R6229 VSS.n6091 VSS.n6093 2.21488
R6230 VSS.n6096 VSS.n6095 0.0732424
R6231 VSS.n6091 VSS.n6096 2.21488
R6232 VSS.n6105 VSS.n6106 4.5005
R6233 VSS.n6108 VSS.n6107 0.0732424
R6234 VSS.n6106 VSS.n6108 2.21488
R6235 VSS.n6111 VSS.n6110 0.0732424
R6236 VSS.n6106 VSS.n6111 2.21488
R6237 VSS.n6120 VSS.n6121 4.5005
R6238 VSS.n6123 VSS.n6122 0.0732424
R6239 VSS.n6121 VSS.n6123 2.21488
R6240 VSS.n6126 VSS.n6125 0.0732424
R6241 VSS.n6121 VSS.n6126 2.21488
R6242 VSS.n6135 VSS.n6136 4.5005
R6243 VSS.n6138 VSS.n6137 0.0732424
R6244 VSS.n6136 VSS.n6138 2.21488
R6245 VSS.n6141 VSS.n6140 0.0732424
R6246 VSS.n6136 VSS.n6141 2.21488
R6247 VSS.n6150 VSS.n6151 4.5005
R6248 VSS.n6153 VSS.n6152 0.0732424
R6249 VSS.n6151 VSS.n6153 2.21488
R6250 VSS.n6156 VSS.n6155 0.0732424
R6251 VSS.n6151 VSS.n6156 2.21488
R6252 VSS.n6165 VSS.n6166 4.5005
R6253 VSS.n6168 VSS.n6167 0.0732424
R6254 VSS.n6166 VSS.n6168 2.21488
R6255 VSS.n6171 VSS.n6170 0.0732424
R6256 VSS.n6166 VSS.n6171 2.21488
R6257 VSS.n6180 VSS.n6181 4.5005
R6258 VSS.n6182 VSS.n6183 0.0732424
R6259 VSS.n6183 VSS.n6181 2.21488
R6260 VSS.n6185 VSS.n6186 0.0732424
R6261 VSS.n6186 VSS.n6181 2.21488
R6262 VSS.n6195 VSS.n6196 4.5005
R6263 VSS.n6198 VSS.n6197 0.0732424
R6264 VSS.n6196 VSS.n6198 2.21488
R6265 VSS.n6201 VSS.n6200 0.0732424
R6266 VSS.n6196 VSS.n6201 2.21488
R6267 VSS.n6210 VSS.n6211 4.5005
R6268 VSS.n6213 VSS.n6212 0.0732424
R6269 VSS.n6211 VSS.n6213 2.21488
R6270 VSS.n6216 VSS.n6215 0.0732424
R6271 VSS.n6211 VSS.n6216 2.21488
R6272 VSS.n6225 VSS.n6226 4.5005
R6273 VSS.n6228 VSS.n6227 0.0732424
R6274 VSS.n6226 VSS.n6228 2.21488
R6275 VSS.n6231 VSS.n6230 0.0732424
R6276 VSS.n6226 VSS.n6231 2.21488
R6277 VSS.n6240 VSS.n6241 4.5005
R6278 VSS.n6242 VSS.n6243 0.0732424
R6279 VSS.n6243 VSS.n6241 2.21488
R6280 VSS.n6245 VSS.n6246 0.0732424
R6281 VSS.n6246 VSS.n6241 2.21488
R6282 VSS.n6255 VSS.n6256 4.5005
R6283 VSS.n6258 VSS.n6257 0.0732424
R6284 VSS.n6256 VSS.n6258 2.21488
R6285 VSS.n6261 VSS.n6260 0.0732424
R6286 VSS.n6256 VSS.n6261 2.21488
R6287 VSS.n6270 VSS.n6271 4.5005
R6288 VSS.n6273 VSS.n6272 0.0732424
R6289 VSS.n6271 VSS.n6273 2.21488
R6290 VSS.n6276 VSS.n6275 0.0732424
R6291 VSS.n6271 VSS.n6276 2.21488
R6292 VSS.n6285 VSS.n6286 4.5005
R6293 VSS.n6288 VSS.n6287 0.0732424
R6294 VSS.n6286 VSS.n6288 2.21488
R6295 VSS.n6291 VSS.n6290 0.0732424
R6296 VSS.n6286 VSS.n6291 2.21488
R6297 VSS.n6300 VSS.n6301 4.5005
R6298 VSS.n6303 VSS.n6302 0.0732424
R6299 VSS.n6301 VSS.n6303 2.21488
R6300 VSS.n6306 VSS.n6305 0.0732424
R6301 VSS.n6301 VSS.n6306 2.21488
R6302 VSS.n6315 VSS.n6316 4.5005
R6303 VSS.n6317 VSS.n6318 0.0732424
R6304 VSS.n6318 VSS.n6316 2.21488
R6305 VSS.n6320 VSS.n6321 0.0732424
R6306 VSS.n6321 VSS.n6316 2.21488
R6307 VSS.n6330 VSS.n6331 4.5005
R6308 VSS.n6333 VSS.n6332 0.0732424
R6309 VSS.n6331 VSS.n6333 2.21488
R6310 VSS.n6336 VSS.n6335 0.0732424
R6311 VSS.n6331 VSS.n6336 2.21488
R6312 VSS.n6345 VSS.n6346 4.5005
R6313 VSS.n6348 VSS.n6347 0.0732424
R6314 VSS.n6346 VSS.n6348 2.21488
R6315 VSS.n6351 VSS.n6350 0.0732424
R6316 VSS.n6346 VSS.n6351 2.21488
R6317 VSS.n6360 VSS.n6361 4.5005
R6318 VSS.n6363 VSS.n6362 0.0732424
R6319 VSS.n6361 VSS.n6363 2.21488
R6320 VSS.n6366 VSS.n6365 0.0732424
R6321 VSS.n6361 VSS.n6366 2.21488
R6322 VSS.n6375 VSS.n6376 4.5005
R6323 VSS.n6377 VSS.n6378 0.0732424
R6324 VSS.n6378 VSS.n6376 2.21488
R6325 VSS.n6380 VSS.n6381 0.0732424
R6326 VSS.n6381 VSS.n6376 2.21488
R6327 VSS.n6390 VSS.n6391 4.5005
R6328 VSS.n6393 VSS.n6392 0.0732424
R6329 VSS.n6391 VSS.n6393 2.21488
R6330 VSS.n6396 VSS.n6395 0.0732424
R6331 VSS.n6391 VSS.n6396 2.21488
R6332 VSS.n6405 VSS.n6406 4.5005
R6333 VSS.n6408 VSS.n6407 0.0732424
R6334 VSS.n6406 VSS.n6408 2.21488
R6335 VSS.n6411 VSS.n6410 0.0732424
R6336 VSS.n6406 VSS.n6411 2.21488
R6337 VSS.n6420 VSS.n6421 4.5005
R6338 VSS.n6423 VSS.n6422 0.0732424
R6339 VSS.n6421 VSS.n6423 2.21488
R6340 VSS.n6426 VSS.n6425 0.0732424
R6341 VSS.n6421 VSS.n6426 2.21488
R6342 VSS.n6435 VSS.n6436 4.5005
R6343 VSS.n6438 VSS.n6437 0.0732424
R6344 VSS.n6436 VSS.n6438 2.21488
R6345 VSS.n6441 VSS.n6440 0.0732424
R6346 VSS.n6436 VSS.n6441 2.21488
R6347 VSS.n6450 VSS.n6451 4.5005
R6348 VSS.n6453 VSS.n6452 0.0732424
R6349 VSS.n6451 VSS.n6453 2.21488
R6350 VSS.n6456 VSS.n6455 0.0732424
R6351 VSS.n6451 VSS.n6456 2.21488
R6352 VSS.n6465 VSS.n6466 4.5005
R6353 VSS.n6468 VSS.n6467 0.0732424
R6354 VSS.n6466 VSS.n6468 2.21488
R6355 VSS.n6471 VSS.n6470 0.0732424
R6356 VSS.n6466 VSS.n6471 2.21488
R6357 VSS.n6480 VSS.n6481 4.5005
R6358 VSS.n6482 VSS.n6483 0.0732424
R6359 VSS.n6483 VSS.n6481 2.21488
R6360 VSS.n6485 VSS.n6486 0.0732424
R6361 VSS.n6486 VSS.n6481 2.21488
R6362 VSS.n6495 VSS.n6496 4.5005
R6363 VSS.n6498 VSS.n6497 0.0732424
R6364 VSS.n6496 VSS.n6498 2.21488
R6365 VSS.n6501 VSS.n6500 0.0732424
R6366 VSS.n6496 VSS.n6501 2.21488
R6367 VSS.n6510 VSS.n6511 4.5005
R6368 VSS.n6513 VSS.n6512 0.0732424
R6369 VSS.n6511 VSS.n6513 2.21488
R6370 VSS.n6516 VSS.n6515 0.0732424
R6371 VSS.n6511 VSS.n6516 2.21488
R6372 VSS.n6525 VSS.n6526 4.5005
R6373 VSS.n6528 VSS.n6527 0.0732424
R6374 VSS.n6526 VSS.n6528 2.21488
R6375 VSS.n6531 VSS.n6530 0.0732424
R6376 VSS.n6526 VSS.n6531 2.21488
R6377 VSS.n6540 VSS.n6541 4.5005
R6378 VSS.n6542 VSS.n6543 0.0732424
R6379 VSS.n6543 VSS.n6541 2.21488
R6380 VSS.n6545 VSS.n6546 0.0732424
R6381 VSS.n6546 VSS.n6541 2.21488
R6382 VSS.n6555 VSS.n6556 4.5005
R6383 VSS.n6558 VSS.n6557 0.0732424
R6384 VSS.n6556 VSS.n6558 2.21488
R6385 VSS.n6561 VSS.n6560 0.0732424
R6386 VSS.n6556 VSS.n6561 2.21488
R6387 VSS.n6570 VSS.n6571 4.5005
R6388 VSS.n6573 VSS.n6572 0.0732424
R6389 VSS.n6571 VSS.n6573 2.21488
R6390 VSS.n6576 VSS.n6575 0.0732424
R6391 VSS.n6571 VSS.n6576 2.21488
R6392 VSS.n6585 VSS.n6586 4.5005
R6393 VSS.n6588 VSS.n6587 0.0732424
R6394 VSS.n6586 VSS.n6588 2.21488
R6395 VSS.n6591 VSS.n6590 0.0732424
R6396 VSS.n6586 VSS.n6591 2.21488
R6397 VSS.n6600 VSS.n6601 4.5005
R6398 VSS.n6603 VSS.n6602 0.0732424
R6399 VSS.n6601 VSS.n6603 2.21488
R6400 VSS.n6606 VSS.n6605 0.0732424
R6401 VSS.n6601 VSS.n6606 2.21488
R6402 VSS.n6615 VSS.n6616 4.5005
R6403 VSS.n6617 VSS.n6618 0.0732424
R6404 VSS.n6618 VSS.n6616 2.21488
R6405 VSS.n6620 VSS.n6621 0.0732424
R6406 VSS.n6621 VSS.n6616 2.21488
R6407 VSS.n6630 VSS.n6631 4.5005
R6408 VSS.n6633 VSS.n6632 0.0732424
R6409 VSS.n6631 VSS.n6633 2.21488
R6410 VSS.n6636 VSS.n6635 0.0732424
R6411 VSS.n6631 VSS.n6636 2.21488
R6412 VSS.n6645 VSS.n6646 4.5005
R6413 VSS.n6648 VSS.n6647 0.0732424
R6414 VSS.n6646 VSS.n6648 2.21488
R6415 VSS.n6651 VSS.n6650 0.0732424
R6416 VSS.n6646 VSS.n6651 2.21488
R6417 VSS.n6660 VSS.n6661 4.5005
R6418 VSS.n6663 VSS.n6662 0.0732424
R6419 VSS.n6661 VSS.n6663 2.21488
R6420 VSS.n6666 VSS.n6665 0.0732424
R6421 VSS.n6661 VSS.n6666 2.21488
R6422 VSS.n6675 VSS.n6676 4.5005
R6423 VSS.n6677 VSS.n6678 0.0732424
R6424 VSS.n6678 VSS.n6676 2.21488
R6425 VSS.n6680 VSS.n6681 0.0732424
R6426 VSS.n6681 VSS.n6676 2.21488
R6427 VSS.n6690 VSS.n6691 4.5005
R6428 VSS.n6693 VSS.n6692 0.0732424
R6429 VSS.n6691 VSS.n6693 2.21488
R6430 VSS.n6696 VSS.n6695 0.0732424
R6431 VSS.n6691 VSS.n6696 2.21488
R6432 VSS.n6705 VSS.n6706 4.5005
R6433 VSS.n6708 VSS.n6707 0.0732424
R6434 VSS.n6706 VSS.n6708 2.21488
R6435 VSS.n6711 VSS.n6710 0.0732424
R6436 VSS.n6706 VSS.n6711 2.21488
R6437 VSS.n6720 VSS.n6721 4.5005
R6438 VSS.n6723 VSS.n6722 0.0732424
R6439 VSS.n6721 VSS.n6723 2.21488
R6440 VSS.n6726 VSS.n6725 0.0732424
R6441 VSS.n6721 VSS.n6726 2.21488
R6442 VSS.n6735 VSS.n6736 4.5005
R6443 VSS.n6738 VSS.n6737 0.0732424
R6444 VSS.n6736 VSS.n6738 2.21488
R6445 VSS.n6741 VSS.n6740 0.0732424
R6446 VSS.n6736 VSS.n6741 2.21488
R6447 VSS.n6750 VSS.n6751 4.5005
R6448 VSS.n6753 VSS.n6752 0.0732424
R6449 VSS.n6751 VSS.n6753 2.21488
R6450 VSS.n6756 VSS.n6755 0.0732424
R6451 VSS.n6751 VSS.n6756 2.21488
R6452 VSS.n6765 VSS.n6766 4.5005
R6453 VSS.n6768 VSS.n6767 0.0732424
R6454 VSS.n6766 VSS.n6768 2.21488
R6455 VSS.n6771 VSS.n6770 0.0732424
R6456 VSS.n6766 VSS.n6771 2.21488
R6457 VSS.n6780 VSS.n6781 4.5005
R6458 VSS.n6782 VSS.n6783 0.0732424
R6459 VSS.n6783 VSS.n6781 2.21488
R6460 VSS.n6785 VSS.n6786 0.0732424
R6461 VSS.n6786 VSS.n6781 2.21488
R6462 VSS.n6795 VSS.n6796 4.5005
R6463 VSS.n6798 VSS.n6797 0.0732424
R6464 VSS.n6796 VSS.n6798 2.21488
R6465 VSS.n6801 VSS.n6800 0.0732424
R6466 VSS.n6796 VSS.n6801 2.21488
R6467 VSS.n6810 VSS.n6811 4.5005
R6468 VSS.n6813 VSS.n6812 0.0732424
R6469 VSS.n6811 VSS.n6813 2.21488
R6470 VSS.n6816 VSS.n6815 0.0732424
R6471 VSS.n6811 VSS.n6816 2.21488
R6472 VSS.n6825 VSS.n6826 4.5005
R6473 VSS.n6828 VSS.n6827 0.0732424
R6474 VSS.n6826 VSS.n6828 2.21488
R6475 VSS.n6831 VSS.n6830 0.0732424
R6476 VSS.n6826 VSS.n6831 2.21488
R6477 VSS.n6840 VSS.n6841 4.5005
R6478 VSS.n6842 VSS.n6843 0.0732424
R6479 VSS.n6843 VSS.n6841 2.21488
R6480 VSS.n6845 VSS.n6846 0.0732424
R6481 VSS.n6846 VSS.n6841 2.21488
R6482 VSS.n6855 VSS.n6856 4.5005
R6483 VSS.n6858 VSS.n6857 0.0732424
R6484 VSS.n6856 VSS.n6858 2.21488
R6485 VSS.n6861 VSS.n6860 0.0732424
R6486 VSS.n6856 VSS.n6861 2.21488
R6487 VSS.n6870 VSS.n6871 4.5005
R6488 VSS.n6873 VSS.n6872 0.0732424
R6489 VSS.n6871 VSS.n6873 2.21488
R6490 VSS.n6876 VSS.n6875 0.0732424
R6491 VSS.n6871 VSS.n6876 2.21488
R6492 VSS.n6885 VSS.n6886 4.5005
R6493 VSS.n6888 VSS.n6887 0.0732424
R6494 VSS.n6886 VSS.n6888 2.21488
R6495 VSS.n6891 VSS.n6890 0.0732424
R6496 VSS.n6886 VSS.n6891 2.21488
R6497 VSS.n6900 VSS.n6901 4.5005
R6498 VSS.n6903 VSS.n6902 0.0732424
R6499 VSS.n6901 VSS.n6903 2.21488
R6500 VSS.n6906 VSS.n6905 0.0732424
R6501 VSS.n6901 VSS.n6906 2.21488
R6502 VSS.n6915 VSS.n6916 4.5005
R6503 VSS.n6917 VSS.n6918 0.0732424
R6504 VSS.n6918 VSS.n6916 2.21488
R6505 VSS.n6920 VSS.n6921 0.0732424
R6506 VSS.n6921 VSS.n6916 2.21488
R6507 VSS.n6930 VSS.n6931 4.5005
R6508 VSS.n6933 VSS.n6932 0.0732424
R6509 VSS.n6931 VSS.n6933 2.21488
R6510 VSS.n6936 VSS.n6935 0.0732424
R6511 VSS.n6931 VSS.n6936 2.21488
R6512 VSS.n6945 VSS.n6946 4.5005
R6513 VSS.n6948 VSS.n6947 0.0732424
R6514 VSS.n6946 VSS.n6948 2.21488
R6515 VSS.n6951 VSS.n6950 0.0732424
R6516 VSS.n6946 VSS.n6951 2.21488
R6517 VSS.n6960 VSS.n6961 4.5005
R6518 VSS.n6963 VSS.n6962 0.0732424
R6519 VSS.n6961 VSS.n6963 2.21488
R6520 VSS.n6966 VSS.n6965 0.0732424
R6521 VSS.n6961 VSS.n6966 2.21488
R6522 VSS.n6975 VSS.n6976 4.5005
R6523 VSS.n6977 VSS.n6978 0.0732424
R6524 VSS.n6978 VSS.n6976 2.21488
R6525 VSS.n6980 VSS.n6981 0.0732424
R6526 VSS.n6981 VSS.n6976 2.21488
R6527 VSS.n6990 VSS.n6991 4.5005
R6528 VSS.n6993 VSS.n6992 0.0732424
R6529 VSS.n6991 VSS.n6993 2.21488
R6530 VSS.n6996 VSS.n6995 0.0732424
R6531 VSS.n6991 VSS.n6996 2.21488
R6532 VSS.n7005 VSS.n7006 4.5005
R6533 VSS.n7008 VSS.n7007 0.0732424
R6534 VSS.n7006 VSS.n7008 2.21488
R6535 VSS.n7011 VSS.n7010 0.0732424
R6536 VSS.n7006 VSS.n7011 2.21488
R6537 VSS.n7020 VSS.n7021 4.5005
R6538 VSS.n7023 VSS.n7022 0.0732424
R6539 VSS.n7021 VSS.n7023 2.21488
R6540 VSS.n7026 VSS.n7025 0.0732424
R6541 VSS.n7021 VSS.n7026 2.21488
R6542 VSS.n7035 VSS.n7036 4.5005
R6543 VSS.n7038 VSS.n7037 0.0732424
R6544 VSS.n7036 VSS.n7038 2.21488
R6545 VSS.n7041 VSS.n7040 0.0732424
R6546 VSS.n7036 VSS.n7041 2.21488
R6547 VSS.n7050 VSS.n7051 4.5005
R6548 VSS.n7053 VSS.n7052 0.0732424
R6549 VSS.n7051 VSS.n7053 2.21488
R6550 VSS.n7056 VSS.n7055 0.0732424
R6551 VSS.n7051 VSS.n7056 2.21488
R6552 VSS.n7065 VSS.n7066 4.5005
R6553 VSS.n7068 VSS.n7067 0.0732424
R6554 VSS.n7066 VSS.n7068 2.21488
R6555 VSS.n7071 VSS.n7070 0.0732424
R6556 VSS.n7066 VSS.n7071 2.21488
R6557 VSS.n7080 VSS.n7081 4.5005
R6558 VSS.n7082 VSS.n7083 0.0732424
R6559 VSS.n7083 VSS.n7081 2.21488
R6560 VSS.n7085 VSS.n7086 0.0732424
R6561 VSS.n7086 VSS.n7081 2.21488
R6562 VSS.n7095 VSS.n7096 4.5005
R6563 VSS.n7098 VSS.n7097 0.0732424
R6564 VSS.n7096 VSS.n7098 2.21488
R6565 VSS.n7101 VSS.n7100 0.0732424
R6566 VSS.n7096 VSS.n7101 2.21488
R6567 VSS.n7110 VSS.n7111 4.5005
R6568 VSS.n7113 VSS.n7112 0.0732424
R6569 VSS.n7111 VSS.n7113 2.21488
R6570 VSS.n7116 VSS.n7115 0.0732424
R6571 VSS.n7111 VSS.n7116 2.21488
R6572 VSS.n7125 VSS.n7126 4.5005
R6573 VSS.n7128 VSS.n7127 0.0732424
R6574 VSS.n7126 VSS.n7128 2.21488
R6575 VSS.n7131 VSS.n7130 0.0732424
R6576 VSS.n7126 VSS.n7131 2.21488
R6577 VSS.n7140 VSS.n7141 4.5005
R6578 VSS.n7143 VSS.n7142 0.0732424
R6579 VSS.n7141 VSS.n7143 2.21488
R6580 VSS.n7146 VSS.n7145 0.0732424
R6581 VSS.n7141 VSS.n7146 2.21488
R6582 VSS.n7155 VSS.n7156 4.5005
R6583 VSS.n7158 VSS.n7157 0.0732424
R6584 VSS.n7156 VSS.n7158 2.21488
R6585 VSS.n7161 VSS.n7160 0.0732424
R6586 VSS.n7156 VSS.n7161 2.21488
R6587 VSS.n7141 VSS.n7156 0.0584021
R6588 VSS.n4784 VSS.n7141 0.0596608
R6589 VSS.n4784 VSS.n7126 0.0244161
R6590 VSS.n7126 VSS.n7111 0.0585594
R6591 VSS.n7111 VSS.n7096 0.0584021
R6592 VSS.n7081 VSS.n7096 0.0596608
R6593 VSS.n7081 VSS.n7066 0.0244161
R6594 VSS.n7066 VSS.n7051 0.0585594
R6595 VSS.n7051 VSS.n7036 0.0584021
R6596 VSS.n7036 VSS 0.16272
R6597 VSS VSS.n7021 0.143052
R6598 VSS.n7006 VSS.n7021 0.0584021
R6599 VSS.n6991 VSS.n7006 0.0584021
R6600 VSS.n6976 VSS.n6991 0.0244161
R6601 VSS.n6976 VSS.n6961 0.0598182
R6602 VSS.n6961 VSS.n6946 0.0584021
R6603 VSS.n6931 VSS.n6946 0.0584021
R6604 VSS.n6916 VSS.n6931 0.0244161
R6605 VSS.n6916 VSS.n6901 0.0598182
R6606 VSS.n6901 VSS.n6886 0.0584021
R6607 VSS.n6886 VSS.n6871 0.0231573
R6608 VSS.n6856 VSS.n6871 0.0584021
R6609 VSS.n6841 VSS.n6856 0.0596608
R6610 VSS.n6841 VSS.n6826 0.0244161
R6611 VSS.n6826 VSS.n6811 0.0585594
R6612 VSS.n6811 VSS.n6796 0.0584021
R6613 VSS.n6781 VSS.n6796 0.0596608
R6614 VSS.n6781 VSS.n6766 0.0244161
R6615 VSS.n6766 VSS.n6751 0.0585594
R6616 VSS.n6751 VSS.n6736 0.0584021
R6617 VSS.n6736 VSS 0.16272
R6618 VSS VSS.n6721 0.143052
R6619 VSS.n6706 VSS.n6721 0.0584021
R6620 VSS.n6691 VSS.n6706 0.0584021
R6621 VSS.n6676 VSS.n6691 0.0244161
R6622 VSS.n6676 VSS.n6661 0.0598182
R6623 VSS.n6661 VSS.n6646 0.0584021
R6624 VSS.n6631 VSS.n6646 0.0584021
R6625 VSS.n6616 VSS.n6631 0.0244161
R6626 VSS.n6616 VSS.n6601 0.0598182
R6627 VSS.n6601 VSS.n6586 0.0584021
R6628 VSS.n6586 VSS.n6571 0.0231573
R6629 VSS.n6556 VSS.n6571 0.0584021
R6630 VSS.n6541 VSS.n6556 0.0596608
R6631 VSS.n6541 VSS.n6526 0.0244161
R6632 VSS.n6526 VSS.n6511 0.0585594
R6633 VSS.n6511 VSS.n6496 0.0584021
R6634 VSS.n6481 VSS.n6496 0.0596608
R6635 VSS.n6481 VSS.n6466 0.0244161
R6636 VSS.n6466 VSS.n6451 0.0585594
R6637 VSS.n6451 VSS.n6436 0.0584021
R6638 VSS.n6436 VSS 0.16272
R6639 VSS VSS.n6421 0.143052
R6640 VSS.n6406 VSS.n6421 0.0584021
R6641 VSS.n6391 VSS.n6406 0.0584021
R6642 VSS.n6376 VSS.n6391 0.0244161
R6643 VSS.n6376 VSS.n6361 0.0598182
R6644 VSS.n6361 VSS.n6346 0.0584021
R6645 VSS.n6331 VSS.n6346 0.0584021
R6646 VSS.n6316 VSS.n6331 0.0244161
R6647 VSS.n6316 VSS.n6301 0.0598182
R6648 VSS.n6301 VSS.n6286 0.0584021
R6649 VSS.n6286 VSS.n6271 0.0231573
R6650 VSS.n6256 VSS.n6271 0.0584021
R6651 VSS.n6241 VSS.n6256 0.0596608
R6652 VSS.n6241 VSS.n6226 0.0244161
R6653 VSS.n6226 VSS.n6211 0.0585594
R6654 VSS.n6211 VSS.n6196 0.0584021
R6655 VSS.n6181 VSS.n6196 0.0596608
R6656 VSS.n6181 VSS.n6166 0.0244161
R6657 VSS.n6166 VSS.n6151 0.0585594
R6658 VSS.n6151 VSS.n6136 0.0584021
R6659 VSS.n6136 VSS 0.16272
R6660 VSS VSS.n6121 0.143052
R6661 VSS.n6106 VSS.n6121 0.0584021
R6662 VSS.n6091 VSS.n6106 0.0584021
R6663 VSS.n6076 VSS.n6091 0.0244161
R6664 VSS.n6076 VSS.n6061 0.0598182
R6665 VSS.n6061 VSS.n6046 0.0584021
R6666 VSS.n6031 VSS.n6046 0.0584021
R6667 VSS.n6016 VSS.n6031 0.0244161
R6668 VSS.n6016 VSS.n6001 0.0598182
R6669 VSS.n6001 VSS.n5986 0.0584021
R6670 VSS.n5986 VSS.n5971 0.0231573
R6671 VSS.n5956 VSS.n5971 0.0584021
R6672 VSS.n5941 VSS.n5956 0.0596608
R6673 VSS.n5941 VSS.n5926 0.0244161
R6674 VSS.n5926 VSS.n5911 0.0585594
R6675 VSS.n5911 VSS.n5896 0.0584021
R6676 VSS.n5881 VSS.n5896 0.0596608
R6677 VSS.n5881 VSS.n5866 0.0244161
R6678 VSS.n5866 VSS.n5851 0.0585594
R6679 VSS.n5851 VSS.n5836 0.0584021
R6680 VSS.n5836 VSS 0.16272
R6681 VSS VSS.n5821 0.143052
R6682 VSS.n5806 VSS.n5821 0.0584021
R6683 VSS.n5791 VSS.n5806 0.0584021
R6684 VSS.n5776 VSS.n5791 0.0244161
R6685 VSS.n5776 VSS.n5761 0.0598182
R6686 VSS.n5761 VSS.n5746 0.0584021
R6687 VSS.n5731 VSS.n5746 0.0584021
R6688 VSS.n5716 VSS.n5731 0.0244161
R6689 VSS.n5716 VSS.n5701 0.0598182
R6690 VSS.n5701 VSS.n5686 0.0584021
R6691 VSS.n5686 VSS.n5671 0.0231573
R6692 VSS.n5656 VSS.n5671 0.0584021
R6693 VSS.n5641 VSS.n5656 0.0596608
R6694 VSS.n5641 VSS.n5626 0.0244161
R6695 VSS.n5626 VSS.n5611 0.0585594
R6696 VSS.n5611 VSS.n5596 0.0584021
R6697 VSS.n5581 VSS.n5596 0.0596608
R6698 VSS.n5581 VSS.n5566 0.0244161
R6699 VSS.n5566 VSS.n5551 0.0585594
R6700 VSS.n5551 VSS.n5536 0.0584021
R6701 VSS.n5536 VSS 0.16272
R6702 VSS VSS.n5521 0.143052
R6703 VSS.n5506 VSS.n5521 0.0584021
R6704 VSS.n5491 VSS.n5506 0.0584021
R6705 VSS.n5476 VSS.n5491 0.0244161
R6706 VSS.n5476 VSS.n5461 0.0598182
R6707 VSS.n5461 VSS.n5446 0.0584021
R6708 VSS.n5431 VSS.n5446 0.0584021
R6709 VSS.n5416 VSS.n5431 0.0244161
R6710 VSS.n5416 VSS.n5401 0.0598182
R6711 VSS.n5401 VSS.n5386 0.0584021
R6712 VSS.n5386 VSS.n5371 0.0231573
R6713 VSS.n5356 VSS.n5371 0.0584021
R6714 VSS.n5341 VSS.n5356 0.0596608
R6715 VSS.n5341 VSS.n5326 0.0244161
R6716 VSS.n5326 VSS.n5311 0.0585594
R6717 VSS.n5311 VSS.n5296 0.0584021
R6718 VSS.n5281 VSS.n5296 0.0596608
R6719 VSS.n5281 VSS.n5266 0.0244161
R6720 VSS.n5266 VSS.n5251 0.0585594
R6721 VSS.n5251 VSS.n5236 0.0584021
R6722 VSS.n5236 VSS 0.16272
R6723 VSS VSS.n5221 0.143052
R6724 VSS.n5206 VSS.n5221 0.0584021
R6725 VSS.n5191 VSS.n5206 0.0584021
R6726 VSS.n5176 VSS.n5191 0.0244161
R6727 VSS.n5176 VSS.n5161 0.0598182
R6728 VSS.n5161 VSS.n5146 0.0584021
R6729 VSS.n5131 VSS.n5146 0.0584021
R6730 VSS.n5116 VSS.n5131 0.0244161
R6731 VSS.n5116 VSS.n5101 0.0598182
R6732 VSS.n5101 VSS.n5086 0.0584021
R6733 VSS.n5086 VSS.n5071 0.0231573
R6734 VSS.n5056 VSS.n5071 0.0584021
R6735 VSS.n5041 VSS.n5056 0.0596608
R6736 VSS.n5041 VSS.n5026 0.0244161
R6737 VSS.n5026 VSS.n5011 0.0585594
R6738 VSS.n5011 VSS.n4996 0.0584021
R6739 VSS.n4981 VSS.n4996 0.0596608
R6740 VSS.n4981 VSS.n4966 0.0244161
R6741 VSS.n4966 VSS.n4951 0.0585594
R6742 VSS.n4951 VSS.n4936 0.0584021
R6743 VSS.n4936 VSS 0.16272
R6744 VSS VSS.n4921 0.143052
R6745 VSS.n4906 VSS.n4921 0.0584021
R6746 VSS.n4891 VSS.n4906 0.0584021
R6747 VSS.n4876 VSS.n4891 0.0244161
R6748 VSS.n4876 VSS.n4861 0.0598182
R6749 VSS.n4861 VSS.n4846 0.0584021
R6750 VSS.n4831 VSS.n4846 0.0584021
R6751 VSS.n4816 VSS.n4831 0.0244161
R6752 VSS.n4816 VSS.n4801 0.0598182
R6753 VSS.n4801 VSS.n4786 0.0584021
R6754 VSS.n7157 VSS.n7162 4.5005
R6755 VSS.n7159 VSS.n7163 4.5005
R6756 VSS.n7160 VSS.n7164 4.5005
R6757 VSS.n7161 VSS.n7165 4.57324
R6758 VSS.n7157 VSS.n7155 0.147342
R6759 VSS.n7158 VSS.n7159 0.0732424
R6760 VSS.n7159 VSS.n7160 0.147342
R6761 VSS.n7162 VSS.n7166 0.0721009
R6762 VSS.n7167 VSS.n7163 4.5005
R6763 VSS.n7168 VSS.n7164 4.5005
R6764 VSS.n7169 VSS.n7165 4.5005
R6765 VSS.n7155 VSS.n7166 4.57442
R6766 VSS.n7162 VSS.n7163 0.147342
R6767 VSS.n7163 VSS.n7164 0.147342
R6768 VSS.n7164 VSS.n7165 0.147342
R6769 VSS.n7166 VSS.n7167 2.39784
R6770 VSS.n7167 VSS.n7168 0.147342
R6771 VSS.n7168 VSS.n7169 0.147342
R6772 VSS.n7169 VSS.t350 3.13212
R6773 VSS.n7142 VSS.n7147 4.5005
R6774 VSS.n7144 VSS.n7148 4.5005
R6775 VSS.n7145 VSS.n7149 4.5005
R6776 VSS.n7146 VSS.n7150 4.57324
R6777 VSS.n7142 VSS.n7140 0.147342
R6778 VSS.n7143 VSS.n7144 0.0732424
R6779 VSS.n7144 VSS.n7145 0.147342
R6780 VSS.n7147 VSS.n7151 0.0721009
R6781 VSS.n7152 VSS.n7148 4.5005
R6782 VSS.n7153 VSS.n7149 4.5005
R6783 VSS.n7154 VSS.n7150 4.5005
R6784 VSS.n7140 VSS.n7151 4.57442
R6785 VSS.n7147 VSS.n7148 0.147342
R6786 VSS.n7148 VSS.n7149 0.147342
R6787 VSS.n7149 VSS.n7150 0.147342
R6788 VSS.n7151 VSS.n7152 2.39784
R6789 VSS.n7152 VSS.n7153 0.147342
R6790 VSS.n7153 VSS.n7154 0.147342
R6791 VSS.n7154 VSS.t297 3.13212
R6792 VSS.n7127 VSS.n7132 4.5005
R6793 VSS.n7129 VSS.n7133 4.5005
R6794 VSS.n7130 VSS.n7134 4.5005
R6795 VSS.n7131 VSS.n7135 4.57324
R6796 VSS.n7127 VSS.n7125 0.147342
R6797 VSS.n7128 VSS.n7129 0.0732424
R6798 VSS.n7129 VSS.n7130 0.147342
R6799 VSS.n7132 VSS.n7136 0.0721009
R6800 VSS.n7137 VSS.n7133 4.5005
R6801 VSS.n7138 VSS.n7134 4.5005
R6802 VSS.n7139 VSS.n7135 4.5005
R6803 VSS.n7125 VSS.n7136 4.57442
R6804 VSS.n7132 VSS.n7133 0.147342
R6805 VSS.n7133 VSS.n7134 0.147342
R6806 VSS.n7134 VSS.n7135 0.147342
R6807 VSS.n7136 VSS.n7137 2.39784
R6808 VSS.n7137 VSS.n7138 0.147342
R6809 VSS.n7138 VSS.n7139 0.147342
R6810 VSS.n7139 VSS.t547 3.13212
R6811 VSS.n7112 VSS.n7117 4.5005
R6812 VSS.n7114 VSS.n7118 4.5005
R6813 VSS.n7115 VSS.n7119 4.5005
R6814 VSS.n7116 VSS.n7120 4.57324
R6815 VSS.n7112 VSS.n7110 0.147342
R6816 VSS.n7113 VSS.n7114 0.0732424
R6817 VSS.n7114 VSS.n7115 0.147342
R6818 VSS.n7117 VSS.n7121 0.0721009
R6819 VSS.n7122 VSS.n7118 4.5005
R6820 VSS.n7123 VSS.n7119 4.5005
R6821 VSS.n7124 VSS.n7120 4.5005
R6822 VSS.n7110 VSS.n7121 4.57442
R6823 VSS.n7117 VSS.n7118 0.147342
R6824 VSS.n7118 VSS.n7119 0.147342
R6825 VSS.n7119 VSS.n7120 0.147342
R6826 VSS.n7121 VSS.n7122 2.39784
R6827 VSS.n7122 VSS.n7123 0.147342
R6828 VSS.n7123 VSS.n7124 0.147342
R6829 VSS.n7124 VSS.t281 3.13212
R6830 VSS.n7097 VSS.n7102 4.5005
R6831 VSS.n7099 VSS.n7103 4.5005
R6832 VSS.n7100 VSS.n7104 4.5005
R6833 VSS.n7101 VSS.n7105 4.57324
R6834 VSS.n7097 VSS.n7095 0.147342
R6835 VSS.n7098 VSS.n7099 0.0732424
R6836 VSS.n7099 VSS.n7100 0.147342
R6837 VSS.n7102 VSS.n7106 0.0721009
R6838 VSS.n7107 VSS.n7103 4.5005
R6839 VSS.n7108 VSS.n7104 4.5005
R6840 VSS.n7109 VSS.n7105 4.5005
R6841 VSS.n7095 VSS.n7106 4.57442
R6842 VSS.n7102 VSS.n7103 0.147342
R6843 VSS.n7103 VSS.n7104 0.147342
R6844 VSS.n7104 VSS.n7105 0.147342
R6845 VSS.n7106 VSS.n7107 2.39784
R6846 VSS.n7107 VSS.n7108 0.147342
R6847 VSS.n7108 VSS.n7109 0.147342
R6848 VSS.n7109 VSS.t163 3.13212
R6849 VSS.n7087 VSS.n7082 4.5005
R6850 VSS.n7088 VSS.n7084 4.5005
R6851 VSS.n7089 VSS.n7085 4.5005
R6852 VSS.n7090 VSS.n7086 4.57324
R6853 VSS.n7080 VSS.n7082 0.147342
R6854 VSS.n7083 VSS.n7084 0.0732424
R6855 VSS.n7084 VSS.n7085 0.147342
R6856 VSS.n7091 VSS.n7087 0.0722544
R6857 VSS.n7092 VSS.n7088 4.5005
R6858 VSS.n7093 VSS.n7089 4.5005
R6859 VSS.n7094 VSS.n7090 4.5005
R6860 VSS.n7091 VSS.n7080 4.57426
R6861 VSS.n7087 VSS.n7088 0.147342
R6862 VSS.n7088 VSS.n7089 0.147342
R6863 VSS.n7089 VSS.n7090 0.147342
R6864 VSS.n7092 VSS.n7091 2.37296
R6865 VSS.n7093 VSS.n7092 0.127318
R6866 VSS.n7094 VSS.n7093 0.127318
R6867 VSS.t0 VSS.n7094 2.73618
R6868 VSS.n7067 VSS.n7072 4.5005
R6869 VSS.n7069 VSS.n7073 4.5005
R6870 VSS.n7070 VSS.n7074 4.5005
R6871 VSS.n7071 VSS.n7075 4.57324
R6872 VSS.n7067 VSS.n7065 0.147342
R6873 VSS.n7068 VSS.n7069 0.0732424
R6874 VSS.n7069 VSS.n7070 0.147342
R6875 VSS.n7072 VSS.n7076 0.0721009
R6876 VSS.n7077 VSS.n7073 4.5005
R6877 VSS.n7078 VSS.n7074 4.5005
R6878 VSS.n7079 VSS.n7075 4.5005
R6879 VSS.n7065 VSS.n7076 4.57442
R6880 VSS.n7072 VSS.n7073 0.147342
R6881 VSS.n7073 VSS.n7074 0.147342
R6882 VSS.n7074 VSS.n7075 0.147342
R6883 VSS.n7076 VSS.n7077 2.39784
R6884 VSS.n7077 VSS.n7078 0.147342
R6885 VSS.n7078 VSS.n7079 0.147342
R6886 VSS.n7079 VSS.t443 3.13212
R6887 VSS.n7052 VSS.n7057 4.5005
R6888 VSS.n7054 VSS.n7058 4.5005
R6889 VSS.n7055 VSS.n7059 4.5005
R6890 VSS.n7056 VSS.n7060 4.57324
R6891 VSS.n7052 VSS.n7050 0.147342
R6892 VSS.n7053 VSS.n7054 0.0732424
R6893 VSS.n7054 VSS.n7055 0.147342
R6894 VSS.n7057 VSS.n7061 0.0721009
R6895 VSS.n7062 VSS.n7058 4.5005
R6896 VSS.n7063 VSS.n7059 4.5005
R6897 VSS.n7064 VSS.n7060 4.5005
R6898 VSS.n7050 VSS.n7061 4.57442
R6899 VSS.n7057 VSS.n7058 0.147342
R6900 VSS.n7058 VSS.n7059 0.147342
R6901 VSS.n7059 VSS.n7060 0.147342
R6902 VSS.n7061 VSS.n7062 2.39784
R6903 VSS.n7062 VSS.n7063 0.147342
R6904 VSS.n7063 VSS.n7064 0.147342
R6905 VSS.n7064 VSS.t157 3.13212
R6906 VSS.n7037 VSS.n7042 4.5005
R6907 VSS.n7039 VSS.n7043 4.5005
R6908 VSS.n7040 VSS.n7044 4.5005
R6909 VSS.n7041 VSS.n7045 4.57324
R6910 VSS.n7037 VSS.n7035 0.147342
R6911 VSS.n7038 VSS.n7039 0.0732424
R6912 VSS.n7039 VSS.n7040 0.147342
R6913 VSS.n7042 VSS.n7046 0.0721009
R6914 VSS.n7047 VSS.n7043 4.5005
R6915 VSS.n7048 VSS.n7044 4.5005
R6916 VSS.n7049 VSS.n7045 4.5005
R6917 VSS.n7035 VSS.n7046 4.57442
R6918 VSS.n7042 VSS.n7043 0.147342
R6919 VSS.n7043 VSS.n7044 0.147342
R6920 VSS.n7044 VSS.n7045 0.147342
R6921 VSS.n7046 VSS.n7047 2.39784
R6922 VSS.n7047 VSS.n7048 0.147342
R6923 VSS.n7048 VSS.n7049 0.147342
R6924 VSS.n7049 VSS.t180 3.13212
R6925 VSS.n7022 VSS.n7027 4.5005
R6926 VSS.n7024 VSS.n7028 4.5005
R6927 VSS.n7025 VSS.n7029 4.5005
R6928 VSS.n7026 VSS.n7030 4.57324
R6929 VSS.n7022 VSS.n7020 0.147342
R6930 VSS.n7023 VSS.n7024 0.0732424
R6931 VSS.n7024 VSS.n7025 0.147342
R6932 VSS.n7027 VSS.n7031 0.0721009
R6933 VSS.n7032 VSS.n7028 4.5005
R6934 VSS.n7033 VSS.n7029 4.5005
R6935 VSS.n7034 VSS.n7030 4.5005
R6936 VSS.n7020 VSS.n7031 4.57442
R6937 VSS.n7027 VSS.n7028 0.147342
R6938 VSS.n7028 VSS.n7029 0.147342
R6939 VSS.n7029 VSS.n7030 0.147342
R6940 VSS.n7031 VSS.n7032 2.39784
R6941 VSS.n7032 VSS.n7033 0.147342
R6942 VSS.n7033 VSS.n7034 0.147342
R6943 VSS.n7034 VSS.t94 3.13212
R6944 VSS.n7007 VSS.n7012 4.5005
R6945 VSS.n7009 VSS.n7013 4.5005
R6946 VSS.n7010 VSS.n7014 4.5005
R6947 VSS.n7011 VSS.n7015 4.57324
R6948 VSS.n7007 VSS.n7005 0.147342
R6949 VSS.n7008 VSS.n7009 0.0732424
R6950 VSS.n7009 VSS.n7010 0.147342
R6951 VSS.n7012 VSS.n7016 0.0721009
R6952 VSS.n7017 VSS.n7013 4.5005
R6953 VSS.n7018 VSS.n7014 4.5005
R6954 VSS.n7019 VSS.n7015 4.5005
R6955 VSS.n7005 VSS.n7016 4.57442
R6956 VSS.n7012 VSS.n7013 0.147342
R6957 VSS.n7013 VSS.n7014 0.147342
R6958 VSS.n7014 VSS.n7015 0.147342
R6959 VSS.n7016 VSS.n7017 2.39784
R6960 VSS.n7017 VSS.n7018 0.147342
R6961 VSS.n7018 VSS.n7019 0.147342
R6962 VSS.n7019 VSS.t484 3.13212
R6963 VSS.n6992 VSS.n6997 4.5005
R6964 VSS.n6994 VSS.n6998 4.5005
R6965 VSS.n6995 VSS.n6999 4.5005
R6966 VSS.n6996 VSS.n7000 4.57324
R6967 VSS.n6992 VSS.n6990 0.147342
R6968 VSS.n6993 VSS.n6994 0.0732424
R6969 VSS.n6994 VSS.n6995 0.147342
R6970 VSS.n6997 VSS.n7001 0.0721009
R6971 VSS.n7002 VSS.n6998 4.5005
R6972 VSS.n7003 VSS.n6999 4.5005
R6973 VSS.n7004 VSS.n7000 4.5005
R6974 VSS.n6990 VSS.n7001 4.57442
R6975 VSS.n6997 VSS.n6998 0.147342
R6976 VSS.n6998 VSS.n6999 0.147342
R6977 VSS.n6999 VSS.n7000 0.147342
R6978 VSS.n7001 VSS.n7002 2.39784
R6979 VSS.n7002 VSS.n7003 0.147342
R6980 VSS.n7003 VSS.n7004 0.147342
R6981 VSS.n7004 VSS.t511 3.13212
R6982 VSS.n6982 VSS.n6977 4.5005
R6983 VSS.n6983 VSS.n6979 4.5005
R6984 VSS.n6984 VSS.n6980 4.5005
R6985 VSS.n6985 VSS.n6981 4.57324
R6986 VSS.n6975 VSS.n6977 0.147342
R6987 VSS.n6978 VSS.n6979 0.0732424
R6988 VSS.n6979 VSS.n6980 0.147342
R6989 VSS.n6986 VSS.n6982 0.0722544
R6990 VSS.n6987 VSS.n6983 4.5005
R6991 VSS.n6988 VSS.n6984 4.5005
R6992 VSS.n6989 VSS.n6985 4.5005
R6993 VSS.n6986 VSS.n6975 4.57426
R6994 VSS.n6982 VSS.n6983 0.147342
R6995 VSS.n6983 VSS.n6984 0.147342
R6996 VSS.n6984 VSS.n6985 0.147342
R6997 VSS.n6987 VSS.n6986 2.37296
R6998 VSS.n6988 VSS.n6987 0.127318
R6999 VSS.n6989 VSS.n6988 0.127318
R7000 VSS.t0 VSS.n6989 2.73618
R7001 VSS.n6962 VSS.n6967 4.5005
R7002 VSS.n6964 VSS.n6968 4.5005
R7003 VSS.n6965 VSS.n6969 4.5005
R7004 VSS.n6966 VSS.n6970 4.57324
R7005 VSS.n6962 VSS.n6960 0.147342
R7006 VSS.n6963 VSS.n6964 0.0732424
R7007 VSS.n6964 VSS.n6965 0.147342
R7008 VSS.n6967 VSS.n6971 0.0721009
R7009 VSS.n6972 VSS.n6968 4.5005
R7010 VSS.n6973 VSS.n6969 4.5005
R7011 VSS.n6974 VSS.n6970 4.5005
R7012 VSS.n6960 VSS.n6971 4.57442
R7013 VSS.n6967 VSS.n6968 0.147342
R7014 VSS.n6968 VSS.n6969 0.147342
R7015 VSS.n6969 VSS.n6970 0.147342
R7016 VSS.n6971 VSS.n6972 2.39784
R7017 VSS.n6972 VSS.n6973 0.147342
R7018 VSS.n6973 VSS.n6974 0.147342
R7019 VSS.n6974 VSS.t35 3.13212
R7020 VSS.n6947 VSS.n6952 4.5005
R7021 VSS.n6949 VSS.n6953 4.5005
R7022 VSS.n6950 VSS.n6954 4.5005
R7023 VSS.n6951 VSS.n6955 4.57324
R7024 VSS.n6947 VSS.n6945 0.147342
R7025 VSS.n6948 VSS.n6949 0.0732424
R7026 VSS.n6949 VSS.n6950 0.147342
R7027 VSS.n6952 VSS.n6956 0.0721009
R7028 VSS.n6957 VSS.n6953 4.5005
R7029 VSS.n6958 VSS.n6954 4.5005
R7030 VSS.n6959 VSS.n6955 4.5005
R7031 VSS.n6945 VSS.n6956 4.57442
R7032 VSS.n6952 VSS.n6953 0.147342
R7033 VSS.n6953 VSS.n6954 0.147342
R7034 VSS.n6954 VSS.n6955 0.147342
R7035 VSS.n6956 VSS.n6957 2.39784
R7036 VSS.n6957 VSS.n6958 0.147342
R7037 VSS.n6958 VSS.n6959 0.147342
R7038 VSS.n6959 VSS.t105 3.13212
R7039 VSS.n6932 VSS.n6937 4.5005
R7040 VSS.n6934 VSS.n6938 4.5005
R7041 VSS.n6935 VSS.n6939 4.5005
R7042 VSS.n6936 VSS.n6940 4.57324
R7043 VSS.n6932 VSS.n6930 0.147342
R7044 VSS.n6933 VSS.n6934 0.0732424
R7045 VSS.n6934 VSS.n6935 0.147342
R7046 VSS.n6937 VSS.n6941 0.0721009
R7047 VSS.n6942 VSS.n6938 4.5005
R7048 VSS.n6943 VSS.n6939 4.5005
R7049 VSS.n6944 VSS.n6940 4.5005
R7050 VSS.n6930 VSS.n6941 4.57442
R7051 VSS.n6937 VSS.n6938 0.147342
R7052 VSS.n6938 VSS.n6939 0.147342
R7053 VSS.n6939 VSS.n6940 0.147342
R7054 VSS.n6941 VSS.n6942 2.39784
R7055 VSS.n6942 VSS.n6943 0.147342
R7056 VSS.n6943 VSS.n6944 0.147342
R7057 VSS.n6944 VSS.t238 3.13212
R7058 VSS.n6922 VSS.n6917 4.5005
R7059 VSS.n6923 VSS.n6919 4.5005
R7060 VSS.n6924 VSS.n6920 4.5005
R7061 VSS.n6925 VSS.n6921 4.57324
R7062 VSS.n6915 VSS.n6917 0.147342
R7063 VSS.n6918 VSS.n6919 0.0732424
R7064 VSS.n6919 VSS.n6920 0.147342
R7065 VSS.n6926 VSS.n6922 0.0722544
R7066 VSS.n6927 VSS.n6923 4.5005
R7067 VSS.n6928 VSS.n6924 4.5005
R7068 VSS.n6929 VSS.n6925 4.5005
R7069 VSS.n6926 VSS.n6915 4.57426
R7070 VSS.n6922 VSS.n6923 0.147342
R7071 VSS.n6923 VSS.n6924 0.147342
R7072 VSS.n6924 VSS.n6925 0.147342
R7073 VSS.n6927 VSS.n6926 2.37296
R7074 VSS.n6928 VSS.n6927 0.127318
R7075 VSS.n6929 VSS.n6928 0.127318
R7076 VSS.t0 VSS.n6929 2.73618
R7077 VSS.n6902 VSS.n6907 4.5005
R7078 VSS.n6904 VSS.n6908 4.5005
R7079 VSS.n6905 VSS.n6909 4.5005
R7080 VSS.n6906 VSS.n6910 4.57324
R7081 VSS.n6902 VSS.n6900 0.147342
R7082 VSS.n6903 VSS.n6904 0.0732424
R7083 VSS.n6904 VSS.n6905 0.147342
R7084 VSS.n6907 VSS.n6911 0.0721009
R7085 VSS.n6912 VSS.n6908 4.5005
R7086 VSS.n6913 VSS.n6909 4.5005
R7087 VSS.n6914 VSS.n6910 4.5005
R7088 VSS.n6900 VSS.n6911 4.57442
R7089 VSS.n6907 VSS.n6908 0.147342
R7090 VSS.n6908 VSS.n6909 0.147342
R7091 VSS.n6909 VSS.n6910 0.147342
R7092 VSS.n6911 VSS.n6912 2.39784
R7093 VSS.n6912 VSS.n6913 0.147342
R7094 VSS.n6913 VSS.n6914 0.147342
R7095 VSS.n6914 VSS.t134 3.13212
R7096 VSS.n6887 VSS.n6892 4.5005
R7097 VSS.n6889 VSS.n6893 4.5005
R7098 VSS.n6890 VSS.n6894 4.5005
R7099 VSS.n6891 VSS.n6895 4.57324
R7100 VSS.n6887 VSS.n6885 0.147342
R7101 VSS.n6888 VSS.n6889 0.0732424
R7102 VSS.n6889 VSS.n6890 0.147342
R7103 VSS.n6892 VSS.n6896 0.0721009
R7104 VSS.n6897 VSS.n6893 4.5005
R7105 VSS.n6898 VSS.n6894 4.5005
R7106 VSS.n6899 VSS.n6895 4.5005
R7107 VSS.n6885 VSS.n6896 4.57442
R7108 VSS.n6892 VSS.n6893 0.147342
R7109 VSS.n6893 VSS.n6894 0.147342
R7110 VSS.n6894 VSS.n6895 0.147342
R7111 VSS.n6896 VSS.n6897 2.39784
R7112 VSS.n6897 VSS.n6898 0.147342
R7113 VSS.n6898 VSS.n6899 0.147342
R7114 VSS.n6899 VSS.t137 3.13212
R7115 VSS.n6872 VSS.n6877 4.5005
R7116 VSS.n6874 VSS.n6878 4.5005
R7117 VSS.n6875 VSS.n6879 4.5005
R7118 VSS.n6876 VSS.n6880 4.57324
R7119 VSS.n6872 VSS.n6870 0.147342
R7120 VSS.n6873 VSS.n6874 0.0732424
R7121 VSS.n6874 VSS.n6875 0.147342
R7122 VSS.n6877 VSS.n6881 0.0721009
R7123 VSS.n6882 VSS.n6878 4.5005
R7124 VSS.n6883 VSS.n6879 4.5005
R7125 VSS.n6884 VSS.n6880 4.5005
R7126 VSS.n6870 VSS.n6881 4.57442
R7127 VSS.n6877 VSS.n6878 0.147342
R7128 VSS.n6878 VSS.n6879 0.147342
R7129 VSS.n6879 VSS.n6880 0.147342
R7130 VSS.n6881 VSS.n6882 2.39784
R7131 VSS.n6882 VSS.n6883 0.147342
R7132 VSS.n6883 VSS.n6884 0.147342
R7133 VSS.n6884 VSS.t351 3.13212
R7134 VSS.n6857 VSS.n6862 4.5005
R7135 VSS.n6859 VSS.n6863 4.5005
R7136 VSS.n6860 VSS.n6864 4.5005
R7137 VSS.n6861 VSS.n6865 4.57324
R7138 VSS.n6857 VSS.n6855 0.147342
R7139 VSS.n6858 VSS.n6859 0.0732424
R7140 VSS.n6859 VSS.n6860 0.147342
R7141 VSS.n6862 VSS.n6866 0.0721009
R7142 VSS.n6867 VSS.n6863 4.5005
R7143 VSS.n6868 VSS.n6864 4.5005
R7144 VSS.n6869 VSS.n6865 4.5005
R7145 VSS.n6855 VSS.n6866 4.57442
R7146 VSS.n6862 VSS.n6863 0.147342
R7147 VSS.n6863 VSS.n6864 0.147342
R7148 VSS.n6864 VSS.n6865 0.147342
R7149 VSS.n6866 VSS.n6867 2.39784
R7150 VSS.n6867 VSS.n6868 0.147342
R7151 VSS.n6868 VSS.n6869 0.147342
R7152 VSS.n6869 VSS.t307 3.13212
R7153 VSS.n6847 VSS.n6842 4.5005
R7154 VSS.n6848 VSS.n6844 4.5005
R7155 VSS.n6849 VSS.n6845 4.5005
R7156 VSS.n6850 VSS.n6846 4.57324
R7157 VSS.n6840 VSS.n6842 0.147342
R7158 VSS.n6843 VSS.n6844 0.0732424
R7159 VSS.n6844 VSS.n6845 0.147342
R7160 VSS.n6851 VSS.n6847 0.0722544
R7161 VSS.n6852 VSS.n6848 4.5005
R7162 VSS.n6853 VSS.n6849 4.5005
R7163 VSS.n6854 VSS.n6850 4.5005
R7164 VSS.n6851 VSS.n6840 4.57426
R7165 VSS.n6847 VSS.n6848 0.147342
R7166 VSS.n6848 VSS.n6849 0.147342
R7167 VSS.n6849 VSS.n6850 0.147342
R7168 VSS.n6852 VSS.n6851 2.37296
R7169 VSS.n6853 VSS.n6852 0.127318
R7170 VSS.n6854 VSS.n6853 0.127318
R7171 VSS.t0 VSS.n6854 2.73618
R7172 VSS.n6827 VSS.n6832 4.5005
R7173 VSS.n6829 VSS.n6833 4.5005
R7174 VSS.n6830 VSS.n6834 4.5005
R7175 VSS.n6831 VSS.n6835 4.57324
R7176 VSS.n6827 VSS.n6825 0.147342
R7177 VSS.n6828 VSS.n6829 0.0732424
R7178 VSS.n6829 VSS.n6830 0.147342
R7179 VSS.n6832 VSS.n6836 0.0721009
R7180 VSS.n6837 VSS.n6833 4.5005
R7181 VSS.n6838 VSS.n6834 4.5005
R7182 VSS.n6839 VSS.n6835 4.5005
R7183 VSS.n6825 VSS.n6836 4.57442
R7184 VSS.n6832 VSS.n6833 0.147342
R7185 VSS.n6833 VSS.n6834 0.147342
R7186 VSS.n6834 VSS.n6835 0.147342
R7187 VSS.n6836 VSS.n6837 2.39784
R7188 VSS.n6837 VSS.n6838 0.147342
R7189 VSS.n6838 VSS.n6839 0.147342
R7190 VSS.n6839 VSS.t550 3.13212
R7191 VSS.n6812 VSS.n6817 4.5005
R7192 VSS.n6814 VSS.n6818 4.5005
R7193 VSS.n6815 VSS.n6819 4.5005
R7194 VSS.n6816 VSS.n6820 4.57324
R7195 VSS.n6812 VSS.n6810 0.147342
R7196 VSS.n6813 VSS.n6814 0.0732424
R7197 VSS.n6814 VSS.n6815 0.147342
R7198 VSS.n6817 VSS.n6821 0.0721009
R7199 VSS.n6822 VSS.n6818 4.5005
R7200 VSS.n6823 VSS.n6819 4.5005
R7201 VSS.n6824 VSS.n6820 4.5005
R7202 VSS.n6810 VSS.n6821 4.57442
R7203 VSS.n6817 VSS.n6818 0.147342
R7204 VSS.n6818 VSS.n6819 0.147342
R7205 VSS.n6819 VSS.n6820 0.147342
R7206 VSS.n6821 VSS.n6822 2.39784
R7207 VSS.n6822 VSS.n6823 0.147342
R7208 VSS.n6823 VSS.n6824 0.147342
R7209 VSS.n6824 VSS.t279 3.13212
R7210 VSS.n6797 VSS.n6802 4.5005
R7211 VSS.n6799 VSS.n6803 4.5005
R7212 VSS.n6800 VSS.n6804 4.5005
R7213 VSS.n6801 VSS.n6805 4.57324
R7214 VSS.n6797 VSS.n6795 0.147342
R7215 VSS.n6798 VSS.n6799 0.0732424
R7216 VSS.n6799 VSS.n6800 0.147342
R7217 VSS.n6802 VSS.n6806 0.0721009
R7218 VSS.n6807 VSS.n6803 4.5005
R7219 VSS.n6808 VSS.n6804 4.5005
R7220 VSS.n6809 VSS.n6805 4.5005
R7221 VSS.n6795 VSS.n6806 4.57442
R7222 VSS.n6802 VSS.n6803 0.147342
R7223 VSS.n6803 VSS.n6804 0.147342
R7224 VSS.n6804 VSS.n6805 0.147342
R7225 VSS.n6806 VSS.n6807 2.39784
R7226 VSS.n6807 VSS.n6808 0.147342
R7227 VSS.n6808 VSS.n6809 0.147342
R7228 VSS.n6809 VSS.t599 3.13212
R7229 VSS.n6787 VSS.n6782 4.5005
R7230 VSS.n6788 VSS.n6784 4.5005
R7231 VSS.n6789 VSS.n6785 4.5005
R7232 VSS.n6790 VSS.n6786 4.57324
R7233 VSS.n6780 VSS.n6782 0.147342
R7234 VSS.n6783 VSS.n6784 0.0732424
R7235 VSS.n6784 VSS.n6785 0.147342
R7236 VSS.n6791 VSS.n6787 0.0722544
R7237 VSS.n6792 VSS.n6788 4.5005
R7238 VSS.n6793 VSS.n6789 4.5005
R7239 VSS.n6794 VSS.n6790 4.5005
R7240 VSS.n6791 VSS.n6780 4.57426
R7241 VSS.n6787 VSS.n6788 0.147342
R7242 VSS.n6788 VSS.n6789 0.147342
R7243 VSS.n6789 VSS.n6790 0.147342
R7244 VSS.n6792 VSS.n6791 2.37296
R7245 VSS.n6793 VSS.n6792 0.127318
R7246 VSS.n6794 VSS.n6793 0.127318
R7247 VSS.t0 VSS.n6794 2.73618
R7248 VSS.n6767 VSS.n6772 4.5005
R7249 VSS.n6769 VSS.n6773 4.5005
R7250 VSS.n6770 VSS.n6774 4.5005
R7251 VSS.n6771 VSS.n6775 4.57324
R7252 VSS.n6767 VSS.n6765 0.147342
R7253 VSS.n6768 VSS.n6769 0.0732424
R7254 VSS.n6769 VSS.n6770 0.147342
R7255 VSS.n6772 VSS.n6776 0.0721009
R7256 VSS.n6777 VSS.n6773 4.5005
R7257 VSS.n6778 VSS.n6774 4.5005
R7258 VSS.n6779 VSS.n6775 4.5005
R7259 VSS.n6765 VSS.n6776 4.57442
R7260 VSS.n6772 VSS.n6773 0.147342
R7261 VSS.n6773 VSS.n6774 0.147342
R7262 VSS.n6774 VSS.n6775 0.147342
R7263 VSS.n6776 VSS.n6777 2.39784
R7264 VSS.n6777 VSS.n6778 0.147342
R7265 VSS.n6778 VSS.n6779 0.147342
R7266 VSS.n6779 VSS.t441 3.13212
R7267 VSS.n6752 VSS.n6757 4.5005
R7268 VSS.n6754 VSS.n6758 4.5005
R7269 VSS.n6755 VSS.n6759 4.5005
R7270 VSS.n6756 VSS.n6760 4.57324
R7271 VSS.n6752 VSS.n6750 0.147342
R7272 VSS.n6753 VSS.n6754 0.0732424
R7273 VSS.n6754 VSS.n6755 0.147342
R7274 VSS.n6757 VSS.n6761 0.0721009
R7275 VSS.n6762 VSS.n6758 4.5005
R7276 VSS.n6763 VSS.n6759 4.5005
R7277 VSS.n6764 VSS.n6760 4.5005
R7278 VSS.n6750 VSS.n6761 4.57442
R7279 VSS.n6757 VSS.n6758 0.147342
R7280 VSS.n6758 VSS.n6759 0.147342
R7281 VSS.n6759 VSS.n6760 0.147342
R7282 VSS.n6761 VSS.n6762 2.39784
R7283 VSS.n6762 VSS.n6763 0.147342
R7284 VSS.n6763 VSS.n6764 0.147342
R7285 VSS.n6764 VSS.t154 3.13212
R7286 VSS.n6737 VSS.n6742 4.5005
R7287 VSS.n6739 VSS.n6743 4.5005
R7288 VSS.n6740 VSS.n6744 4.5005
R7289 VSS.n6741 VSS.n6745 4.57324
R7290 VSS.n6737 VSS.n6735 0.147342
R7291 VSS.n6738 VSS.n6739 0.0732424
R7292 VSS.n6739 VSS.n6740 0.147342
R7293 VSS.n6742 VSS.n6746 0.0721009
R7294 VSS.n6747 VSS.n6743 4.5005
R7295 VSS.n6748 VSS.n6744 4.5005
R7296 VSS.n6749 VSS.n6745 4.5005
R7297 VSS.n6735 VSS.n6746 4.57442
R7298 VSS.n6742 VSS.n6743 0.147342
R7299 VSS.n6743 VSS.n6744 0.147342
R7300 VSS.n6744 VSS.n6745 0.147342
R7301 VSS.n6746 VSS.n6747 2.39784
R7302 VSS.n6747 VSS.n6748 0.147342
R7303 VSS.n6748 VSS.n6749 0.147342
R7304 VSS.n6749 VSS.t178 3.13212
R7305 VSS.n6722 VSS.n6727 4.5005
R7306 VSS.n6724 VSS.n6728 4.5005
R7307 VSS.n6725 VSS.n6729 4.5005
R7308 VSS.n6726 VSS.n6730 4.57324
R7309 VSS.n6722 VSS.n6720 0.147342
R7310 VSS.n6723 VSS.n6724 0.0732424
R7311 VSS.n6724 VSS.n6725 0.147342
R7312 VSS.n6727 VSS.n6731 0.0721009
R7313 VSS.n6732 VSS.n6728 4.5005
R7314 VSS.n6733 VSS.n6729 4.5005
R7315 VSS.n6734 VSS.n6730 4.5005
R7316 VSS.n6720 VSS.n6731 4.57442
R7317 VSS.n6727 VSS.n6728 0.147342
R7318 VSS.n6728 VSS.n6729 0.147342
R7319 VSS.n6729 VSS.n6730 0.147342
R7320 VSS.n6731 VSS.n6732 2.39784
R7321 VSS.n6732 VSS.n6733 0.147342
R7322 VSS.n6733 VSS.n6734 0.147342
R7323 VSS.n6734 VSS.t266 3.13212
R7324 VSS.n6707 VSS.n6712 4.5005
R7325 VSS.n6709 VSS.n6713 4.5005
R7326 VSS.n6710 VSS.n6714 4.5005
R7327 VSS.n6711 VSS.n6715 4.57324
R7328 VSS.n6707 VSS.n6705 0.147342
R7329 VSS.n6708 VSS.n6709 0.0732424
R7330 VSS.n6709 VSS.n6710 0.147342
R7331 VSS.n6712 VSS.n6716 0.0721009
R7332 VSS.n6717 VSS.n6713 4.5005
R7333 VSS.n6718 VSS.n6714 4.5005
R7334 VSS.n6719 VSS.n6715 4.5005
R7335 VSS.n6705 VSS.n6716 4.57442
R7336 VSS.n6712 VSS.n6713 0.147342
R7337 VSS.n6713 VSS.n6714 0.147342
R7338 VSS.n6714 VSS.n6715 0.147342
R7339 VSS.n6716 VSS.n6717 2.39784
R7340 VSS.n6717 VSS.n6718 0.147342
R7341 VSS.n6718 VSS.n6719 0.147342
R7342 VSS.n6719 VSS.t482 3.13212
R7343 VSS.n6692 VSS.n6697 4.5005
R7344 VSS.n6694 VSS.n6698 4.5005
R7345 VSS.n6695 VSS.n6699 4.5005
R7346 VSS.n6696 VSS.n6700 4.57324
R7347 VSS.n6692 VSS.n6690 0.147342
R7348 VSS.n6693 VSS.n6694 0.0732424
R7349 VSS.n6694 VSS.n6695 0.147342
R7350 VSS.n6697 VSS.n6701 0.0721009
R7351 VSS.n6702 VSS.n6698 4.5005
R7352 VSS.n6703 VSS.n6699 4.5005
R7353 VSS.n6704 VSS.n6700 4.5005
R7354 VSS.n6690 VSS.n6701 4.57442
R7355 VSS.n6697 VSS.n6698 0.147342
R7356 VSS.n6698 VSS.n6699 0.147342
R7357 VSS.n6699 VSS.n6700 0.147342
R7358 VSS.n6701 VSS.n6702 2.39784
R7359 VSS.n6702 VSS.n6703 0.147342
R7360 VSS.n6703 VSS.n6704 0.147342
R7361 VSS.n6704 VSS.t64 3.13212
R7362 VSS.n6682 VSS.n6677 4.5005
R7363 VSS.n6683 VSS.n6679 4.5005
R7364 VSS.n6684 VSS.n6680 4.5005
R7365 VSS.n6685 VSS.n6681 4.57324
R7366 VSS.n6675 VSS.n6677 0.147342
R7367 VSS.n6678 VSS.n6679 0.0732424
R7368 VSS.n6679 VSS.n6680 0.147342
R7369 VSS.n6686 VSS.n6682 0.0722544
R7370 VSS.n6687 VSS.n6683 4.5005
R7371 VSS.n6688 VSS.n6684 4.5005
R7372 VSS.n6689 VSS.n6685 4.5005
R7373 VSS.n6686 VSS.n6675 4.57426
R7374 VSS.n6682 VSS.n6683 0.147342
R7375 VSS.n6683 VSS.n6684 0.147342
R7376 VSS.n6684 VSS.n6685 0.147342
R7377 VSS.n6687 VSS.n6686 2.37296
R7378 VSS.n6688 VSS.n6687 0.127318
R7379 VSS.n6689 VSS.n6688 0.127318
R7380 VSS.t0 VSS.n6689 2.73618
R7381 VSS.n6662 VSS.n6667 4.5005
R7382 VSS.n6664 VSS.n6668 4.5005
R7383 VSS.n6665 VSS.n6669 4.5005
R7384 VSS.n6666 VSS.n6670 4.57324
R7385 VSS.n6662 VSS.n6660 0.147342
R7386 VSS.n6663 VSS.n6664 0.0732424
R7387 VSS.n6664 VSS.n6665 0.147342
R7388 VSS.n6667 VSS.n6671 0.0721009
R7389 VSS.n6672 VSS.n6668 4.5005
R7390 VSS.n6673 VSS.n6669 4.5005
R7391 VSS.n6674 VSS.n6670 4.5005
R7392 VSS.n6660 VSS.n6671 4.57442
R7393 VSS.n6667 VSS.n6668 0.147342
R7394 VSS.n6668 VSS.n6669 0.147342
R7395 VSS.n6669 VSS.n6670 0.147342
R7396 VSS.n6671 VSS.n6672 2.39784
R7397 VSS.n6672 VSS.n6673 0.147342
R7398 VSS.n6673 VSS.n6674 0.147342
R7399 VSS.n6674 VSS.t215 3.13212
R7400 VSS.n6647 VSS.n6652 4.5005
R7401 VSS.n6649 VSS.n6653 4.5005
R7402 VSS.n6650 VSS.n6654 4.5005
R7403 VSS.n6651 VSS.n6655 4.57324
R7404 VSS.n6647 VSS.n6645 0.147342
R7405 VSS.n6648 VSS.n6649 0.0732424
R7406 VSS.n6649 VSS.n6650 0.147342
R7407 VSS.n6652 VSS.n6656 0.0721009
R7408 VSS.n6657 VSS.n6653 4.5005
R7409 VSS.n6658 VSS.n6654 4.5005
R7410 VSS.n6659 VSS.n6655 4.5005
R7411 VSS.n6645 VSS.n6656 4.57442
R7412 VSS.n6652 VSS.n6653 0.147342
R7413 VSS.n6653 VSS.n6654 0.147342
R7414 VSS.n6654 VSS.n6655 0.147342
R7415 VSS.n6656 VSS.n6657 2.39784
R7416 VSS.n6657 VSS.n6658 0.147342
R7417 VSS.n6658 VSS.n6659 0.147342
R7418 VSS.n6659 VSS.t211 3.13212
R7419 VSS.n6632 VSS.n6637 4.5005
R7420 VSS.n6634 VSS.n6638 4.5005
R7421 VSS.n6635 VSS.n6639 4.5005
R7422 VSS.n6636 VSS.n6640 4.57324
R7423 VSS.n6632 VSS.n6630 0.147342
R7424 VSS.n6633 VSS.n6634 0.0732424
R7425 VSS.n6634 VSS.n6635 0.147342
R7426 VSS.n6637 VSS.n6641 0.0721009
R7427 VSS.n6642 VSS.n6638 4.5005
R7428 VSS.n6643 VSS.n6639 4.5005
R7429 VSS.n6644 VSS.n6640 4.5005
R7430 VSS.n6630 VSS.n6641 4.57442
R7431 VSS.n6637 VSS.n6638 0.147342
R7432 VSS.n6638 VSS.n6639 0.147342
R7433 VSS.n6639 VSS.n6640 0.147342
R7434 VSS.n6641 VSS.n6642 2.39784
R7435 VSS.n6642 VSS.n6643 0.147342
R7436 VSS.n6643 VSS.n6644 0.147342
R7437 VSS.n6644 VSS.t130 3.13212
R7438 VSS.n6622 VSS.n6617 4.5005
R7439 VSS.n6623 VSS.n6619 4.5005
R7440 VSS.n6624 VSS.n6620 4.5005
R7441 VSS.n6625 VSS.n6621 4.57324
R7442 VSS.n6615 VSS.n6617 0.147342
R7443 VSS.n6618 VSS.n6619 0.0732424
R7444 VSS.n6619 VSS.n6620 0.147342
R7445 VSS.n6626 VSS.n6622 0.0722544
R7446 VSS.n6627 VSS.n6623 4.5005
R7447 VSS.n6628 VSS.n6624 4.5005
R7448 VSS.n6629 VSS.n6625 4.5005
R7449 VSS.n6626 VSS.n6615 4.57426
R7450 VSS.n6622 VSS.n6623 0.147342
R7451 VSS.n6623 VSS.n6624 0.147342
R7452 VSS.n6624 VSS.n6625 0.147342
R7453 VSS.n6627 VSS.n6626 2.37296
R7454 VSS.n6628 VSS.n6627 0.127318
R7455 VSS.n6629 VSS.n6628 0.127318
R7456 VSS.t0 VSS.n6629 2.73618
R7457 VSS.n6602 VSS.n6607 4.5005
R7458 VSS.n6604 VSS.n6608 4.5005
R7459 VSS.n6605 VSS.n6609 4.5005
R7460 VSS.n6606 VSS.n6610 4.57324
R7461 VSS.n6602 VSS.n6600 0.147342
R7462 VSS.n6603 VSS.n6604 0.0732424
R7463 VSS.n6604 VSS.n6605 0.147342
R7464 VSS.n6607 VSS.n6611 0.0721009
R7465 VSS.n6612 VSS.n6608 4.5005
R7466 VSS.n6613 VSS.n6609 4.5005
R7467 VSS.n6614 VSS.n6610 4.5005
R7468 VSS.n6600 VSS.n6611 4.57442
R7469 VSS.n6607 VSS.n6608 0.147342
R7470 VSS.n6608 VSS.n6609 0.147342
R7471 VSS.n6609 VSS.n6610 0.147342
R7472 VSS.n6611 VSS.n6612 2.39784
R7473 VSS.n6612 VSS.n6613 0.147342
R7474 VSS.n6613 VSS.n6614 0.147342
R7475 VSS.n6614 VSS.t141 3.13212
R7476 VSS.n6587 VSS.n6592 4.5005
R7477 VSS.n6589 VSS.n6593 4.5005
R7478 VSS.n6590 VSS.n6594 4.5005
R7479 VSS.n6591 VSS.n6595 4.57324
R7480 VSS.n6587 VSS.n6585 0.147342
R7481 VSS.n6588 VSS.n6589 0.0732424
R7482 VSS.n6589 VSS.n6590 0.147342
R7483 VSS.n6592 VSS.n6596 0.0721009
R7484 VSS.n6597 VSS.n6593 4.5005
R7485 VSS.n6598 VSS.n6594 4.5005
R7486 VSS.n6599 VSS.n6595 4.5005
R7487 VSS.n6585 VSS.n6596 4.57442
R7488 VSS.n6592 VSS.n6593 0.147342
R7489 VSS.n6593 VSS.n6594 0.147342
R7490 VSS.n6594 VSS.n6595 0.147342
R7491 VSS.n6596 VSS.n6597 2.39784
R7492 VSS.n6597 VSS.n6598 0.147342
R7493 VSS.n6598 VSS.n6599 0.147342
R7494 VSS.n6599 VSS.t100 3.13212
R7495 VSS.n6572 VSS.n6577 4.5005
R7496 VSS.n6574 VSS.n6578 4.5005
R7497 VSS.n6575 VSS.n6579 4.5005
R7498 VSS.n6576 VSS.n6580 4.57324
R7499 VSS.n6572 VSS.n6570 0.147342
R7500 VSS.n6573 VSS.n6574 0.0732424
R7501 VSS.n6574 VSS.n6575 0.147342
R7502 VSS.n6577 VSS.n6581 0.0721009
R7503 VSS.n6582 VSS.n6578 4.5005
R7504 VSS.n6583 VSS.n6579 4.5005
R7505 VSS.n6584 VSS.n6580 4.5005
R7506 VSS.n6570 VSS.n6581 4.57442
R7507 VSS.n6577 VSS.n6578 0.147342
R7508 VSS.n6578 VSS.n6579 0.147342
R7509 VSS.n6579 VSS.n6580 0.147342
R7510 VSS.n6581 VSS.n6582 2.39784
R7511 VSS.n6582 VSS.n6583 0.147342
R7512 VSS.n6583 VSS.n6584 0.147342
R7513 VSS.n6584 VSS.t287 3.13212
R7514 VSS.n6557 VSS.n6562 4.5005
R7515 VSS.n6559 VSS.n6563 4.5005
R7516 VSS.n6560 VSS.n6564 4.5005
R7517 VSS.n6561 VSS.n6565 4.57324
R7518 VSS.n6557 VSS.n6555 0.147342
R7519 VSS.n6558 VSS.n6559 0.0732424
R7520 VSS.n6559 VSS.n6560 0.147342
R7521 VSS.n6562 VSS.n6566 0.0721009
R7522 VSS.n6567 VSS.n6563 4.5005
R7523 VSS.n6568 VSS.n6564 4.5005
R7524 VSS.n6569 VSS.n6565 4.5005
R7525 VSS.n6555 VSS.n6566 4.57442
R7526 VSS.n6562 VSS.n6563 0.147342
R7527 VSS.n6563 VSS.n6564 0.147342
R7528 VSS.n6564 VSS.n6565 0.147342
R7529 VSS.n6566 VSS.n6567 2.39784
R7530 VSS.n6567 VSS.n6568 0.147342
R7531 VSS.n6568 VSS.n6569 0.147342
R7532 VSS.n6569 VSS.t310 3.13212
R7533 VSS.n6547 VSS.n6542 4.5005
R7534 VSS.n6548 VSS.n6544 4.5005
R7535 VSS.n6549 VSS.n6545 4.5005
R7536 VSS.n6550 VSS.n6546 4.57324
R7537 VSS.n6540 VSS.n6542 0.147342
R7538 VSS.n6543 VSS.n6544 0.0732424
R7539 VSS.n6544 VSS.n6545 0.147342
R7540 VSS.n6551 VSS.n6547 0.0722544
R7541 VSS.n6552 VSS.n6548 4.5005
R7542 VSS.n6553 VSS.n6549 4.5005
R7543 VSS.n6554 VSS.n6550 4.5005
R7544 VSS.n6551 VSS.n6540 4.57426
R7545 VSS.n6547 VSS.n6548 0.147342
R7546 VSS.n6548 VSS.n6549 0.147342
R7547 VSS.n6549 VSS.n6550 0.147342
R7548 VSS.n6552 VSS.n6551 2.37296
R7549 VSS.n6553 VSS.n6552 0.127318
R7550 VSS.n6554 VSS.n6553 0.127318
R7551 VSS.t0 VSS.n6554 2.73618
R7552 VSS.n6527 VSS.n6532 4.5005
R7553 VSS.n6529 VSS.n6533 4.5005
R7554 VSS.n6530 VSS.n6534 4.5005
R7555 VSS.n6531 VSS.n6535 4.57324
R7556 VSS.n6527 VSS.n6525 0.147342
R7557 VSS.n6528 VSS.n6529 0.0732424
R7558 VSS.n6529 VSS.n6530 0.147342
R7559 VSS.n6532 VSS.n6536 0.0721009
R7560 VSS.n6537 VSS.n6533 4.5005
R7561 VSS.n6538 VSS.n6534 4.5005
R7562 VSS.n6539 VSS.n6535 4.5005
R7563 VSS.n6525 VSS.n6536 4.57442
R7564 VSS.n6532 VSS.n6533 0.147342
R7565 VSS.n6533 VSS.n6534 0.147342
R7566 VSS.n6534 VSS.n6535 0.147342
R7567 VSS.n6536 VSS.n6537 2.39784
R7568 VSS.n6537 VSS.n6538 0.147342
R7569 VSS.n6538 VSS.n6539 0.147342
R7570 VSS.n6539 VSS.t548 3.13212
R7571 VSS.n6512 VSS.n6517 4.5005
R7572 VSS.n6514 VSS.n6518 4.5005
R7573 VSS.n6515 VSS.n6519 4.5005
R7574 VSS.n6516 VSS.n6520 4.57324
R7575 VSS.n6512 VSS.n6510 0.147342
R7576 VSS.n6513 VSS.n6514 0.0732424
R7577 VSS.n6514 VSS.n6515 0.147342
R7578 VSS.n6517 VSS.n6521 0.0721009
R7579 VSS.n6522 VSS.n6518 4.5005
R7580 VSS.n6523 VSS.n6519 4.5005
R7581 VSS.n6524 VSS.n6520 4.5005
R7582 VSS.n6510 VSS.n6521 4.57442
R7583 VSS.n6517 VSS.n6518 0.147342
R7584 VSS.n6518 VSS.n6519 0.147342
R7585 VSS.n6519 VSS.n6520 0.147342
R7586 VSS.n6521 VSS.n6522 2.39784
R7587 VSS.n6522 VSS.n6523 0.147342
R7588 VSS.n6523 VSS.n6524 0.147342
R7589 VSS.n6524 VSS.t256 3.13212
R7590 VSS.n6497 VSS.n6502 4.5005
R7591 VSS.n6499 VSS.n6503 4.5005
R7592 VSS.n6500 VSS.n6504 4.5005
R7593 VSS.n6501 VSS.n6505 4.57324
R7594 VSS.n6497 VSS.n6495 0.147342
R7595 VSS.n6498 VSS.n6499 0.0732424
R7596 VSS.n6499 VSS.n6500 0.147342
R7597 VSS.n6502 VSS.n6506 0.0721009
R7598 VSS.n6507 VSS.n6503 4.5005
R7599 VSS.n6508 VSS.n6504 4.5005
R7600 VSS.n6509 VSS.n6505 4.5005
R7601 VSS.n6495 VSS.n6506 4.57442
R7602 VSS.n6502 VSS.n6503 0.147342
R7603 VSS.n6503 VSS.n6504 0.147342
R7604 VSS.n6504 VSS.n6505 0.147342
R7605 VSS.n6506 VSS.n6507 2.39784
R7606 VSS.n6507 VSS.n6508 0.147342
R7607 VSS.n6508 VSS.n6509 0.147342
R7608 VSS.n6509 VSS.t435 3.13212
R7609 VSS.n6487 VSS.n6482 4.5005
R7610 VSS.n6488 VSS.n6484 4.5005
R7611 VSS.n6489 VSS.n6485 4.5005
R7612 VSS.n6490 VSS.n6486 4.57324
R7613 VSS.n6480 VSS.n6482 0.147342
R7614 VSS.n6483 VSS.n6484 0.0732424
R7615 VSS.n6484 VSS.n6485 0.147342
R7616 VSS.n6491 VSS.n6487 0.0722544
R7617 VSS.n6492 VSS.n6488 4.5005
R7618 VSS.n6493 VSS.n6489 4.5005
R7619 VSS.n6494 VSS.n6490 4.5005
R7620 VSS.n6491 VSS.n6480 4.57426
R7621 VSS.n6487 VSS.n6488 0.147342
R7622 VSS.n6488 VSS.n6489 0.147342
R7623 VSS.n6489 VSS.n6490 0.147342
R7624 VSS.n6492 VSS.n6491 2.37296
R7625 VSS.n6493 VSS.n6492 0.127318
R7626 VSS.n6494 VSS.n6493 0.127318
R7627 VSS.t0 VSS.n6494 2.73618
R7628 VSS.n6467 VSS.n6472 4.5005
R7629 VSS.n6469 VSS.n6473 4.5005
R7630 VSS.n6470 VSS.n6474 4.5005
R7631 VSS.n6471 VSS.n6475 4.57324
R7632 VSS.n6467 VSS.n6465 0.147342
R7633 VSS.n6468 VSS.n6469 0.0732424
R7634 VSS.n6469 VSS.n6470 0.147342
R7635 VSS.n6472 VSS.n6476 0.0721009
R7636 VSS.n6477 VSS.n6473 4.5005
R7637 VSS.n6478 VSS.n6474 4.5005
R7638 VSS.n6479 VSS.n6475 4.5005
R7639 VSS.n6465 VSS.n6476 4.57442
R7640 VSS.n6472 VSS.n6473 0.147342
R7641 VSS.n6473 VSS.n6474 0.147342
R7642 VSS.n6474 VSS.n6475 0.147342
R7643 VSS.n6476 VSS.n6477 2.39784
R7644 VSS.n6477 VSS.n6478 0.147342
R7645 VSS.n6478 VSS.n6479 0.147342
R7646 VSS.n6479 VSS.t3 3.13212
R7647 VSS.n6452 VSS.n6457 4.5005
R7648 VSS.n6454 VSS.n6458 4.5005
R7649 VSS.n6455 VSS.n6459 4.5005
R7650 VSS.n6456 VSS.n6460 4.57324
R7651 VSS.n6452 VSS.n6450 0.147342
R7652 VSS.n6453 VSS.n6454 0.0732424
R7653 VSS.n6454 VSS.n6455 0.147342
R7654 VSS.n6457 VSS.n6461 0.0721009
R7655 VSS.n6462 VSS.n6458 4.5005
R7656 VSS.n6463 VSS.n6459 4.5005
R7657 VSS.n6464 VSS.n6460 4.5005
R7658 VSS.n6450 VSS.n6461 4.57442
R7659 VSS.n6457 VSS.n6458 0.147342
R7660 VSS.n6458 VSS.n6459 0.147342
R7661 VSS.n6459 VSS.n6460 0.147342
R7662 VSS.n6461 VSS.n6462 2.39784
R7663 VSS.n6462 VSS.n6463 0.147342
R7664 VSS.n6463 VSS.n6464 0.147342
R7665 VSS.n6464 VSS.t407 3.13212
R7666 VSS.n6437 VSS.n6442 4.5005
R7667 VSS.n6439 VSS.n6443 4.5005
R7668 VSS.n6440 VSS.n6444 4.5005
R7669 VSS.n6441 VSS.n6445 4.57324
R7670 VSS.n6437 VSS.n6435 0.147342
R7671 VSS.n6438 VSS.n6439 0.0732424
R7672 VSS.n6439 VSS.n6440 0.147342
R7673 VSS.n6442 VSS.n6446 0.0721009
R7674 VSS.n6447 VSS.n6443 4.5005
R7675 VSS.n6448 VSS.n6444 4.5005
R7676 VSS.n6449 VSS.n6445 4.5005
R7677 VSS.n6435 VSS.n6446 4.57442
R7678 VSS.n6442 VSS.n6443 0.147342
R7679 VSS.n6443 VSS.n6444 0.147342
R7680 VSS.n6444 VSS.n6445 0.147342
R7681 VSS.n6446 VSS.n6447 2.39784
R7682 VSS.n6447 VSS.n6448 0.147342
R7683 VSS.n6448 VSS.n6449 0.147342
R7684 VSS.n6449 VSS.t260 3.13212
R7685 VSS.n6422 VSS.n6427 4.5005
R7686 VSS.n6424 VSS.n6428 4.5005
R7687 VSS.n6425 VSS.n6429 4.5005
R7688 VSS.n6426 VSS.n6430 4.57324
R7689 VSS.n6422 VSS.n6420 0.147342
R7690 VSS.n6423 VSS.n6424 0.0732424
R7691 VSS.n6424 VSS.n6425 0.147342
R7692 VSS.n6427 VSS.n6431 0.0721009
R7693 VSS.n6432 VSS.n6428 4.5005
R7694 VSS.n6433 VSS.n6429 4.5005
R7695 VSS.n6434 VSS.n6430 4.5005
R7696 VSS.n6420 VSS.n6431 4.57442
R7697 VSS.n6427 VSS.n6428 0.147342
R7698 VSS.n6428 VSS.n6429 0.147342
R7699 VSS.n6429 VSS.n6430 0.147342
R7700 VSS.n6431 VSS.n6432 2.39784
R7701 VSS.n6432 VSS.n6433 0.147342
R7702 VSS.n6433 VSS.n6434 0.147342
R7703 VSS.n6434 VSS.t268 3.13212
R7704 VSS.n6407 VSS.n6412 4.5005
R7705 VSS.n6409 VSS.n6413 4.5005
R7706 VSS.n6410 VSS.n6414 4.5005
R7707 VSS.n6411 VSS.n6415 4.57324
R7708 VSS.n6407 VSS.n6405 0.147342
R7709 VSS.n6408 VSS.n6409 0.0732424
R7710 VSS.n6409 VSS.n6410 0.147342
R7711 VSS.n6412 VSS.n6416 0.0721009
R7712 VSS.n6417 VSS.n6413 4.5005
R7713 VSS.n6418 VSS.n6414 4.5005
R7714 VSS.n6419 VSS.n6415 4.5005
R7715 VSS.n6405 VSS.n6416 4.57442
R7716 VSS.n6412 VSS.n6413 0.147342
R7717 VSS.n6413 VSS.n6414 0.147342
R7718 VSS.n6414 VSS.n6415 0.147342
R7719 VSS.n6416 VSS.n6417 2.39784
R7720 VSS.n6417 VSS.n6418 0.147342
R7721 VSS.n6418 VSS.n6419 0.147342
R7722 VSS.n6419 VSS.t480 3.13212
R7723 VSS.n6392 VSS.n6397 4.5005
R7724 VSS.n6394 VSS.n6398 4.5005
R7725 VSS.n6395 VSS.n6399 4.5005
R7726 VSS.n6396 VSS.n6400 4.57324
R7727 VSS.n6392 VSS.n6390 0.147342
R7728 VSS.n6393 VSS.n6394 0.0732424
R7729 VSS.n6394 VSS.n6395 0.147342
R7730 VSS.n6397 VSS.n6401 0.0721009
R7731 VSS.n6402 VSS.n6398 4.5005
R7732 VSS.n6403 VSS.n6399 4.5005
R7733 VSS.n6404 VSS.n6400 4.5005
R7734 VSS.n6390 VSS.n6401 4.57442
R7735 VSS.n6397 VSS.n6398 0.147342
R7736 VSS.n6398 VSS.n6399 0.147342
R7737 VSS.n6399 VSS.n6400 0.147342
R7738 VSS.n6401 VSS.n6402 2.39784
R7739 VSS.n6402 VSS.n6403 0.147342
R7740 VSS.n6403 VSS.n6404 0.147342
R7741 VSS.n6404 VSS.t62 3.13212
R7742 VSS.n6382 VSS.n6377 4.5005
R7743 VSS.n6383 VSS.n6379 4.5005
R7744 VSS.n6384 VSS.n6380 4.5005
R7745 VSS.n6385 VSS.n6381 4.57324
R7746 VSS.n6375 VSS.n6377 0.147342
R7747 VSS.n6378 VSS.n6379 0.0732424
R7748 VSS.n6379 VSS.n6380 0.147342
R7749 VSS.n6386 VSS.n6382 0.0722544
R7750 VSS.n6387 VSS.n6383 4.5005
R7751 VSS.n6388 VSS.n6384 4.5005
R7752 VSS.n6389 VSS.n6385 4.5005
R7753 VSS.n6386 VSS.n6375 4.57426
R7754 VSS.n6382 VSS.n6383 0.147342
R7755 VSS.n6383 VSS.n6384 0.147342
R7756 VSS.n6384 VSS.n6385 0.147342
R7757 VSS.n6387 VSS.n6386 2.37296
R7758 VSS.n6388 VSS.n6387 0.127318
R7759 VSS.n6389 VSS.n6388 0.127318
R7760 VSS.t0 VSS.n6389 2.73618
R7761 VSS.n6362 VSS.n6367 4.5005
R7762 VSS.n6364 VSS.n6368 4.5005
R7763 VSS.n6365 VSS.n6369 4.5005
R7764 VSS.n6366 VSS.n6370 4.57324
R7765 VSS.n6362 VSS.n6360 0.147342
R7766 VSS.n6363 VSS.n6364 0.0732424
R7767 VSS.n6364 VSS.n6365 0.147342
R7768 VSS.n6367 VSS.n6371 0.0721009
R7769 VSS.n6372 VSS.n6368 4.5005
R7770 VSS.n6373 VSS.n6369 4.5005
R7771 VSS.n6374 VSS.n6370 4.5005
R7772 VSS.n6360 VSS.n6371 4.57442
R7773 VSS.n6367 VSS.n6368 0.147342
R7774 VSS.n6368 VSS.n6369 0.147342
R7775 VSS.n6369 VSS.n6370 0.147342
R7776 VSS.n6371 VSS.n6372 2.39784
R7777 VSS.n6372 VSS.n6373 0.147342
R7778 VSS.n6373 VSS.n6374 0.147342
R7779 VSS.n6374 VSS.t217 3.13212
R7780 VSS.n6347 VSS.n6352 4.5005
R7781 VSS.n6349 VSS.n6353 4.5005
R7782 VSS.n6350 VSS.n6354 4.5005
R7783 VSS.n6351 VSS.n6355 4.57324
R7784 VSS.n6347 VSS.n6345 0.147342
R7785 VSS.n6348 VSS.n6349 0.0732424
R7786 VSS.n6349 VSS.n6350 0.147342
R7787 VSS.n6352 VSS.n6356 0.0721009
R7788 VSS.n6357 VSS.n6353 4.5005
R7789 VSS.n6358 VSS.n6354 4.5005
R7790 VSS.n6359 VSS.n6355 4.5005
R7791 VSS.n6345 VSS.n6356 4.57442
R7792 VSS.n6352 VSS.n6353 0.147342
R7793 VSS.n6353 VSS.n6354 0.147342
R7794 VSS.n6354 VSS.n6355 0.147342
R7795 VSS.n6356 VSS.n6357 2.39784
R7796 VSS.n6357 VSS.n6358 0.147342
R7797 VSS.n6358 VSS.n6359 0.147342
R7798 VSS.n6359 VSS.t103 3.13212
R7799 VSS.n6332 VSS.n6337 4.5005
R7800 VSS.n6334 VSS.n6338 4.5005
R7801 VSS.n6335 VSS.n6339 4.5005
R7802 VSS.n6336 VSS.n6340 4.57324
R7803 VSS.n6332 VSS.n6330 0.147342
R7804 VSS.n6333 VSS.n6334 0.0732424
R7805 VSS.n6334 VSS.n6335 0.147342
R7806 VSS.n6337 VSS.n6341 0.0721009
R7807 VSS.n6342 VSS.n6338 4.5005
R7808 VSS.n6343 VSS.n6339 4.5005
R7809 VSS.n6344 VSS.n6340 4.5005
R7810 VSS.n6330 VSS.n6341 4.57442
R7811 VSS.n6337 VSS.n6338 0.147342
R7812 VSS.n6338 VSS.n6339 0.147342
R7813 VSS.n6339 VSS.n6340 0.147342
R7814 VSS.n6341 VSS.n6342 2.39784
R7815 VSS.n6342 VSS.n6343 0.147342
R7816 VSS.n6343 VSS.n6344 0.147342
R7817 VSS.n6344 VSS.t132 3.13212
R7818 VSS.n6322 VSS.n6317 4.5005
R7819 VSS.n6323 VSS.n6319 4.5005
R7820 VSS.n6324 VSS.n6320 4.5005
R7821 VSS.n6325 VSS.n6321 4.57324
R7822 VSS.n6315 VSS.n6317 0.147342
R7823 VSS.n6318 VSS.n6319 0.0732424
R7824 VSS.n6319 VSS.n6320 0.147342
R7825 VSS.n6326 VSS.n6322 0.0722544
R7826 VSS.n6327 VSS.n6323 4.5005
R7827 VSS.n6328 VSS.n6324 4.5005
R7828 VSS.n6329 VSS.n6325 4.5005
R7829 VSS.n6326 VSS.n6315 4.57426
R7830 VSS.n6322 VSS.n6323 0.147342
R7831 VSS.n6323 VSS.n6324 0.147342
R7832 VSS.n6324 VSS.n6325 0.147342
R7833 VSS.n6327 VSS.n6326 2.37296
R7834 VSS.n6328 VSS.n6327 0.127318
R7835 VSS.n6329 VSS.n6328 0.127318
R7836 VSS.t0 VSS.n6329 2.73618
R7837 VSS.n6302 VSS.n6307 4.5005
R7838 VSS.n6304 VSS.n6308 4.5005
R7839 VSS.n6305 VSS.n6309 4.5005
R7840 VSS.n6306 VSS.n6310 4.57324
R7841 VSS.n6302 VSS.n6300 0.147342
R7842 VSS.n6303 VSS.n6304 0.0732424
R7843 VSS.n6304 VSS.n6305 0.147342
R7844 VSS.n6307 VSS.n6311 0.0721009
R7845 VSS.n6312 VSS.n6308 4.5005
R7846 VSS.n6313 VSS.n6309 4.5005
R7847 VSS.n6314 VSS.n6310 4.5005
R7848 VSS.n6300 VSS.n6311 4.57442
R7849 VSS.n6307 VSS.n6308 0.147342
R7850 VSS.n6308 VSS.n6309 0.147342
R7851 VSS.n6309 VSS.n6310 0.147342
R7852 VSS.n6311 VSS.n6312 2.39784
R7853 VSS.n6312 VSS.n6313 0.147342
R7854 VSS.n6313 VSS.n6314 0.147342
R7855 VSS.n6314 VSS.t133 3.13212
R7856 VSS.n6287 VSS.n6292 4.5005
R7857 VSS.n6289 VSS.n6293 4.5005
R7858 VSS.n6290 VSS.n6294 4.5005
R7859 VSS.n6291 VSS.n6295 4.57324
R7860 VSS.n6287 VSS.n6285 0.147342
R7861 VSS.n6288 VSS.n6289 0.0732424
R7862 VSS.n6289 VSS.n6290 0.147342
R7863 VSS.n6292 VSS.n6296 0.0721009
R7864 VSS.n6297 VSS.n6293 4.5005
R7865 VSS.n6298 VSS.n6294 4.5005
R7866 VSS.n6299 VSS.n6295 4.5005
R7867 VSS.n6285 VSS.n6296 4.57442
R7868 VSS.n6292 VSS.n6293 0.147342
R7869 VSS.n6293 VSS.n6294 0.147342
R7870 VSS.n6294 VSS.n6295 0.147342
R7871 VSS.n6296 VSS.n6297 2.39784
R7872 VSS.n6297 VSS.n6298 0.147342
R7873 VSS.n6298 VSS.n6299 0.147342
R7874 VSS.n6299 VSS.t102 3.13212
R7875 VSS.n6272 VSS.n6277 4.5005
R7876 VSS.n6274 VSS.n6278 4.5005
R7877 VSS.n6275 VSS.n6279 4.5005
R7878 VSS.n6276 VSS.n6280 4.57324
R7879 VSS.n6272 VSS.n6270 0.147342
R7880 VSS.n6273 VSS.n6274 0.0732424
R7881 VSS.n6274 VSS.n6275 0.147342
R7882 VSS.n6277 VSS.n6281 0.0721009
R7883 VSS.n6282 VSS.n6278 4.5005
R7884 VSS.n6283 VSS.n6279 4.5005
R7885 VSS.n6284 VSS.n6280 4.5005
R7886 VSS.n6270 VSS.n6281 4.57442
R7887 VSS.n6277 VSS.n6278 0.147342
R7888 VSS.n6278 VSS.n6279 0.147342
R7889 VSS.n6279 VSS.n6280 0.147342
R7890 VSS.n6281 VSS.n6282 2.39784
R7891 VSS.n6282 VSS.n6283 0.147342
R7892 VSS.n6283 VSS.n6284 0.147342
R7893 VSS.n6284 VSS.t285 3.13212
R7894 VSS.n6257 VSS.n6262 4.5005
R7895 VSS.n6259 VSS.n6263 4.5005
R7896 VSS.n6260 VSS.n6264 4.5005
R7897 VSS.n6261 VSS.n6265 4.57324
R7898 VSS.n6257 VSS.n6255 0.147342
R7899 VSS.n6258 VSS.n6259 0.0732424
R7900 VSS.n6259 VSS.n6260 0.147342
R7901 VSS.n6262 VSS.n6266 0.0721009
R7902 VSS.n6267 VSS.n6263 4.5005
R7903 VSS.n6268 VSS.n6264 4.5005
R7904 VSS.n6269 VSS.n6265 4.5005
R7905 VSS.n6255 VSS.n6266 4.57442
R7906 VSS.n6262 VSS.n6263 0.147342
R7907 VSS.n6263 VSS.n6264 0.147342
R7908 VSS.n6264 VSS.n6265 0.147342
R7909 VSS.n6266 VSS.n6267 2.39784
R7910 VSS.n6267 VSS.n6268 0.147342
R7911 VSS.n6268 VSS.n6269 0.147342
R7912 VSS.n6269 VSS.t295 3.13212
R7913 VSS.n6247 VSS.n6242 4.5005
R7914 VSS.n6248 VSS.n6244 4.5005
R7915 VSS.n6249 VSS.n6245 4.5005
R7916 VSS.n6250 VSS.n6246 4.57324
R7917 VSS.n6240 VSS.n6242 0.147342
R7918 VSS.n6243 VSS.n6244 0.0732424
R7919 VSS.n6244 VSS.n6245 0.147342
R7920 VSS.n6251 VSS.n6247 0.0722544
R7921 VSS.n6252 VSS.n6248 4.5005
R7922 VSS.n6253 VSS.n6249 4.5005
R7923 VSS.n6254 VSS.n6250 4.5005
R7924 VSS.n6251 VSS.n6240 4.57426
R7925 VSS.n6247 VSS.n6248 0.147342
R7926 VSS.n6248 VSS.n6249 0.147342
R7927 VSS.n6249 VSS.n6250 0.147342
R7928 VSS.n6252 VSS.n6251 2.37296
R7929 VSS.n6253 VSS.n6252 0.127318
R7930 VSS.n6254 VSS.n6253 0.127318
R7931 VSS.t0 VSS.n6254 2.73618
R7932 VSS.n6227 VSS.n6232 4.5005
R7933 VSS.n6229 VSS.n6233 4.5005
R7934 VSS.n6230 VSS.n6234 4.5005
R7935 VSS.n6231 VSS.n6235 4.57324
R7936 VSS.n6227 VSS.n6225 0.147342
R7937 VSS.n6228 VSS.n6229 0.0732424
R7938 VSS.n6229 VSS.n6230 0.147342
R7939 VSS.n6232 VSS.n6236 0.0721009
R7940 VSS.n6237 VSS.n6233 4.5005
R7941 VSS.n6238 VSS.n6234 4.5005
R7942 VSS.n6239 VSS.n6235 4.5005
R7943 VSS.n6225 VSS.n6236 4.57442
R7944 VSS.n6232 VSS.n6233 0.147342
R7945 VSS.n6233 VSS.n6234 0.147342
R7946 VSS.n6234 VSS.n6235 0.147342
R7947 VSS.n6236 VSS.n6237 2.39784
R7948 VSS.n6237 VSS.n6238 0.147342
R7949 VSS.n6238 VSS.n6239 0.147342
R7950 VSS.n6239 VSS.t542 3.13212
R7951 VSS.n6212 VSS.n6217 4.5005
R7952 VSS.n6214 VSS.n6218 4.5005
R7953 VSS.n6215 VSS.n6219 4.5005
R7954 VSS.n6216 VSS.n6220 4.57324
R7955 VSS.n6212 VSS.n6210 0.147342
R7956 VSS.n6213 VSS.n6214 0.0732424
R7957 VSS.n6214 VSS.n6215 0.147342
R7958 VSS.n6217 VSS.n6221 0.0721009
R7959 VSS.n6222 VSS.n6218 4.5005
R7960 VSS.n6223 VSS.n6219 4.5005
R7961 VSS.n6224 VSS.n6220 4.5005
R7962 VSS.n6210 VSS.n6221 4.57442
R7963 VSS.n6217 VSS.n6218 0.147342
R7964 VSS.n6218 VSS.n6219 0.147342
R7965 VSS.n6219 VSS.n6220 0.147342
R7966 VSS.n6221 VSS.n6222 2.39784
R7967 VSS.n6222 VSS.n6223 0.147342
R7968 VSS.n6223 VSS.n6224 0.147342
R7969 VSS.n6224 VSS.t278 3.13212
R7970 VSS.n6197 VSS.n6202 4.5005
R7971 VSS.n6199 VSS.n6203 4.5005
R7972 VSS.n6200 VSS.n6204 4.5005
R7973 VSS.n6201 VSS.n6205 4.57324
R7974 VSS.n6197 VSS.n6195 0.147342
R7975 VSS.n6198 VSS.n6199 0.0732424
R7976 VSS.n6199 VSS.n6200 0.147342
R7977 VSS.n6202 VSS.n6206 0.0721009
R7978 VSS.n6207 VSS.n6203 4.5005
R7979 VSS.n6208 VSS.n6204 4.5005
R7980 VSS.n6209 VSS.n6205 4.5005
R7981 VSS.n6195 VSS.n6206 4.57442
R7982 VSS.n6202 VSS.n6203 0.147342
R7983 VSS.n6203 VSS.n6204 0.147342
R7984 VSS.n6204 VSS.n6205 0.147342
R7985 VSS.n6206 VSS.n6207 2.39784
R7986 VSS.n6207 VSS.n6208 0.147342
R7987 VSS.n6208 VSS.n6209 0.147342
R7988 VSS.n6209 VSS.t439 3.13212
R7989 VSS.n6187 VSS.n6182 4.5005
R7990 VSS.n6188 VSS.n6184 4.5005
R7991 VSS.n6189 VSS.n6185 4.5005
R7992 VSS.n6190 VSS.n6186 4.57324
R7993 VSS.n6180 VSS.n6182 0.147342
R7994 VSS.n6183 VSS.n6184 0.0732424
R7995 VSS.n6184 VSS.n6185 0.147342
R7996 VSS.n6191 VSS.n6187 0.0722544
R7997 VSS.n6192 VSS.n6188 4.5005
R7998 VSS.n6193 VSS.n6189 4.5005
R7999 VSS.n6194 VSS.n6190 4.5005
R8000 VSS.n6191 VSS.n6180 4.57426
R8001 VSS.n6187 VSS.n6188 0.147342
R8002 VSS.n6188 VSS.n6189 0.147342
R8003 VSS.n6189 VSS.n6190 0.147342
R8004 VSS.n6192 VSS.n6191 2.37296
R8005 VSS.n6193 VSS.n6192 0.127318
R8006 VSS.n6194 VSS.n6193 0.127318
R8007 VSS.t0 VSS.n6194 2.73618
R8008 VSS.n6167 VSS.n6172 4.5005
R8009 VSS.n6169 VSS.n6173 4.5005
R8010 VSS.n6170 VSS.n6174 4.5005
R8011 VSS.n6171 VSS.n6175 4.57324
R8012 VSS.n6167 VSS.n6165 0.147342
R8013 VSS.n6168 VSS.n6169 0.0732424
R8014 VSS.n6169 VSS.n6170 0.147342
R8015 VSS.n6172 VSS.n6176 0.0721009
R8016 VSS.n6177 VSS.n6173 4.5005
R8017 VSS.n6178 VSS.n6174 4.5005
R8018 VSS.n6179 VSS.n6175 4.5005
R8019 VSS.n6165 VSS.n6176 4.57442
R8020 VSS.n6172 VSS.n6173 0.147342
R8021 VSS.n6173 VSS.n6174 0.147342
R8022 VSS.n6174 VSS.n6175 0.147342
R8023 VSS.n6176 VSS.n6177 2.39784
R8024 VSS.n6177 VSS.n6178 0.147342
R8025 VSS.n6178 VSS.n6179 0.147342
R8026 VSS.n6179 VSS.t444 3.13212
R8027 VSS.n6152 VSS.n6157 4.5005
R8028 VSS.n6154 VSS.n6158 4.5005
R8029 VSS.n6155 VSS.n6159 4.5005
R8030 VSS.n6156 VSS.n6160 4.57324
R8031 VSS.n6152 VSS.n6150 0.147342
R8032 VSS.n6153 VSS.n6154 0.0732424
R8033 VSS.n6154 VSS.n6155 0.147342
R8034 VSS.n6157 VSS.n6161 0.0721009
R8035 VSS.n6162 VSS.n6158 4.5005
R8036 VSS.n6163 VSS.n6159 4.5005
R8037 VSS.n6164 VSS.n6160 4.5005
R8038 VSS.n6150 VSS.n6161 4.57442
R8039 VSS.n6157 VSS.n6158 0.147342
R8040 VSS.n6158 VSS.n6159 0.147342
R8041 VSS.n6159 VSS.n6160 0.147342
R8042 VSS.n6161 VSS.n6162 2.39784
R8043 VSS.n6162 VSS.n6163 0.147342
R8044 VSS.n6163 VSS.n6164 0.147342
R8045 VSS.n6164 VSS.t408 3.13212
R8046 VSS.n6137 VSS.n6142 4.5005
R8047 VSS.n6139 VSS.n6143 4.5005
R8048 VSS.n6140 VSS.n6144 4.5005
R8049 VSS.n6141 VSS.n6145 4.57324
R8050 VSS.n6137 VSS.n6135 0.147342
R8051 VSS.n6138 VSS.n6139 0.0732424
R8052 VSS.n6139 VSS.n6140 0.147342
R8053 VSS.n6142 VSS.n6146 0.0721009
R8054 VSS.n6147 VSS.n6143 4.5005
R8055 VSS.n6148 VSS.n6144 4.5005
R8056 VSS.n6149 VSS.n6145 4.5005
R8057 VSS.n6135 VSS.n6146 4.57442
R8058 VSS.n6142 VSS.n6143 0.147342
R8059 VSS.n6143 VSS.n6144 0.147342
R8060 VSS.n6144 VSS.n6145 0.147342
R8061 VSS.n6146 VSS.n6147 2.39784
R8062 VSS.n6147 VSS.n6148 0.147342
R8063 VSS.n6148 VSS.n6149 0.147342
R8064 VSS.n6149 VSS.t261 3.13212
R8065 VSS.n6122 VSS.n6127 4.5005
R8066 VSS.n6124 VSS.n6128 4.5005
R8067 VSS.n6125 VSS.n6129 4.5005
R8068 VSS.n6126 VSS.n6130 4.57324
R8069 VSS.n6122 VSS.n6120 0.147342
R8070 VSS.n6123 VSS.n6124 0.0732424
R8071 VSS.n6124 VSS.n6125 0.147342
R8072 VSS.n6127 VSS.n6131 0.0721009
R8073 VSS.n6132 VSS.n6128 4.5005
R8074 VSS.n6133 VSS.n6129 4.5005
R8075 VSS.n6134 VSS.n6130 4.5005
R8076 VSS.n6120 VSS.n6131 4.57442
R8077 VSS.n6127 VSS.n6128 0.147342
R8078 VSS.n6128 VSS.n6129 0.147342
R8079 VSS.n6129 VSS.n6130 0.147342
R8080 VSS.n6131 VSS.n6132 2.39784
R8081 VSS.n6132 VSS.n6133 0.147342
R8082 VSS.n6133 VSS.n6134 0.147342
R8083 VSS.n6134 VSS.t96 3.13212
R8084 VSS.n6107 VSS.n6112 4.5005
R8085 VSS.n6109 VSS.n6113 4.5005
R8086 VSS.n6110 VSS.n6114 4.5005
R8087 VSS.n6111 VSS.n6115 4.57324
R8088 VSS.n6107 VSS.n6105 0.147342
R8089 VSS.n6108 VSS.n6109 0.0732424
R8090 VSS.n6109 VSS.n6110 0.147342
R8091 VSS.n6112 VSS.n6116 0.0721009
R8092 VSS.n6117 VSS.n6113 4.5005
R8093 VSS.n6118 VSS.n6114 4.5005
R8094 VSS.n6119 VSS.n6115 4.5005
R8095 VSS.n6105 VSS.n6116 4.57442
R8096 VSS.n6112 VSS.n6113 0.147342
R8097 VSS.n6113 VSS.n6114 0.147342
R8098 VSS.n6114 VSS.n6115 0.147342
R8099 VSS.n6116 VSS.n6117 2.39784
R8100 VSS.n6117 VSS.n6118 0.147342
R8101 VSS.n6118 VSS.n6119 0.147342
R8102 VSS.n6119 VSS.t470 3.13212
R8103 VSS.n6092 VSS.n6097 4.5005
R8104 VSS.n6094 VSS.n6098 4.5005
R8105 VSS.n6095 VSS.n6099 4.5005
R8106 VSS.n6096 VSS.n6100 4.57324
R8107 VSS.n6092 VSS.n6090 0.147342
R8108 VSS.n6093 VSS.n6094 0.0732424
R8109 VSS.n6094 VSS.n6095 0.147342
R8110 VSS.n6097 VSS.n6101 0.0721009
R8111 VSS.n6102 VSS.n6098 4.5005
R8112 VSS.n6103 VSS.n6099 4.5005
R8113 VSS.n6104 VSS.n6100 4.5005
R8114 VSS.n6090 VSS.n6101 4.57442
R8115 VSS.n6097 VSS.n6098 0.147342
R8116 VSS.n6098 VSS.n6099 0.147342
R8117 VSS.n6099 VSS.n6100 0.147342
R8118 VSS.n6101 VSS.n6102 2.39784
R8119 VSS.n6102 VSS.n6103 0.147342
R8120 VSS.n6103 VSS.n6104 0.147342
R8121 VSS.n6104 VSS.t512 3.13212
R8122 VSS.n6082 VSS.n6077 4.5005
R8123 VSS.n6083 VSS.n6079 4.5005
R8124 VSS.n6084 VSS.n6080 4.5005
R8125 VSS.n6085 VSS.n6081 4.57324
R8126 VSS.n6075 VSS.n6077 0.147342
R8127 VSS.n6078 VSS.n6079 0.0732424
R8128 VSS.n6079 VSS.n6080 0.147342
R8129 VSS.n6086 VSS.n6082 0.0722544
R8130 VSS.n6087 VSS.n6083 4.5005
R8131 VSS.n6088 VSS.n6084 4.5005
R8132 VSS.n6089 VSS.n6085 4.5005
R8133 VSS.n6086 VSS.n6075 4.57426
R8134 VSS.n6082 VSS.n6083 0.147342
R8135 VSS.n6083 VSS.n6084 0.147342
R8136 VSS.n6084 VSS.n6085 0.147342
R8137 VSS.n6087 VSS.n6086 2.37296
R8138 VSS.n6088 VSS.n6087 0.127318
R8139 VSS.n6089 VSS.n6088 0.127318
R8140 VSS.t0 VSS.n6089 2.73618
R8141 VSS.n6062 VSS.n6067 4.5005
R8142 VSS.n6064 VSS.n6068 4.5005
R8143 VSS.n6065 VSS.n6069 4.5005
R8144 VSS.n6066 VSS.n6070 4.57324
R8145 VSS.n6062 VSS.n6060 0.147342
R8146 VSS.n6063 VSS.n6064 0.0732424
R8147 VSS.n6064 VSS.n6065 0.147342
R8148 VSS.n6067 VSS.n6071 0.0721009
R8149 VSS.n6072 VSS.n6068 4.5005
R8150 VSS.n6073 VSS.n6069 4.5005
R8151 VSS.n6074 VSS.n6070 4.5005
R8152 VSS.n6060 VSS.n6071 4.57442
R8153 VSS.n6067 VSS.n6068 0.147342
R8154 VSS.n6068 VSS.n6069 0.147342
R8155 VSS.n6069 VSS.n6070 0.147342
R8156 VSS.n6071 VSS.n6072 2.39784
R8157 VSS.n6072 VSS.n6073 0.147342
R8158 VSS.n6073 VSS.n6074 0.147342
R8159 VSS.n6074 VSS.t213 3.13212
R8160 VSS.n6047 VSS.n6052 4.5005
R8161 VSS.n6049 VSS.n6053 4.5005
R8162 VSS.n6050 VSS.n6054 4.5005
R8163 VSS.n6051 VSS.n6055 4.57324
R8164 VSS.n6047 VSS.n6045 0.147342
R8165 VSS.n6048 VSS.n6049 0.0732424
R8166 VSS.n6049 VSS.n6050 0.147342
R8167 VSS.n6052 VSS.n6056 0.0721009
R8168 VSS.n6057 VSS.n6053 4.5005
R8169 VSS.n6058 VSS.n6054 4.5005
R8170 VSS.n6059 VSS.n6055 4.5005
R8171 VSS.n6045 VSS.n6056 4.57442
R8172 VSS.n6052 VSS.n6053 0.147342
R8173 VSS.n6053 VSS.n6054 0.147342
R8174 VSS.n6054 VSS.n6055 0.147342
R8175 VSS.n6056 VSS.n6057 2.39784
R8176 VSS.n6057 VSS.n6058 0.147342
R8177 VSS.n6058 VSS.n6059 0.147342
R8178 VSS.n6059 VSS.t104 3.13212
R8179 VSS.n6032 VSS.n6037 4.5005
R8180 VSS.n6034 VSS.n6038 4.5005
R8181 VSS.n6035 VSS.n6039 4.5005
R8182 VSS.n6036 VSS.n6040 4.57324
R8183 VSS.n6032 VSS.n6030 0.147342
R8184 VSS.n6033 VSS.n6034 0.0732424
R8185 VSS.n6034 VSS.n6035 0.147342
R8186 VSS.n6037 VSS.n6041 0.0721009
R8187 VSS.n6042 VSS.n6038 4.5005
R8188 VSS.n6043 VSS.n6039 4.5005
R8189 VSS.n6044 VSS.n6040 4.5005
R8190 VSS.n6030 VSS.n6041 4.57442
R8191 VSS.n6037 VSS.n6038 0.147342
R8192 VSS.n6038 VSS.n6039 0.147342
R8193 VSS.n6039 VSS.n6040 0.147342
R8194 VSS.n6041 VSS.n6042 2.39784
R8195 VSS.n6042 VSS.n6043 0.147342
R8196 VSS.n6043 VSS.n6044 0.147342
R8197 VSS.n6044 VSS.t237 3.13212
R8198 VSS.n6022 VSS.n6017 4.5005
R8199 VSS.n6023 VSS.n6019 4.5005
R8200 VSS.n6024 VSS.n6020 4.5005
R8201 VSS.n6025 VSS.n6021 4.57324
R8202 VSS.n6015 VSS.n6017 0.147342
R8203 VSS.n6018 VSS.n6019 0.0732424
R8204 VSS.n6019 VSS.n6020 0.147342
R8205 VSS.n6026 VSS.n6022 0.0722544
R8206 VSS.n6027 VSS.n6023 4.5005
R8207 VSS.n6028 VSS.n6024 4.5005
R8208 VSS.n6029 VSS.n6025 4.5005
R8209 VSS.n6026 VSS.n6015 4.57426
R8210 VSS.n6022 VSS.n6023 0.147342
R8211 VSS.n6023 VSS.n6024 0.147342
R8212 VSS.n6024 VSS.n6025 0.147342
R8213 VSS.n6027 VSS.n6026 2.37296
R8214 VSS.n6028 VSS.n6027 0.127318
R8215 VSS.n6029 VSS.n6028 0.127318
R8216 VSS.t0 VSS.n6029 2.73618
R8217 VSS.n6002 VSS.n6007 4.5005
R8218 VSS.n6004 VSS.n6008 4.5005
R8219 VSS.n6005 VSS.n6009 4.5005
R8220 VSS.n6006 VSS.n6010 4.57324
R8221 VSS.n6002 VSS.n6000 0.147342
R8222 VSS.n6003 VSS.n6004 0.0732424
R8223 VSS.n6004 VSS.n6005 0.147342
R8224 VSS.n6007 VSS.n6011 0.0721009
R8225 VSS.n6012 VSS.n6008 4.5005
R8226 VSS.n6013 VSS.n6009 4.5005
R8227 VSS.n6014 VSS.n6010 4.5005
R8228 VSS.n6000 VSS.n6011 4.57442
R8229 VSS.n6007 VSS.n6008 0.147342
R8230 VSS.n6008 VSS.n6009 0.147342
R8231 VSS.n6009 VSS.n6010 0.147342
R8232 VSS.n6011 VSS.n6012 2.39784
R8233 VSS.n6012 VSS.n6013 0.147342
R8234 VSS.n6013 VSS.n6014 0.147342
R8235 VSS.n6014 VSS.t138 3.13212
R8236 VSS.n5987 VSS.n5992 4.5005
R8237 VSS.n5989 VSS.n5993 4.5005
R8238 VSS.n5990 VSS.n5994 4.5005
R8239 VSS.n5991 VSS.n5995 4.57324
R8240 VSS.n5987 VSS.n5985 0.147342
R8241 VSS.n5988 VSS.n5989 0.0732424
R8242 VSS.n5989 VSS.n5990 0.147342
R8243 VSS.n5992 VSS.n5996 0.0721009
R8244 VSS.n5997 VSS.n5993 4.5005
R8245 VSS.n5998 VSS.n5994 4.5005
R8246 VSS.n5999 VSS.n5995 4.5005
R8247 VSS.n5985 VSS.n5996 4.57442
R8248 VSS.n5992 VSS.n5993 0.147342
R8249 VSS.n5993 VSS.n5994 0.147342
R8250 VSS.n5994 VSS.n5995 0.147342
R8251 VSS.n5996 VSS.n5997 2.39784
R8252 VSS.n5997 VSS.n5998 0.147342
R8253 VSS.n5998 VSS.n5999 0.147342
R8254 VSS.n5999 VSS.t136 3.13212
R8255 VSS.n5972 VSS.n5977 4.5005
R8256 VSS.n5974 VSS.n5978 4.5005
R8257 VSS.n5975 VSS.n5979 4.5005
R8258 VSS.n5976 VSS.n5980 4.57324
R8259 VSS.n5972 VSS.n5970 0.147342
R8260 VSS.n5973 VSS.n5974 0.0732424
R8261 VSS.n5974 VSS.n5975 0.147342
R8262 VSS.n5977 VSS.n5981 0.0721009
R8263 VSS.n5982 VSS.n5978 4.5005
R8264 VSS.n5983 VSS.n5979 4.5005
R8265 VSS.n5984 VSS.n5980 4.5005
R8266 VSS.n5970 VSS.n5981 4.57442
R8267 VSS.n5977 VSS.n5978 0.147342
R8268 VSS.n5978 VSS.n5979 0.147342
R8269 VSS.n5979 VSS.n5980 0.147342
R8270 VSS.n5981 VSS.n5982 2.39784
R8271 VSS.n5982 VSS.n5983 0.147342
R8272 VSS.n5983 VSS.n5984 0.147342
R8273 VSS.n5984 VSS.t349 3.13212
R8274 VSS.n5957 VSS.n5962 4.5005
R8275 VSS.n5959 VSS.n5963 4.5005
R8276 VSS.n5960 VSS.n5964 4.5005
R8277 VSS.n5961 VSS.n5965 4.57324
R8278 VSS.n5957 VSS.n5955 0.147342
R8279 VSS.n5958 VSS.n5959 0.0732424
R8280 VSS.n5959 VSS.n5960 0.147342
R8281 VSS.n5962 VSS.n5966 0.0721009
R8282 VSS.n5967 VSS.n5963 4.5005
R8283 VSS.n5968 VSS.n5964 4.5005
R8284 VSS.n5969 VSS.n5965 4.5005
R8285 VSS.n5955 VSS.n5966 4.57442
R8286 VSS.n5962 VSS.n5963 0.147342
R8287 VSS.n5963 VSS.n5964 0.147342
R8288 VSS.n5964 VSS.n5965 0.147342
R8289 VSS.n5966 VSS.n5967 2.39784
R8290 VSS.n5967 VSS.n5968 0.147342
R8291 VSS.n5968 VSS.n5969 0.147342
R8292 VSS.n5969 VSS.t296 3.13212
R8293 VSS.n5947 VSS.n5942 4.5005
R8294 VSS.n5948 VSS.n5944 4.5005
R8295 VSS.n5949 VSS.n5945 4.5005
R8296 VSS.n5950 VSS.n5946 4.57324
R8297 VSS.n5940 VSS.n5942 0.147342
R8298 VSS.n5943 VSS.n5944 0.0732424
R8299 VSS.n5944 VSS.n5945 0.147342
R8300 VSS.n5951 VSS.n5947 0.0722544
R8301 VSS.n5952 VSS.n5948 4.5005
R8302 VSS.n5953 VSS.n5949 4.5005
R8303 VSS.n5954 VSS.n5950 4.5005
R8304 VSS.n5951 VSS.n5940 4.57426
R8305 VSS.n5947 VSS.n5948 0.147342
R8306 VSS.n5948 VSS.n5949 0.147342
R8307 VSS.n5949 VSS.n5950 0.147342
R8308 VSS.n5952 VSS.n5951 2.37296
R8309 VSS.n5953 VSS.n5952 0.127318
R8310 VSS.n5954 VSS.n5953 0.127318
R8311 VSS.t0 VSS.n5954 2.73618
R8312 VSS.n5927 VSS.n5932 4.5005
R8313 VSS.n5929 VSS.n5933 4.5005
R8314 VSS.n5930 VSS.n5934 4.5005
R8315 VSS.n5931 VSS.n5935 4.57324
R8316 VSS.n5927 VSS.n5925 0.147342
R8317 VSS.n5928 VSS.n5929 0.0732424
R8318 VSS.n5929 VSS.n5930 0.147342
R8319 VSS.n5932 VSS.n5936 0.0721009
R8320 VSS.n5937 VSS.n5933 4.5005
R8321 VSS.n5938 VSS.n5934 4.5005
R8322 VSS.n5939 VSS.n5935 4.5005
R8323 VSS.n5925 VSS.n5936 4.57442
R8324 VSS.n5932 VSS.n5933 0.147342
R8325 VSS.n5933 VSS.n5934 0.147342
R8326 VSS.n5934 VSS.n5935 0.147342
R8327 VSS.n5936 VSS.n5937 2.39784
R8328 VSS.n5937 VSS.n5938 0.147342
R8329 VSS.n5938 VSS.n5939 0.147342
R8330 VSS.n5939 VSS.t545 3.13212
R8331 VSS.n5912 VSS.n5917 4.5005
R8332 VSS.n5914 VSS.n5918 4.5005
R8333 VSS.n5915 VSS.n5919 4.5005
R8334 VSS.n5916 VSS.n5920 4.57324
R8335 VSS.n5912 VSS.n5910 0.147342
R8336 VSS.n5913 VSS.n5914 0.0732424
R8337 VSS.n5914 VSS.n5915 0.147342
R8338 VSS.n5917 VSS.n5921 0.0721009
R8339 VSS.n5922 VSS.n5918 4.5005
R8340 VSS.n5923 VSS.n5919 4.5005
R8341 VSS.n5924 VSS.n5920 4.5005
R8342 VSS.n5910 VSS.n5921 4.57442
R8343 VSS.n5917 VSS.n5918 0.147342
R8344 VSS.n5918 VSS.n5919 0.147342
R8345 VSS.n5919 VSS.n5920 0.147342
R8346 VSS.n5921 VSS.n5922 2.39784
R8347 VSS.n5922 VSS.n5923 0.147342
R8348 VSS.n5923 VSS.n5924 0.147342
R8349 VSS.n5924 VSS.t282 3.13212
R8350 VSS.n5897 VSS.n5902 4.5005
R8351 VSS.n5899 VSS.n5903 4.5005
R8352 VSS.n5900 VSS.n5904 4.5005
R8353 VSS.n5901 VSS.n5905 4.57324
R8354 VSS.n5897 VSS.n5895 0.147342
R8355 VSS.n5898 VSS.n5899 0.0732424
R8356 VSS.n5899 VSS.n5900 0.147342
R8357 VSS.n5902 VSS.n5906 0.0721009
R8358 VSS.n5907 VSS.n5903 4.5005
R8359 VSS.n5908 VSS.n5904 4.5005
R8360 VSS.n5909 VSS.n5905 4.5005
R8361 VSS.n5895 VSS.n5906 4.57442
R8362 VSS.n5902 VSS.n5903 0.147342
R8363 VSS.n5903 VSS.n5904 0.147342
R8364 VSS.n5904 VSS.n5905 0.147342
R8365 VSS.n5906 VSS.n5907 2.39784
R8366 VSS.n5907 VSS.n5908 0.147342
R8367 VSS.n5908 VSS.n5909 0.147342
R8368 VSS.n5909 VSS.t600 3.13212
R8369 VSS.n5887 VSS.n5882 4.5005
R8370 VSS.n5888 VSS.n5884 4.5005
R8371 VSS.n5889 VSS.n5885 4.5005
R8372 VSS.n5890 VSS.n5886 4.57324
R8373 VSS.n5880 VSS.n5882 0.147342
R8374 VSS.n5883 VSS.n5884 0.0732424
R8375 VSS.n5884 VSS.n5885 0.147342
R8376 VSS.n5891 VSS.n5887 0.0722544
R8377 VSS.n5892 VSS.n5888 4.5005
R8378 VSS.n5893 VSS.n5889 4.5005
R8379 VSS.n5894 VSS.n5890 4.5005
R8380 VSS.n5891 VSS.n5880 4.57426
R8381 VSS.n5887 VSS.n5888 0.147342
R8382 VSS.n5888 VSS.n5889 0.147342
R8383 VSS.n5889 VSS.n5890 0.147342
R8384 VSS.n5892 VSS.n5891 2.37296
R8385 VSS.n5893 VSS.n5892 0.127318
R8386 VSS.n5894 VSS.n5893 0.127318
R8387 VSS.t0 VSS.n5894 2.73618
R8388 VSS.n5867 VSS.n5872 4.5005
R8389 VSS.n5869 VSS.n5873 4.5005
R8390 VSS.n5870 VSS.n5874 4.5005
R8391 VSS.n5871 VSS.n5875 4.57324
R8392 VSS.n5867 VSS.n5865 0.147342
R8393 VSS.n5868 VSS.n5869 0.0732424
R8394 VSS.n5869 VSS.n5870 0.147342
R8395 VSS.n5872 VSS.n5876 0.0721009
R8396 VSS.n5877 VSS.n5873 4.5005
R8397 VSS.n5878 VSS.n5874 4.5005
R8398 VSS.n5879 VSS.n5875 4.5005
R8399 VSS.n5865 VSS.n5876 4.57442
R8400 VSS.n5872 VSS.n5873 0.147342
R8401 VSS.n5873 VSS.n5874 0.147342
R8402 VSS.n5874 VSS.n5875 0.147342
R8403 VSS.n5876 VSS.n5877 2.39784
R8404 VSS.n5877 VSS.n5878 0.147342
R8405 VSS.n5878 VSS.n5879 0.147342
R8406 VSS.n5879 VSS.t2 3.13212
R8407 VSS.n5852 VSS.n5857 4.5005
R8408 VSS.n5854 VSS.n5858 4.5005
R8409 VSS.n5855 VSS.n5859 4.5005
R8410 VSS.n5856 VSS.n5860 4.57324
R8411 VSS.n5852 VSS.n5850 0.147342
R8412 VSS.n5853 VSS.n5854 0.0732424
R8413 VSS.n5854 VSS.n5855 0.147342
R8414 VSS.n5857 VSS.n5861 0.0721009
R8415 VSS.n5862 VSS.n5858 4.5005
R8416 VSS.n5863 VSS.n5859 4.5005
R8417 VSS.n5864 VSS.n5860 4.5005
R8418 VSS.n5850 VSS.n5861 4.57442
R8419 VSS.n5857 VSS.n5858 0.147342
R8420 VSS.n5858 VSS.n5859 0.147342
R8421 VSS.n5859 VSS.n5860 0.147342
R8422 VSS.n5861 VSS.n5862 2.39784
R8423 VSS.n5862 VSS.n5863 0.147342
R8424 VSS.n5863 VSS.n5864 0.147342
R8425 VSS.n5864 VSS.t153 3.13212
R8426 VSS.n5837 VSS.n5842 4.5005
R8427 VSS.n5839 VSS.n5843 4.5005
R8428 VSS.n5840 VSS.n5844 4.5005
R8429 VSS.n5841 VSS.n5845 4.57324
R8430 VSS.n5837 VSS.n5835 0.147342
R8431 VSS.n5838 VSS.n5839 0.0732424
R8432 VSS.n5839 VSS.n5840 0.147342
R8433 VSS.n5842 VSS.n5846 0.0721009
R8434 VSS.n5847 VSS.n5843 4.5005
R8435 VSS.n5848 VSS.n5844 4.5005
R8436 VSS.n5849 VSS.n5845 4.5005
R8437 VSS.n5835 VSS.n5846 4.57442
R8438 VSS.n5842 VSS.n5843 0.147342
R8439 VSS.n5843 VSS.n5844 0.147342
R8440 VSS.n5844 VSS.n5845 0.147342
R8441 VSS.n5846 VSS.n5847 2.39784
R8442 VSS.n5847 VSS.n5848 0.147342
R8443 VSS.n5848 VSS.n5849 0.147342
R8444 VSS.n5849 VSS.t264 3.13212
R8445 VSS.n5822 VSS.n5827 4.5005
R8446 VSS.n5824 VSS.n5828 4.5005
R8447 VSS.n5825 VSS.n5829 4.5005
R8448 VSS.n5826 VSS.n5830 4.57324
R8449 VSS.n5822 VSS.n5820 0.147342
R8450 VSS.n5823 VSS.n5824 0.0732424
R8451 VSS.n5824 VSS.n5825 0.147342
R8452 VSS.n5827 VSS.n5831 0.0721009
R8453 VSS.n5832 VSS.n5828 4.5005
R8454 VSS.n5833 VSS.n5829 4.5005
R8455 VSS.n5834 VSS.n5830 4.5005
R8456 VSS.n5820 VSS.n5831 4.57442
R8457 VSS.n5827 VSS.n5828 0.147342
R8458 VSS.n5828 VSS.n5829 0.147342
R8459 VSS.n5829 VSS.n5830 0.147342
R8460 VSS.n5831 VSS.n5832 2.39784
R8461 VSS.n5832 VSS.n5833 0.147342
R8462 VSS.n5833 VSS.n5834 0.147342
R8463 VSS.n5834 VSS.t97 3.13212
R8464 VSS.n5807 VSS.n5812 4.5005
R8465 VSS.n5809 VSS.n5813 4.5005
R8466 VSS.n5810 VSS.n5814 4.5005
R8467 VSS.n5811 VSS.n5815 4.57324
R8468 VSS.n5807 VSS.n5805 0.147342
R8469 VSS.n5808 VSS.n5809 0.0732424
R8470 VSS.n5809 VSS.n5810 0.147342
R8471 VSS.n5812 VSS.n5816 0.0721009
R8472 VSS.n5817 VSS.n5813 4.5005
R8473 VSS.n5818 VSS.n5814 4.5005
R8474 VSS.n5819 VSS.n5815 4.5005
R8475 VSS.n5805 VSS.n5816 4.57442
R8476 VSS.n5812 VSS.n5813 0.147342
R8477 VSS.n5813 VSS.n5814 0.147342
R8478 VSS.n5814 VSS.n5815 0.147342
R8479 VSS.n5816 VSS.n5817 2.39784
R8480 VSS.n5817 VSS.n5818 0.147342
R8481 VSS.n5818 VSS.n5819 0.147342
R8482 VSS.n5819 VSS.t471 3.13212
R8483 VSS.n5792 VSS.n5797 4.5005
R8484 VSS.n5794 VSS.n5798 4.5005
R8485 VSS.n5795 VSS.n5799 4.5005
R8486 VSS.n5796 VSS.n5800 4.57324
R8487 VSS.n5792 VSS.n5790 0.147342
R8488 VSS.n5793 VSS.n5794 0.0732424
R8489 VSS.n5794 VSS.n5795 0.147342
R8490 VSS.n5797 VSS.n5801 0.0721009
R8491 VSS.n5802 VSS.n5798 4.5005
R8492 VSS.n5803 VSS.n5799 4.5005
R8493 VSS.n5804 VSS.n5800 4.5005
R8494 VSS.n5790 VSS.n5801 4.57442
R8495 VSS.n5797 VSS.n5798 0.147342
R8496 VSS.n5798 VSS.n5799 0.147342
R8497 VSS.n5799 VSS.n5800 0.147342
R8498 VSS.n5801 VSS.n5802 2.39784
R8499 VSS.n5802 VSS.n5803 0.147342
R8500 VSS.n5803 VSS.n5804 0.147342
R8501 VSS.n5804 VSS.t60 3.13212
R8502 VSS.n5782 VSS.n5777 4.5005
R8503 VSS.n5783 VSS.n5779 4.5005
R8504 VSS.n5784 VSS.n5780 4.5005
R8505 VSS.n5785 VSS.n5781 4.57324
R8506 VSS.n5775 VSS.n5777 0.147342
R8507 VSS.n5778 VSS.n5779 0.0732424
R8508 VSS.n5779 VSS.n5780 0.147342
R8509 VSS.n5786 VSS.n5782 0.0722544
R8510 VSS.n5787 VSS.n5783 4.5005
R8511 VSS.n5788 VSS.n5784 4.5005
R8512 VSS.n5789 VSS.n5785 4.5005
R8513 VSS.n5786 VSS.n5775 4.57426
R8514 VSS.n5782 VSS.n5783 0.147342
R8515 VSS.n5783 VSS.n5784 0.147342
R8516 VSS.n5784 VSS.n5785 0.147342
R8517 VSS.n5787 VSS.n5786 2.37296
R8518 VSS.n5788 VSS.n5787 0.127318
R8519 VSS.n5789 VSS.n5788 0.127318
R8520 VSS.t0 VSS.n5789 2.73618
R8521 VSS.n5762 VSS.n5767 4.5005
R8522 VSS.n5764 VSS.n5768 4.5005
R8523 VSS.n5765 VSS.n5769 4.5005
R8524 VSS.n5766 VSS.n5770 4.57324
R8525 VSS.n5762 VSS.n5760 0.147342
R8526 VSS.n5763 VSS.n5764 0.0732424
R8527 VSS.n5764 VSS.n5765 0.147342
R8528 VSS.n5767 VSS.n5771 0.0721009
R8529 VSS.n5772 VSS.n5768 4.5005
R8530 VSS.n5773 VSS.n5769 4.5005
R8531 VSS.n5774 VSS.n5770 4.5005
R8532 VSS.n5760 VSS.n5771 4.57442
R8533 VSS.n5767 VSS.n5768 0.147342
R8534 VSS.n5768 VSS.n5769 0.147342
R8535 VSS.n5769 VSS.n5770 0.147342
R8536 VSS.n5771 VSS.n5772 2.39784
R8537 VSS.n5772 VSS.n5773 0.147342
R8538 VSS.n5773 VSS.n5774 0.147342
R8539 VSS.n5774 VSS.t214 3.13212
R8540 VSS.n5747 VSS.n5752 4.5005
R8541 VSS.n5749 VSS.n5753 4.5005
R8542 VSS.n5750 VSS.n5754 4.5005
R8543 VSS.n5751 VSS.n5755 4.57324
R8544 VSS.n5747 VSS.n5745 0.147342
R8545 VSS.n5748 VSS.n5749 0.0732424
R8546 VSS.n5749 VSS.n5750 0.147342
R8547 VSS.n5752 VSS.n5756 0.0721009
R8548 VSS.n5757 VSS.n5753 4.5005
R8549 VSS.n5758 VSS.n5754 4.5005
R8550 VSS.n5759 VSS.n5755 4.5005
R8551 VSS.n5745 VSS.n5756 4.57442
R8552 VSS.n5752 VSS.n5753 0.147342
R8553 VSS.n5753 VSS.n5754 0.147342
R8554 VSS.n5754 VSS.n5755 0.147342
R8555 VSS.n5756 VSS.n5757 2.39784
R8556 VSS.n5757 VSS.n5758 0.147342
R8557 VSS.n5758 VSS.n5759 0.147342
R8558 VSS.n5759 VSS.t208 3.13212
R8559 VSS.n5732 VSS.n5737 4.5005
R8560 VSS.n5734 VSS.n5738 4.5005
R8561 VSS.n5735 VSS.n5739 4.5005
R8562 VSS.n5736 VSS.n5740 4.57324
R8563 VSS.n5732 VSS.n5730 0.147342
R8564 VSS.n5733 VSS.n5734 0.0732424
R8565 VSS.n5734 VSS.n5735 0.147342
R8566 VSS.n5737 VSS.n5741 0.0721009
R8567 VSS.n5742 VSS.n5738 4.5005
R8568 VSS.n5743 VSS.n5739 4.5005
R8569 VSS.n5744 VSS.n5740 4.5005
R8570 VSS.n5730 VSS.n5741 4.57442
R8571 VSS.n5737 VSS.n5738 0.147342
R8572 VSS.n5738 VSS.n5739 0.147342
R8573 VSS.n5739 VSS.n5740 0.147342
R8574 VSS.n5741 VSS.n5742 2.39784
R8575 VSS.n5742 VSS.n5743 0.147342
R8576 VSS.n5743 VSS.n5744 0.147342
R8577 VSS.n5744 VSS.t129 3.13212
R8578 VSS.n5722 VSS.n5717 4.5005
R8579 VSS.n5723 VSS.n5719 4.5005
R8580 VSS.n5724 VSS.n5720 4.5005
R8581 VSS.n5725 VSS.n5721 4.57324
R8582 VSS.n5715 VSS.n5717 0.147342
R8583 VSS.n5718 VSS.n5719 0.0732424
R8584 VSS.n5719 VSS.n5720 0.147342
R8585 VSS.n5726 VSS.n5722 0.0722544
R8586 VSS.n5727 VSS.n5723 4.5005
R8587 VSS.n5728 VSS.n5724 4.5005
R8588 VSS.n5729 VSS.n5725 4.5005
R8589 VSS.n5726 VSS.n5715 4.57426
R8590 VSS.n5722 VSS.n5723 0.147342
R8591 VSS.n5723 VSS.n5724 0.147342
R8592 VSS.n5724 VSS.n5725 0.147342
R8593 VSS.n5727 VSS.n5726 2.37296
R8594 VSS.n5728 VSS.n5727 0.127318
R8595 VSS.n5729 VSS.n5728 0.127318
R8596 VSS.t0 VSS.n5729 2.73618
R8597 VSS.n5702 VSS.n5707 4.5005
R8598 VSS.n5704 VSS.n5708 4.5005
R8599 VSS.n5705 VSS.n5709 4.5005
R8600 VSS.n5706 VSS.n5710 4.57324
R8601 VSS.n5702 VSS.n5700 0.147342
R8602 VSS.n5703 VSS.n5704 0.0732424
R8603 VSS.n5704 VSS.n5705 0.147342
R8604 VSS.n5707 VSS.n5711 0.0721009
R8605 VSS.n5712 VSS.n5708 4.5005
R8606 VSS.n5713 VSS.n5709 4.5005
R8607 VSS.n5714 VSS.n5710 4.5005
R8608 VSS.n5700 VSS.n5711 4.57442
R8609 VSS.n5707 VSS.n5708 0.147342
R8610 VSS.n5708 VSS.n5709 0.147342
R8611 VSS.n5709 VSS.n5710 0.147342
R8612 VSS.n5711 VSS.n5712 2.39784
R8613 VSS.n5712 VSS.n5713 0.147342
R8614 VSS.n5713 VSS.n5714 0.147342
R8615 VSS.n5714 VSS.t38 3.13212
R8616 VSS.n5687 VSS.n5692 4.5005
R8617 VSS.n5689 VSS.n5693 4.5005
R8618 VSS.n5690 VSS.n5694 4.5005
R8619 VSS.n5691 VSS.n5695 4.57324
R8620 VSS.n5687 VSS.n5685 0.147342
R8621 VSS.n5688 VSS.n5689 0.0732424
R8622 VSS.n5689 VSS.n5690 0.147342
R8623 VSS.n5692 VSS.n5696 0.0721009
R8624 VSS.n5697 VSS.n5693 4.5005
R8625 VSS.n5698 VSS.n5694 4.5005
R8626 VSS.n5699 VSS.n5695 4.5005
R8627 VSS.n5685 VSS.n5696 4.57442
R8628 VSS.n5692 VSS.n5693 0.147342
R8629 VSS.n5693 VSS.n5694 0.147342
R8630 VSS.n5694 VSS.n5695 0.147342
R8631 VSS.n5696 VSS.n5697 2.39784
R8632 VSS.n5697 VSS.n5698 0.147342
R8633 VSS.n5698 VSS.n5699 0.147342
R8634 VSS.n5699 VSS.t99 3.13212
R8635 VSS.n5672 VSS.n5677 4.5005
R8636 VSS.n5674 VSS.n5678 4.5005
R8637 VSS.n5675 VSS.n5679 4.5005
R8638 VSS.n5676 VSS.n5680 4.57324
R8639 VSS.n5672 VSS.n5670 0.147342
R8640 VSS.n5673 VSS.n5674 0.0732424
R8641 VSS.n5674 VSS.n5675 0.147342
R8642 VSS.n5677 VSS.n5681 0.0721009
R8643 VSS.n5682 VSS.n5678 4.5005
R8644 VSS.n5683 VSS.n5679 4.5005
R8645 VSS.n5684 VSS.n5680 4.5005
R8646 VSS.n5670 VSS.n5681 4.57442
R8647 VSS.n5677 VSS.n5678 0.147342
R8648 VSS.n5678 VSS.n5679 0.147342
R8649 VSS.n5679 VSS.n5680 0.147342
R8650 VSS.n5681 VSS.n5682 2.39784
R8651 VSS.n5682 VSS.n5683 0.147342
R8652 VSS.n5683 VSS.n5684 0.147342
R8653 VSS.n5684 VSS.t300 3.13212
R8654 VSS.n5657 VSS.n5662 4.5005
R8655 VSS.n5659 VSS.n5663 4.5005
R8656 VSS.n5660 VSS.n5664 4.5005
R8657 VSS.n5661 VSS.n5665 4.57324
R8658 VSS.n5657 VSS.n5655 0.147342
R8659 VSS.n5658 VSS.n5659 0.0732424
R8660 VSS.n5659 VSS.n5660 0.147342
R8661 VSS.n5662 VSS.n5666 0.0721009
R8662 VSS.n5667 VSS.n5663 4.5005
R8663 VSS.n5668 VSS.n5664 4.5005
R8664 VSS.n5669 VSS.n5665 4.5005
R8665 VSS.n5655 VSS.n5666 4.57442
R8666 VSS.n5662 VSS.n5663 0.147342
R8667 VSS.n5663 VSS.n5664 0.147342
R8668 VSS.n5664 VSS.n5665 0.147342
R8669 VSS.n5666 VSS.n5667 2.39784
R8670 VSS.n5667 VSS.n5668 0.147342
R8671 VSS.n5668 VSS.n5669 0.147342
R8672 VSS.n5669 VSS.t308 3.13212
R8673 VSS.n5647 VSS.n5642 4.5005
R8674 VSS.n5648 VSS.n5644 4.5005
R8675 VSS.n5649 VSS.n5645 4.5005
R8676 VSS.n5650 VSS.n5646 4.57324
R8677 VSS.n5640 VSS.n5642 0.147342
R8678 VSS.n5643 VSS.n5644 0.0732424
R8679 VSS.n5644 VSS.n5645 0.147342
R8680 VSS.n5651 VSS.n5647 0.0722544
R8681 VSS.n5652 VSS.n5648 4.5005
R8682 VSS.n5653 VSS.n5649 4.5005
R8683 VSS.n5654 VSS.n5650 4.5005
R8684 VSS.n5651 VSS.n5640 4.57426
R8685 VSS.n5647 VSS.n5648 0.147342
R8686 VSS.n5648 VSS.n5649 0.147342
R8687 VSS.n5649 VSS.n5650 0.147342
R8688 VSS.n5652 VSS.n5651 2.37296
R8689 VSS.n5653 VSS.n5652 0.127318
R8690 VSS.n5654 VSS.n5653 0.127318
R8691 VSS.t0 VSS.n5654 2.73618
R8692 VSS.n5627 VSS.n5632 4.5005
R8693 VSS.n5629 VSS.n5633 4.5005
R8694 VSS.n5630 VSS.n5634 4.5005
R8695 VSS.n5631 VSS.n5635 4.57324
R8696 VSS.n5627 VSS.n5625 0.147342
R8697 VSS.n5628 VSS.n5629 0.0732424
R8698 VSS.n5629 VSS.n5630 0.147342
R8699 VSS.n5632 VSS.n5636 0.0721009
R8700 VSS.n5637 VSS.n5633 4.5005
R8701 VSS.n5638 VSS.n5634 4.5005
R8702 VSS.n5639 VSS.n5635 4.5005
R8703 VSS.n5625 VSS.n5636 4.57442
R8704 VSS.n5632 VSS.n5633 0.147342
R8705 VSS.n5633 VSS.n5634 0.147342
R8706 VSS.n5634 VSS.n5635 0.147342
R8707 VSS.n5636 VSS.n5637 2.39784
R8708 VSS.n5637 VSS.n5638 0.147342
R8709 VSS.n5638 VSS.n5639 0.147342
R8710 VSS.n5639 VSS.t543 3.13212
R8711 VSS.n5612 VSS.n5617 4.5005
R8712 VSS.n5614 VSS.n5618 4.5005
R8713 VSS.n5615 VSS.n5619 4.5005
R8714 VSS.n5616 VSS.n5620 4.57324
R8715 VSS.n5612 VSS.n5610 0.147342
R8716 VSS.n5613 VSS.n5614 0.0732424
R8717 VSS.n5614 VSS.n5615 0.147342
R8718 VSS.n5617 VSS.n5621 0.0721009
R8719 VSS.n5622 VSS.n5618 4.5005
R8720 VSS.n5623 VSS.n5619 4.5005
R8721 VSS.n5624 VSS.n5620 4.5005
R8722 VSS.n5610 VSS.n5621 4.57442
R8723 VSS.n5617 VSS.n5618 0.147342
R8724 VSS.n5618 VSS.n5619 0.147342
R8725 VSS.n5619 VSS.n5620 0.147342
R8726 VSS.n5621 VSS.n5622 2.39784
R8727 VSS.n5622 VSS.n5623 0.147342
R8728 VSS.n5623 VSS.n5624 0.147342
R8729 VSS.n5624 VSS.t280 3.13212
R8730 VSS.n5597 VSS.n5602 4.5005
R8731 VSS.n5599 VSS.n5603 4.5005
R8732 VSS.n5600 VSS.n5604 4.5005
R8733 VSS.n5601 VSS.n5605 4.57324
R8734 VSS.n5597 VSS.n5595 0.147342
R8735 VSS.n5598 VSS.n5599 0.0732424
R8736 VSS.n5599 VSS.n5600 0.147342
R8737 VSS.n5602 VSS.n5606 0.0721009
R8738 VSS.n5607 VSS.n5603 4.5005
R8739 VSS.n5608 VSS.n5604 4.5005
R8740 VSS.n5609 VSS.n5605 4.5005
R8741 VSS.n5595 VSS.n5606 4.57442
R8742 VSS.n5602 VSS.n5603 0.147342
R8743 VSS.n5603 VSS.n5604 0.147342
R8744 VSS.n5604 VSS.n5605 0.147342
R8745 VSS.n5606 VSS.n5607 2.39784
R8746 VSS.n5607 VSS.n5608 0.147342
R8747 VSS.n5608 VSS.n5609 0.147342
R8748 VSS.n5609 VSS.t164 3.13212
R8749 VSS.n5587 VSS.n5582 4.5005
R8750 VSS.n5588 VSS.n5584 4.5005
R8751 VSS.n5589 VSS.n5585 4.5005
R8752 VSS.n5590 VSS.n5586 4.57324
R8753 VSS.n5580 VSS.n5582 0.147342
R8754 VSS.n5583 VSS.n5584 0.0732424
R8755 VSS.n5584 VSS.n5585 0.147342
R8756 VSS.n5591 VSS.n5587 0.0722544
R8757 VSS.n5592 VSS.n5588 4.5005
R8758 VSS.n5593 VSS.n5589 4.5005
R8759 VSS.n5594 VSS.n5590 4.5005
R8760 VSS.n5591 VSS.n5580 4.57426
R8761 VSS.n5587 VSS.n5588 0.147342
R8762 VSS.n5588 VSS.n5589 0.147342
R8763 VSS.n5589 VSS.n5590 0.147342
R8764 VSS.n5592 VSS.n5591 2.37296
R8765 VSS.n5593 VSS.n5592 0.127318
R8766 VSS.n5594 VSS.n5593 0.127318
R8767 VSS.t0 VSS.n5594 2.73618
R8768 VSS.n5567 VSS.n5572 4.5005
R8769 VSS.n5569 VSS.n5573 4.5005
R8770 VSS.n5570 VSS.n5574 4.5005
R8771 VSS.n5571 VSS.n5575 4.57324
R8772 VSS.n5567 VSS.n5565 0.147342
R8773 VSS.n5568 VSS.n5569 0.0732424
R8774 VSS.n5569 VSS.n5570 0.147342
R8775 VSS.n5572 VSS.n5576 0.0721009
R8776 VSS.n5577 VSS.n5573 4.5005
R8777 VSS.n5578 VSS.n5574 4.5005
R8778 VSS.n5579 VSS.n5575 4.5005
R8779 VSS.n5565 VSS.n5576 4.57442
R8780 VSS.n5572 VSS.n5573 0.147342
R8781 VSS.n5573 VSS.n5574 0.147342
R8782 VSS.n5574 VSS.n5575 0.147342
R8783 VSS.n5576 VSS.n5577 2.39784
R8784 VSS.n5577 VSS.n5578 0.147342
R8785 VSS.n5578 VSS.n5579 0.147342
R8786 VSS.n5579 VSS.t440 3.13212
R8787 VSS.n5552 VSS.n5557 4.5005
R8788 VSS.n5554 VSS.n5558 4.5005
R8789 VSS.n5555 VSS.n5559 4.5005
R8790 VSS.n5556 VSS.n5560 4.57324
R8791 VSS.n5552 VSS.n5550 0.147342
R8792 VSS.n5553 VSS.n5554 0.0732424
R8793 VSS.n5554 VSS.n5555 0.147342
R8794 VSS.n5557 VSS.n5561 0.0721009
R8795 VSS.n5562 VSS.n5558 4.5005
R8796 VSS.n5563 VSS.n5559 4.5005
R8797 VSS.n5564 VSS.n5560 4.5005
R8798 VSS.n5550 VSS.n5561 4.57442
R8799 VSS.n5557 VSS.n5558 0.147342
R8800 VSS.n5558 VSS.n5559 0.147342
R8801 VSS.n5559 VSS.n5560 0.147342
R8802 VSS.n5561 VSS.n5562 2.39784
R8803 VSS.n5562 VSS.n5563 0.147342
R8804 VSS.n5563 VSS.n5564 0.147342
R8805 VSS.n5564 VSS.t155 3.13212
R8806 VSS.n5537 VSS.n5542 4.5005
R8807 VSS.n5539 VSS.n5543 4.5005
R8808 VSS.n5540 VSS.n5544 4.5005
R8809 VSS.n5541 VSS.n5545 4.57324
R8810 VSS.n5537 VSS.n5535 0.147342
R8811 VSS.n5538 VSS.n5539 0.0732424
R8812 VSS.n5539 VSS.n5540 0.147342
R8813 VSS.n5542 VSS.n5546 0.0721009
R8814 VSS.n5547 VSS.n5543 4.5005
R8815 VSS.n5548 VSS.n5544 4.5005
R8816 VSS.n5549 VSS.n5545 4.5005
R8817 VSS.n5535 VSS.n5546 4.57442
R8818 VSS.n5542 VSS.n5543 0.147342
R8819 VSS.n5543 VSS.n5544 0.147342
R8820 VSS.n5544 VSS.n5545 0.147342
R8821 VSS.n5546 VSS.n5547 2.39784
R8822 VSS.n5547 VSS.n5548 0.147342
R8823 VSS.n5548 VSS.n5549 0.147342
R8824 VSS.n5549 VSS.t262 3.13212
R8825 VSS.n5522 VSS.n5527 4.5005
R8826 VSS.n5524 VSS.n5528 4.5005
R8827 VSS.n5525 VSS.n5529 4.5005
R8828 VSS.n5526 VSS.n5530 4.57324
R8829 VSS.n5522 VSS.n5520 0.147342
R8830 VSS.n5523 VSS.n5524 0.0732424
R8831 VSS.n5524 VSS.n5525 0.147342
R8832 VSS.n5527 VSS.n5531 0.0721009
R8833 VSS.n5532 VSS.n5528 4.5005
R8834 VSS.n5533 VSS.n5529 4.5005
R8835 VSS.n5534 VSS.n5530 4.5005
R8836 VSS.n5520 VSS.n5531 4.57442
R8837 VSS.n5527 VSS.n5528 0.147342
R8838 VSS.n5528 VSS.n5529 0.147342
R8839 VSS.n5529 VSS.n5530 0.147342
R8840 VSS.n5531 VSS.n5532 2.39784
R8841 VSS.n5532 VSS.n5533 0.147342
R8842 VSS.n5533 VSS.n5534 0.147342
R8843 VSS.n5534 VSS.t267 3.13212
R8844 VSS.n5507 VSS.n5512 4.5005
R8845 VSS.n5509 VSS.n5513 4.5005
R8846 VSS.n5510 VSS.n5514 4.5005
R8847 VSS.n5511 VSS.n5515 4.57324
R8848 VSS.n5507 VSS.n5505 0.147342
R8849 VSS.n5508 VSS.n5509 0.0732424
R8850 VSS.n5509 VSS.n5510 0.147342
R8851 VSS.n5512 VSS.n5516 0.0721009
R8852 VSS.n5517 VSS.n5513 4.5005
R8853 VSS.n5518 VSS.n5514 4.5005
R8854 VSS.n5519 VSS.n5515 4.5005
R8855 VSS.n5505 VSS.n5516 4.57442
R8856 VSS.n5512 VSS.n5513 0.147342
R8857 VSS.n5513 VSS.n5514 0.147342
R8858 VSS.n5514 VSS.n5515 0.147342
R8859 VSS.n5516 VSS.n5517 2.39784
R8860 VSS.n5517 VSS.n5518 0.147342
R8861 VSS.n5518 VSS.n5519 0.147342
R8862 VSS.n5519 VSS.t479 3.13212
R8863 VSS.n5492 VSS.n5497 4.5005
R8864 VSS.n5494 VSS.n5498 4.5005
R8865 VSS.n5495 VSS.n5499 4.5005
R8866 VSS.n5496 VSS.n5500 4.57324
R8867 VSS.n5492 VSS.n5490 0.147342
R8868 VSS.n5493 VSS.n5494 0.0732424
R8869 VSS.n5494 VSS.n5495 0.147342
R8870 VSS.n5497 VSS.n5501 0.0721009
R8871 VSS.n5502 VSS.n5498 4.5005
R8872 VSS.n5503 VSS.n5499 4.5005
R8873 VSS.n5504 VSS.n5500 4.5005
R8874 VSS.n5490 VSS.n5501 4.57442
R8875 VSS.n5497 VSS.n5498 0.147342
R8876 VSS.n5498 VSS.n5499 0.147342
R8877 VSS.n5499 VSS.n5500 0.147342
R8878 VSS.n5501 VSS.n5502 2.39784
R8879 VSS.n5502 VSS.n5503 0.147342
R8880 VSS.n5503 VSS.n5504 0.147342
R8881 VSS.n5504 VSS.t59 3.13212
R8882 VSS.n5482 VSS.n5477 4.5005
R8883 VSS.n5483 VSS.n5479 4.5005
R8884 VSS.n5484 VSS.n5480 4.5005
R8885 VSS.n5485 VSS.n5481 4.57324
R8886 VSS.n5475 VSS.n5477 0.147342
R8887 VSS.n5478 VSS.n5479 0.0732424
R8888 VSS.n5479 VSS.n5480 0.147342
R8889 VSS.n5486 VSS.n5482 0.0722544
R8890 VSS.n5487 VSS.n5483 4.5005
R8891 VSS.n5488 VSS.n5484 4.5005
R8892 VSS.n5489 VSS.n5485 4.5005
R8893 VSS.n5486 VSS.n5475 4.57426
R8894 VSS.n5482 VSS.n5483 0.147342
R8895 VSS.n5483 VSS.n5484 0.147342
R8896 VSS.n5484 VSS.n5485 0.147342
R8897 VSS.n5487 VSS.n5486 2.37296
R8898 VSS.n5488 VSS.n5487 0.127318
R8899 VSS.n5489 VSS.n5488 0.127318
R8900 VSS.t0 VSS.n5489 2.73618
R8901 VSS.n5462 VSS.n5467 4.5005
R8902 VSS.n5464 VSS.n5468 4.5005
R8903 VSS.n5465 VSS.n5469 4.5005
R8904 VSS.n5466 VSS.n5470 4.57324
R8905 VSS.n5462 VSS.n5460 0.147342
R8906 VSS.n5463 VSS.n5464 0.0732424
R8907 VSS.n5464 VSS.n5465 0.147342
R8908 VSS.n5467 VSS.n5471 0.0721009
R8909 VSS.n5472 VSS.n5468 4.5005
R8910 VSS.n5473 VSS.n5469 4.5005
R8911 VSS.n5474 VSS.n5470 4.5005
R8912 VSS.n5460 VSS.n5471 4.57442
R8913 VSS.n5467 VSS.n5468 0.147342
R8914 VSS.n5468 VSS.n5469 0.147342
R8915 VSS.n5469 VSS.n5470 0.147342
R8916 VSS.n5471 VSS.n5472 2.39784
R8917 VSS.n5472 VSS.n5473 0.147342
R8918 VSS.n5473 VSS.n5474 0.147342
R8919 VSS.n5474 VSS.t216 3.13212
R8920 VSS.n5447 VSS.n5452 4.5005
R8921 VSS.n5449 VSS.n5453 4.5005
R8922 VSS.n5450 VSS.n5454 4.5005
R8923 VSS.n5451 VSS.n5455 4.57324
R8924 VSS.n5447 VSS.n5445 0.147342
R8925 VSS.n5448 VSS.n5449 0.0732424
R8926 VSS.n5449 VSS.n5450 0.147342
R8927 VSS.n5452 VSS.n5456 0.0721009
R8928 VSS.n5457 VSS.n5453 4.5005
R8929 VSS.n5458 VSS.n5454 4.5005
R8930 VSS.n5459 VSS.n5455 4.5005
R8931 VSS.n5445 VSS.n5456 4.57442
R8932 VSS.n5452 VSS.n5453 0.147342
R8933 VSS.n5453 VSS.n5454 0.147342
R8934 VSS.n5454 VSS.n5455 0.147342
R8935 VSS.n5456 VSS.n5457 2.39784
R8936 VSS.n5457 VSS.n5458 0.147342
R8937 VSS.n5458 VSS.n5459 0.147342
R8938 VSS.n5459 VSS.t209 3.13212
R8939 VSS.n5432 VSS.n5437 4.5005
R8940 VSS.n5434 VSS.n5438 4.5005
R8941 VSS.n5435 VSS.n5439 4.5005
R8942 VSS.n5436 VSS.n5440 4.57324
R8943 VSS.n5432 VSS.n5430 0.147342
R8944 VSS.n5433 VSS.n5434 0.0732424
R8945 VSS.n5434 VSS.n5435 0.147342
R8946 VSS.n5437 VSS.n5441 0.0721009
R8947 VSS.n5442 VSS.n5438 4.5005
R8948 VSS.n5443 VSS.n5439 4.5005
R8949 VSS.n5444 VSS.n5440 4.5005
R8950 VSS.n5430 VSS.n5441 4.57442
R8951 VSS.n5437 VSS.n5438 0.147342
R8952 VSS.n5438 VSS.n5439 0.147342
R8953 VSS.n5439 VSS.n5440 0.147342
R8954 VSS.n5441 VSS.n5442 2.39784
R8955 VSS.n5442 VSS.n5443 0.147342
R8956 VSS.n5443 VSS.n5444 0.147342
R8957 VSS.n5444 VSS.t131 3.13212
R8958 VSS.n5422 VSS.n5417 4.5005
R8959 VSS.n5423 VSS.n5419 4.5005
R8960 VSS.n5424 VSS.n5420 4.5005
R8961 VSS.n5425 VSS.n5421 4.57324
R8962 VSS.n5415 VSS.n5417 0.147342
R8963 VSS.n5418 VSS.n5419 0.0732424
R8964 VSS.n5419 VSS.n5420 0.147342
R8965 VSS.n5426 VSS.n5422 0.0722544
R8966 VSS.n5427 VSS.n5423 4.5005
R8967 VSS.n5428 VSS.n5424 4.5005
R8968 VSS.n5429 VSS.n5425 4.5005
R8969 VSS.n5426 VSS.n5415 4.57426
R8970 VSS.n5422 VSS.n5423 0.147342
R8971 VSS.n5423 VSS.n5424 0.147342
R8972 VSS.n5424 VSS.n5425 0.147342
R8973 VSS.n5427 VSS.n5426 2.37296
R8974 VSS.n5428 VSS.n5427 0.127318
R8975 VSS.n5429 VSS.n5428 0.127318
R8976 VSS.t0 VSS.n5429 2.73618
R8977 VSS.n5402 VSS.n5407 4.5005
R8978 VSS.n5404 VSS.n5408 4.5005
R8979 VSS.n5405 VSS.n5409 4.5005
R8980 VSS.n5406 VSS.n5410 4.57324
R8981 VSS.n5402 VSS.n5400 0.147342
R8982 VSS.n5403 VSS.n5404 0.0732424
R8983 VSS.n5404 VSS.n5405 0.147342
R8984 VSS.n5407 VSS.n5411 0.0721009
R8985 VSS.n5412 VSS.n5408 4.5005
R8986 VSS.n5413 VSS.n5409 4.5005
R8987 VSS.n5414 VSS.n5410 4.5005
R8988 VSS.n5400 VSS.n5411 4.57442
R8989 VSS.n5407 VSS.n5408 0.147342
R8990 VSS.n5408 VSS.n5409 0.147342
R8991 VSS.n5409 VSS.n5410 0.147342
R8992 VSS.n5411 VSS.n5412 2.39784
R8993 VSS.n5412 VSS.n5413 0.147342
R8994 VSS.n5413 VSS.n5414 0.147342
R8995 VSS.n5414 VSS.t139 3.13212
R8996 VSS.n5387 VSS.n5392 4.5005
R8997 VSS.n5389 VSS.n5393 4.5005
R8998 VSS.n5390 VSS.n5394 4.5005
R8999 VSS.n5391 VSS.n5395 4.57324
R9000 VSS.n5387 VSS.n5385 0.147342
R9001 VSS.n5388 VSS.n5389 0.0732424
R9002 VSS.n5389 VSS.n5390 0.147342
R9003 VSS.n5392 VSS.n5396 0.0721009
R9004 VSS.n5397 VSS.n5393 4.5005
R9005 VSS.n5398 VSS.n5394 4.5005
R9006 VSS.n5399 VSS.n5395 4.5005
R9007 VSS.n5385 VSS.n5396 4.57442
R9008 VSS.n5392 VSS.n5393 0.147342
R9009 VSS.n5393 VSS.n5394 0.147342
R9010 VSS.n5394 VSS.n5395 0.147342
R9011 VSS.n5396 VSS.n5397 2.39784
R9012 VSS.n5397 VSS.n5398 0.147342
R9013 VSS.n5398 VSS.n5399 0.147342
R9014 VSS.n5399 VSS.t101 3.13212
R9015 VSS.n5372 VSS.n5377 4.5005
R9016 VSS.n5374 VSS.n5378 4.5005
R9017 VSS.n5375 VSS.n5379 4.5005
R9018 VSS.n5376 VSS.n5380 4.57324
R9019 VSS.n5372 VSS.n5370 0.147342
R9020 VSS.n5373 VSS.n5374 0.0732424
R9021 VSS.n5374 VSS.n5375 0.147342
R9022 VSS.n5377 VSS.n5381 0.0721009
R9023 VSS.n5382 VSS.n5378 4.5005
R9024 VSS.n5383 VSS.n5379 4.5005
R9025 VSS.n5384 VSS.n5380 4.5005
R9026 VSS.n5370 VSS.n5381 4.57442
R9027 VSS.n5377 VSS.n5378 0.147342
R9028 VSS.n5378 VSS.n5379 0.147342
R9029 VSS.n5379 VSS.n5380 0.147342
R9030 VSS.n5381 VSS.n5382 2.39784
R9031 VSS.n5382 VSS.n5383 0.147342
R9032 VSS.n5383 VSS.n5384 0.147342
R9033 VSS.n5384 VSS.t284 3.13212
R9034 VSS.n5357 VSS.n5362 4.5005
R9035 VSS.n5359 VSS.n5363 4.5005
R9036 VSS.n5360 VSS.n5364 4.5005
R9037 VSS.n5361 VSS.n5365 4.57324
R9038 VSS.n5357 VSS.n5355 0.147342
R9039 VSS.n5358 VSS.n5359 0.0732424
R9040 VSS.n5359 VSS.n5360 0.147342
R9041 VSS.n5362 VSS.n5366 0.0721009
R9042 VSS.n5367 VSS.n5363 4.5005
R9043 VSS.n5368 VSS.n5364 4.5005
R9044 VSS.n5369 VSS.n5365 4.5005
R9045 VSS.n5355 VSS.n5366 4.57442
R9046 VSS.n5362 VSS.n5363 0.147342
R9047 VSS.n5363 VSS.n5364 0.147342
R9048 VSS.n5364 VSS.n5365 0.147342
R9049 VSS.n5366 VSS.n5367 2.39784
R9050 VSS.n5367 VSS.n5368 0.147342
R9051 VSS.n5368 VSS.n5369 0.147342
R9052 VSS.n5369 VSS.t309 3.13212
R9053 VSS.n5347 VSS.n5342 4.5005
R9054 VSS.n5348 VSS.n5344 4.5005
R9055 VSS.n5349 VSS.n5345 4.5005
R9056 VSS.n5350 VSS.n5346 4.57324
R9057 VSS.n5340 VSS.n5342 0.147342
R9058 VSS.n5343 VSS.n5344 0.0732424
R9059 VSS.n5344 VSS.n5345 0.147342
R9060 VSS.n5351 VSS.n5347 0.0722544
R9061 VSS.n5352 VSS.n5348 4.5005
R9062 VSS.n5353 VSS.n5349 4.5005
R9063 VSS.n5354 VSS.n5350 4.5005
R9064 VSS.n5351 VSS.n5340 4.57426
R9065 VSS.n5347 VSS.n5348 0.147342
R9066 VSS.n5348 VSS.n5349 0.147342
R9067 VSS.n5349 VSS.n5350 0.147342
R9068 VSS.n5352 VSS.n5351 2.37296
R9069 VSS.n5353 VSS.n5352 0.127318
R9070 VSS.n5354 VSS.n5353 0.127318
R9071 VSS.t0 VSS.n5354 2.73618
R9072 VSS.n5327 VSS.n5332 4.5005
R9073 VSS.n5329 VSS.n5333 4.5005
R9074 VSS.n5330 VSS.n5334 4.5005
R9075 VSS.n5331 VSS.n5335 4.57324
R9076 VSS.n5327 VSS.n5325 0.147342
R9077 VSS.n5328 VSS.n5329 0.0732424
R9078 VSS.n5329 VSS.n5330 0.147342
R9079 VSS.n5332 VSS.n5336 0.0721009
R9080 VSS.n5337 VSS.n5333 4.5005
R9081 VSS.n5338 VSS.n5334 4.5005
R9082 VSS.n5339 VSS.n5335 4.5005
R9083 VSS.n5325 VSS.n5336 4.57442
R9084 VSS.n5332 VSS.n5333 0.147342
R9085 VSS.n5333 VSS.n5334 0.147342
R9086 VSS.n5334 VSS.n5335 0.147342
R9087 VSS.n5336 VSS.n5337 2.39784
R9088 VSS.n5337 VSS.n5338 0.147342
R9089 VSS.n5338 VSS.n5339 0.147342
R9090 VSS.n5339 VSS.t549 3.13212
R9091 VSS.n5312 VSS.n5317 4.5005
R9092 VSS.n5314 VSS.n5318 4.5005
R9093 VSS.n5315 VSS.n5319 4.5005
R9094 VSS.n5316 VSS.n5320 4.57324
R9095 VSS.n5312 VSS.n5310 0.147342
R9096 VSS.n5313 VSS.n5314 0.0732424
R9097 VSS.n5314 VSS.n5315 0.147342
R9098 VSS.n5317 VSS.n5321 0.0721009
R9099 VSS.n5322 VSS.n5318 4.5005
R9100 VSS.n5323 VSS.n5319 4.5005
R9101 VSS.n5324 VSS.n5320 4.5005
R9102 VSS.n5310 VSS.n5321 4.57442
R9103 VSS.n5317 VSS.n5318 0.147342
R9104 VSS.n5318 VSS.n5319 0.147342
R9105 VSS.n5319 VSS.n5320 0.147342
R9106 VSS.n5321 VSS.n5322 2.39784
R9107 VSS.n5322 VSS.n5323 0.147342
R9108 VSS.n5323 VSS.n5324 0.147342
R9109 VSS.n5324 VSS.t255 3.13212
R9110 VSS.n5297 VSS.n5302 4.5005
R9111 VSS.n5299 VSS.n5303 4.5005
R9112 VSS.n5300 VSS.n5304 4.5005
R9113 VSS.n5301 VSS.n5305 4.57324
R9114 VSS.n5297 VSS.n5295 0.147342
R9115 VSS.n5298 VSS.n5299 0.0732424
R9116 VSS.n5299 VSS.n5300 0.147342
R9117 VSS.n5302 VSS.n5306 0.0721009
R9118 VSS.n5307 VSS.n5303 4.5005
R9119 VSS.n5308 VSS.n5304 4.5005
R9120 VSS.n5309 VSS.n5305 4.5005
R9121 VSS.n5295 VSS.n5306 4.57442
R9122 VSS.n5302 VSS.n5303 0.147342
R9123 VSS.n5303 VSS.n5304 0.147342
R9124 VSS.n5304 VSS.n5305 0.147342
R9125 VSS.n5306 VSS.n5307 2.39784
R9126 VSS.n5307 VSS.n5308 0.147342
R9127 VSS.n5308 VSS.n5309 0.147342
R9128 VSS.n5309 VSS.t432 3.13212
R9129 VSS.n5287 VSS.n5282 4.5005
R9130 VSS.n5288 VSS.n5284 4.5005
R9131 VSS.n5289 VSS.n5285 4.5005
R9132 VSS.n5290 VSS.n5286 4.57324
R9133 VSS.n5280 VSS.n5282 0.147342
R9134 VSS.n5283 VSS.n5284 0.0732424
R9135 VSS.n5284 VSS.n5285 0.147342
R9136 VSS.n5291 VSS.n5287 0.0722544
R9137 VSS.n5292 VSS.n5288 4.5005
R9138 VSS.n5293 VSS.n5289 4.5005
R9139 VSS.n5294 VSS.n5290 4.5005
R9140 VSS.n5291 VSS.n5280 4.57426
R9141 VSS.n5287 VSS.n5288 0.147342
R9142 VSS.n5288 VSS.n5289 0.147342
R9143 VSS.n5289 VSS.n5290 0.147342
R9144 VSS.n5292 VSS.n5291 2.37296
R9145 VSS.n5293 VSS.n5292 0.127318
R9146 VSS.n5294 VSS.n5293 0.127318
R9147 VSS.t0 VSS.n5294 2.73618
R9148 VSS.n5267 VSS.n5272 4.5005
R9149 VSS.n5269 VSS.n5273 4.5005
R9150 VSS.n5270 VSS.n5274 4.5005
R9151 VSS.n5271 VSS.n5275 4.57324
R9152 VSS.n5267 VSS.n5265 0.147342
R9153 VSS.n5268 VSS.n5269 0.0732424
R9154 VSS.n5269 VSS.n5270 0.147342
R9155 VSS.n5272 VSS.n5276 0.0721009
R9156 VSS.n5277 VSS.n5273 4.5005
R9157 VSS.n5278 VSS.n5274 4.5005
R9158 VSS.n5279 VSS.n5275 4.5005
R9159 VSS.n5265 VSS.n5276 4.57442
R9160 VSS.n5272 VSS.n5273 0.147342
R9161 VSS.n5273 VSS.n5274 0.147342
R9162 VSS.n5274 VSS.n5275 0.147342
R9163 VSS.n5276 VSS.n5277 2.39784
R9164 VSS.n5277 VSS.n5278 0.147342
R9165 VSS.n5278 VSS.n5279 0.147342
R9166 VSS.n5279 VSS.t442 3.13212
R9167 VSS.n5252 VSS.n5257 4.5005
R9168 VSS.n5254 VSS.n5258 4.5005
R9169 VSS.n5255 VSS.n5259 4.5005
R9170 VSS.n5256 VSS.n5260 4.57324
R9171 VSS.n5252 VSS.n5250 0.147342
R9172 VSS.n5253 VSS.n5254 0.0732424
R9173 VSS.n5254 VSS.n5255 0.147342
R9174 VSS.n5257 VSS.n5261 0.0721009
R9175 VSS.n5262 VSS.n5258 4.5005
R9176 VSS.n5263 VSS.n5259 4.5005
R9177 VSS.n5264 VSS.n5260 4.5005
R9178 VSS.n5250 VSS.n5261 4.57442
R9179 VSS.n5257 VSS.n5258 0.147342
R9180 VSS.n5258 VSS.n5259 0.147342
R9181 VSS.n5259 VSS.n5260 0.147342
R9182 VSS.n5261 VSS.n5262 2.39784
R9183 VSS.n5262 VSS.n5263 0.147342
R9184 VSS.n5263 VSS.n5264 0.147342
R9185 VSS.n5264 VSS.t156 3.13212
R9186 VSS.n5237 VSS.n5242 4.5005
R9187 VSS.n5239 VSS.n5243 4.5005
R9188 VSS.n5240 VSS.n5244 4.5005
R9189 VSS.n5241 VSS.n5245 4.57324
R9190 VSS.n5237 VSS.n5235 0.147342
R9191 VSS.n5238 VSS.n5239 0.0732424
R9192 VSS.n5239 VSS.n5240 0.147342
R9193 VSS.n5242 VSS.n5246 0.0721009
R9194 VSS.n5247 VSS.n5243 4.5005
R9195 VSS.n5248 VSS.n5244 4.5005
R9196 VSS.n5249 VSS.n5245 4.5005
R9197 VSS.n5235 VSS.n5246 4.57442
R9198 VSS.n5242 VSS.n5243 0.147342
R9199 VSS.n5243 VSS.n5244 0.147342
R9200 VSS.n5244 VSS.n5245 0.147342
R9201 VSS.n5246 VSS.n5247 2.39784
R9202 VSS.n5247 VSS.n5248 0.147342
R9203 VSS.n5248 VSS.n5249 0.147342
R9204 VSS.n5249 VSS.t179 3.13212
R9205 VSS.n5222 VSS.n5227 4.5005
R9206 VSS.n5224 VSS.n5228 4.5005
R9207 VSS.n5225 VSS.n5229 4.5005
R9208 VSS.n5226 VSS.n5230 4.57324
R9209 VSS.n5222 VSS.n5220 0.147342
R9210 VSS.n5223 VSS.n5224 0.0732424
R9211 VSS.n5224 VSS.n5225 0.147342
R9212 VSS.n5227 VSS.n5231 0.0721009
R9213 VSS.n5232 VSS.n5228 4.5005
R9214 VSS.n5233 VSS.n5229 4.5005
R9215 VSS.n5234 VSS.n5230 4.5005
R9216 VSS.n5220 VSS.n5231 4.57442
R9217 VSS.n5227 VSS.n5228 0.147342
R9218 VSS.n5228 VSS.n5229 0.147342
R9219 VSS.n5229 VSS.n5230 0.147342
R9220 VSS.n5231 VSS.n5232 2.39784
R9221 VSS.n5232 VSS.n5233 0.147342
R9222 VSS.n5233 VSS.n5234 0.147342
R9223 VSS.n5234 VSS.t98 3.13212
R9224 VSS.n5207 VSS.n5212 4.5005
R9225 VSS.n5209 VSS.n5213 4.5005
R9226 VSS.n5210 VSS.n5214 4.5005
R9227 VSS.n5211 VSS.n5215 4.57324
R9228 VSS.n5207 VSS.n5205 0.147342
R9229 VSS.n5208 VSS.n5209 0.0732424
R9230 VSS.n5209 VSS.n5210 0.147342
R9231 VSS.n5212 VSS.n5216 0.0721009
R9232 VSS.n5217 VSS.n5213 4.5005
R9233 VSS.n5218 VSS.n5214 4.5005
R9234 VSS.n5219 VSS.n5215 4.5005
R9235 VSS.n5205 VSS.n5216 4.57442
R9236 VSS.n5212 VSS.n5213 0.147342
R9237 VSS.n5213 VSS.n5214 0.147342
R9238 VSS.n5214 VSS.n5215 0.147342
R9239 VSS.n5216 VSS.n5217 2.39784
R9240 VSS.n5217 VSS.n5218 0.147342
R9241 VSS.n5218 VSS.n5219 0.147342
R9242 VSS.n5219 VSS.t481 3.13212
R9243 VSS.n5192 VSS.n5197 4.5005
R9244 VSS.n5194 VSS.n5198 4.5005
R9245 VSS.n5195 VSS.n5199 4.5005
R9246 VSS.n5196 VSS.n5200 4.57324
R9247 VSS.n5192 VSS.n5190 0.147342
R9248 VSS.n5193 VSS.n5194 0.0732424
R9249 VSS.n5194 VSS.n5195 0.147342
R9250 VSS.n5197 VSS.n5201 0.0721009
R9251 VSS.n5202 VSS.n5198 4.5005
R9252 VSS.n5203 VSS.n5199 4.5005
R9253 VSS.n5204 VSS.n5200 4.5005
R9254 VSS.n5190 VSS.n5201 4.57442
R9255 VSS.n5197 VSS.n5198 0.147342
R9256 VSS.n5198 VSS.n5199 0.147342
R9257 VSS.n5199 VSS.n5200 0.147342
R9258 VSS.n5201 VSS.n5202 2.39784
R9259 VSS.n5202 VSS.n5203 0.147342
R9260 VSS.n5203 VSS.n5204 0.147342
R9261 VSS.n5204 VSS.t61 3.13212
R9262 VSS.n5182 VSS.n5177 4.5005
R9263 VSS.n5183 VSS.n5179 4.5005
R9264 VSS.n5184 VSS.n5180 4.5005
R9265 VSS.n5185 VSS.n5181 4.57324
R9266 VSS.n5175 VSS.n5177 0.147342
R9267 VSS.n5178 VSS.n5179 0.0732424
R9268 VSS.n5179 VSS.n5180 0.147342
R9269 VSS.n5186 VSS.n5182 0.0722544
R9270 VSS.n5187 VSS.n5183 4.5005
R9271 VSS.n5188 VSS.n5184 4.5005
R9272 VSS.n5189 VSS.n5185 4.5005
R9273 VSS.n5186 VSS.n5175 4.57426
R9274 VSS.n5182 VSS.n5183 0.147342
R9275 VSS.n5183 VSS.n5184 0.147342
R9276 VSS.n5184 VSS.n5185 0.147342
R9277 VSS.n5187 VSS.n5186 2.37296
R9278 VSS.n5188 VSS.n5187 0.127318
R9279 VSS.n5189 VSS.n5188 0.127318
R9280 VSS.t0 VSS.n5189 2.73618
R9281 VSS.n5162 VSS.n5167 4.5005
R9282 VSS.n5164 VSS.n5168 4.5005
R9283 VSS.n5165 VSS.n5169 4.5005
R9284 VSS.n5166 VSS.n5170 4.57324
R9285 VSS.n5162 VSS.n5160 0.147342
R9286 VSS.n5163 VSS.n5164 0.0732424
R9287 VSS.n5164 VSS.n5165 0.147342
R9288 VSS.n5167 VSS.n5171 0.0721009
R9289 VSS.n5172 VSS.n5168 4.5005
R9290 VSS.n5173 VSS.n5169 4.5005
R9291 VSS.n5174 VSS.n5170 4.5005
R9292 VSS.n5160 VSS.n5171 4.57442
R9293 VSS.n5167 VSS.n5168 0.147342
R9294 VSS.n5168 VSS.n5169 0.147342
R9295 VSS.n5169 VSS.n5170 0.147342
R9296 VSS.n5171 VSS.n5172 2.39784
R9297 VSS.n5172 VSS.n5173 0.147342
R9298 VSS.n5173 VSS.n5174 0.147342
R9299 VSS.n5174 VSS.t218 3.13212
R9300 VSS.n5147 VSS.n5152 4.5005
R9301 VSS.n5149 VSS.n5153 4.5005
R9302 VSS.n5150 VSS.n5154 4.5005
R9303 VSS.n5151 VSS.n5155 4.57324
R9304 VSS.n5147 VSS.n5145 0.147342
R9305 VSS.n5148 VSS.n5149 0.0732424
R9306 VSS.n5149 VSS.n5150 0.147342
R9307 VSS.n5152 VSS.n5156 0.0721009
R9308 VSS.n5157 VSS.n5153 4.5005
R9309 VSS.n5158 VSS.n5154 4.5005
R9310 VSS.n5159 VSS.n5155 4.5005
R9311 VSS.n5145 VSS.n5156 4.57442
R9312 VSS.n5152 VSS.n5153 0.147342
R9313 VSS.n5153 VSS.n5154 0.147342
R9314 VSS.n5154 VSS.n5155 0.147342
R9315 VSS.n5156 VSS.n5157 2.39784
R9316 VSS.n5157 VSS.n5158 0.147342
R9317 VSS.n5158 VSS.n5159 0.147342
R9318 VSS.n5159 VSS.t212 3.13212
R9319 VSS.n5132 VSS.n5137 4.5005
R9320 VSS.n5134 VSS.n5138 4.5005
R9321 VSS.n5135 VSS.n5139 4.5005
R9322 VSS.n5136 VSS.n5140 4.57324
R9323 VSS.n5132 VSS.n5130 0.147342
R9324 VSS.n5133 VSS.n5134 0.0732424
R9325 VSS.n5134 VSS.n5135 0.147342
R9326 VSS.n5137 VSS.n5141 0.0721009
R9327 VSS.n5142 VSS.n5138 4.5005
R9328 VSS.n5143 VSS.n5139 4.5005
R9329 VSS.n5144 VSS.n5140 4.5005
R9330 VSS.n5130 VSS.n5141 4.57442
R9331 VSS.n5137 VSS.n5138 0.147342
R9332 VSS.n5138 VSS.n5139 0.147342
R9333 VSS.n5139 VSS.n5140 0.147342
R9334 VSS.n5141 VSS.n5142 2.39784
R9335 VSS.n5142 VSS.n5143 0.147342
R9336 VSS.n5143 VSS.n5144 0.147342
R9337 VSS.n5144 VSS.t235 3.13212
R9338 VSS.n5122 VSS.n5117 4.5005
R9339 VSS.n5123 VSS.n5119 4.5005
R9340 VSS.n5124 VSS.n5120 4.5005
R9341 VSS.n5125 VSS.n5121 4.57324
R9342 VSS.n5115 VSS.n5117 0.147342
R9343 VSS.n5118 VSS.n5119 0.0732424
R9344 VSS.n5119 VSS.n5120 0.147342
R9345 VSS.n5126 VSS.n5122 0.0722544
R9346 VSS.n5127 VSS.n5123 4.5005
R9347 VSS.n5128 VSS.n5124 4.5005
R9348 VSS.n5129 VSS.n5125 4.5005
R9349 VSS.n5126 VSS.n5115 4.57426
R9350 VSS.n5122 VSS.n5123 0.147342
R9351 VSS.n5123 VSS.n5124 0.147342
R9352 VSS.n5124 VSS.n5125 0.147342
R9353 VSS.n5127 VSS.n5126 2.37296
R9354 VSS.n5128 VSS.n5127 0.127318
R9355 VSS.n5129 VSS.n5128 0.127318
R9356 VSS.t0 VSS.n5129 2.73618
R9357 VSS.n5102 VSS.n5107 4.5005
R9358 VSS.n5104 VSS.n5108 4.5005
R9359 VSS.n5105 VSS.n5109 4.5005
R9360 VSS.n5106 VSS.n5110 4.57324
R9361 VSS.n5102 VSS.n5100 0.147342
R9362 VSS.n5103 VSS.n5104 0.0732424
R9363 VSS.n5104 VSS.n5105 0.147342
R9364 VSS.n5107 VSS.n5111 0.0721009
R9365 VSS.n5112 VSS.n5108 4.5005
R9366 VSS.n5113 VSS.n5109 4.5005
R9367 VSS.n5114 VSS.n5110 4.5005
R9368 VSS.n5100 VSS.n5111 4.57442
R9369 VSS.n5107 VSS.n5108 0.147342
R9370 VSS.n5108 VSS.n5109 0.147342
R9371 VSS.n5109 VSS.n5110 0.147342
R9372 VSS.n5111 VSS.n5112 2.39784
R9373 VSS.n5112 VSS.n5113 0.147342
R9374 VSS.n5113 VSS.n5114 0.147342
R9375 VSS.n5114 VSS.t39 3.13212
R9376 VSS.n5087 VSS.n5092 4.5005
R9377 VSS.n5089 VSS.n5093 4.5005
R9378 VSS.n5090 VSS.n5094 4.5005
R9379 VSS.n5091 VSS.n5095 4.57324
R9380 VSS.n5087 VSS.n5085 0.147342
R9381 VSS.n5088 VSS.n5089 0.0732424
R9382 VSS.n5089 VSS.n5090 0.147342
R9383 VSS.n5092 VSS.n5096 0.0721009
R9384 VSS.n5097 VSS.n5093 4.5005
R9385 VSS.n5098 VSS.n5094 4.5005
R9386 VSS.n5099 VSS.n5095 4.5005
R9387 VSS.n5085 VSS.n5096 4.57442
R9388 VSS.n5092 VSS.n5093 0.147342
R9389 VSS.n5093 VSS.n5094 0.147342
R9390 VSS.n5094 VSS.n5095 0.147342
R9391 VSS.n5096 VSS.n5097 2.39784
R9392 VSS.n5097 VSS.n5098 0.147342
R9393 VSS.n5098 VSS.n5099 0.147342
R9394 VSS.n5099 VSS.t4 3.13212
R9395 VSS.n5072 VSS.n5077 4.5005
R9396 VSS.n5074 VSS.n5078 4.5005
R9397 VSS.n5075 VSS.n5079 4.5005
R9398 VSS.n5076 VSS.n5080 4.57324
R9399 VSS.n5072 VSS.n5070 0.147342
R9400 VSS.n5073 VSS.n5074 0.0732424
R9401 VSS.n5074 VSS.n5075 0.147342
R9402 VSS.n5077 VSS.n5081 0.0721009
R9403 VSS.n5082 VSS.n5078 4.5005
R9404 VSS.n5083 VSS.n5079 4.5005
R9405 VSS.n5084 VSS.n5080 4.5005
R9406 VSS.n5070 VSS.n5081 4.57442
R9407 VSS.n5077 VSS.n5078 0.147342
R9408 VSS.n5078 VSS.n5079 0.147342
R9409 VSS.n5079 VSS.n5080 0.147342
R9410 VSS.n5081 VSS.n5082 2.39784
R9411 VSS.n5082 VSS.n5083 0.147342
R9412 VSS.n5083 VSS.n5084 0.147342
R9413 VSS.n5084 VSS.t286 3.13212
R9414 VSS.n5057 VSS.n5062 4.5005
R9415 VSS.n5059 VSS.n5063 4.5005
R9416 VSS.n5060 VSS.n5064 4.5005
R9417 VSS.n5061 VSS.n5065 4.57324
R9418 VSS.n5057 VSS.n5055 0.147342
R9419 VSS.n5058 VSS.n5059 0.0732424
R9420 VSS.n5059 VSS.n5060 0.147342
R9421 VSS.n5062 VSS.n5066 0.0721009
R9422 VSS.n5067 VSS.n5063 4.5005
R9423 VSS.n5068 VSS.n5064 4.5005
R9424 VSS.n5069 VSS.n5065 4.5005
R9425 VSS.n5055 VSS.n5066 4.57442
R9426 VSS.n5062 VSS.n5063 0.147342
R9427 VSS.n5063 VSS.n5064 0.147342
R9428 VSS.n5064 VSS.n5065 0.147342
R9429 VSS.n5066 VSS.n5067 2.39784
R9430 VSS.n5067 VSS.n5068 0.147342
R9431 VSS.n5068 VSS.n5069 0.147342
R9432 VSS.n5069 VSS.t294 3.13212
R9433 VSS.n5047 VSS.n5042 4.5005
R9434 VSS.n5048 VSS.n5044 4.5005
R9435 VSS.n5049 VSS.n5045 4.5005
R9436 VSS.n5050 VSS.n5046 4.57324
R9437 VSS.n5040 VSS.n5042 0.147342
R9438 VSS.n5043 VSS.n5044 0.0732424
R9439 VSS.n5044 VSS.n5045 0.147342
R9440 VSS.n5051 VSS.n5047 0.0722544
R9441 VSS.n5052 VSS.n5048 4.5005
R9442 VSS.n5053 VSS.n5049 4.5005
R9443 VSS.n5054 VSS.n5050 4.5005
R9444 VSS.n5051 VSS.n5040 4.57426
R9445 VSS.n5047 VSS.n5048 0.147342
R9446 VSS.n5048 VSS.n5049 0.147342
R9447 VSS.n5049 VSS.n5050 0.147342
R9448 VSS.n5052 VSS.n5051 2.37296
R9449 VSS.n5053 VSS.n5052 0.127318
R9450 VSS.n5054 VSS.n5053 0.127318
R9451 VSS.t0 VSS.n5054 2.73618
R9452 VSS.n5027 VSS.n5032 4.5005
R9453 VSS.n5029 VSS.n5033 4.5005
R9454 VSS.n5030 VSS.n5034 4.5005
R9455 VSS.n5031 VSS.n5035 4.57324
R9456 VSS.n5027 VSS.n5025 0.147342
R9457 VSS.n5028 VSS.n5029 0.0732424
R9458 VSS.n5029 VSS.n5030 0.147342
R9459 VSS.n5032 VSS.n5036 0.0721009
R9460 VSS.n5037 VSS.n5033 4.5005
R9461 VSS.n5038 VSS.n5034 4.5005
R9462 VSS.n5039 VSS.n5035 4.5005
R9463 VSS.n5025 VSS.n5036 4.57442
R9464 VSS.n5032 VSS.n5033 0.147342
R9465 VSS.n5033 VSS.n5034 0.147342
R9466 VSS.n5034 VSS.n5035 0.147342
R9467 VSS.n5036 VSS.n5037 2.39784
R9468 VSS.n5037 VSS.n5038 0.147342
R9469 VSS.n5038 VSS.n5039 0.147342
R9470 VSS.n5039 VSS.t544 3.13212
R9471 VSS.n5012 VSS.n5017 4.5005
R9472 VSS.n5014 VSS.n5018 4.5005
R9473 VSS.n5015 VSS.n5019 4.5005
R9474 VSS.n5016 VSS.n5020 4.57324
R9475 VSS.n5012 VSS.n5010 0.147342
R9476 VSS.n5013 VSS.n5014 0.0732424
R9477 VSS.n5014 VSS.n5015 0.147342
R9478 VSS.n5017 VSS.n5021 0.0721009
R9479 VSS.n5022 VSS.n5018 4.5005
R9480 VSS.n5023 VSS.n5019 4.5005
R9481 VSS.n5024 VSS.n5020 4.5005
R9482 VSS.n5010 VSS.n5021 4.57442
R9483 VSS.n5017 VSS.n5018 0.147342
R9484 VSS.n5018 VSS.n5019 0.147342
R9485 VSS.n5019 VSS.n5020 0.147342
R9486 VSS.n5021 VSS.n5022 2.39784
R9487 VSS.n5022 VSS.n5023 0.147342
R9488 VSS.n5023 VSS.n5024 0.147342
R9489 VSS.n5024 VSS.t257 3.13212
R9490 VSS.n4997 VSS.n5002 4.5005
R9491 VSS.n4999 VSS.n5003 4.5005
R9492 VSS.n5000 VSS.n5004 4.5005
R9493 VSS.n5001 VSS.n5005 4.57324
R9494 VSS.n4997 VSS.n4995 0.147342
R9495 VSS.n4998 VSS.n4999 0.0732424
R9496 VSS.n4999 VSS.n5000 0.147342
R9497 VSS.n5002 VSS.n5006 0.0721009
R9498 VSS.n5007 VSS.n5003 4.5005
R9499 VSS.n5008 VSS.n5004 4.5005
R9500 VSS.n5009 VSS.n5005 4.5005
R9501 VSS.n4995 VSS.n5006 4.57442
R9502 VSS.n5002 VSS.n5003 0.147342
R9503 VSS.n5003 VSS.n5004 0.147342
R9504 VSS.n5004 VSS.n5005 0.147342
R9505 VSS.n5006 VSS.n5007 2.39784
R9506 VSS.n5007 VSS.n5008 0.147342
R9507 VSS.n5008 VSS.n5009 0.147342
R9508 VSS.n5009 VSS.t538 3.13212
R9509 VSS.n4987 VSS.n4982 4.5005
R9510 VSS.n4988 VSS.n4984 4.5005
R9511 VSS.n4989 VSS.n4985 4.5005
R9512 VSS.n4990 VSS.n4986 4.57324
R9513 VSS.n4980 VSS.n4982 0.147342
R9514 VSS.n4983 VSS.n4984 0.0732424
R9515 VSS.n4984 VSS.n4985 0.147342
R9516 VSS.n4991 VSS.n4987 0.0722544
R9517 VSS.n4992 VSS.n4988 4.5005
R9518 VSS.n4993 VSS.n4989 4.5005
R9519 VSS.n4994 VSS.n4990 4.5005
R9520 VSS.n4991 VSS.n4980 4.57426
R9521 VSS.n4987 VSS.n4988 0.147342
R9522 VSS.n4988 VSS.n4989 0.147342
R9523 VSS.n4989 VSS.n4990 0.147342
R9524 VSS.n4992 VSS.n4991 2.37296
R9525 VSS.n4993 VSS.n4992 0.127318
R9526 VSS.n4994 VSS.n4993 0.127318
R9527 VSS.t0 VSS.n4994 2.73618
R9528 VSS.n4967 VSS.n4972 4.5005
R9529 VSS.n4969 VSS.n4973 4.5005
R9530 VSS.n4970 VSS.n4974 4.5005
R9531 VSS.n4971 VSS.n4975 4.57324
R9532 VSS.n4967 VSS.n4965 0.147342
R9533 VSS.n4968 VSS.n4969 0.0732424
R9534 VSS.n4969 VSS.n4970 0.147342
R9535 VSS.n4972 VSS.n4976 0.0721009
R9536 VSS.n4977 VSS.n4973 4.5005
R9537 VSS.n4978 VSS.n4974 4.5005
R9538 VSS.n4979 VSS.n4975 4.5005
R9539 VSS.n4965 VSS.n4976 4.57442
R9540 VSS.n4972 VSS.n4973 0.147342
R9541 VSS.n4973 VSS.n4974 0.147342
R9542 VSS.n4974 VSS.n4975 0.147342
R9543 VSS.n4976 VSS.n4977 2.39784
R9544 VSS.n4977 VSS.n4978 0.147342
R9545 VSS.n4978 VSS.n4979 0.147342
R9546 VSS.n4979 VSS.t1 3.13212
R9547 VSS.n4952 VSS.n4957 4.5005
R9548 VSS.n4954 VSS.n4958 4.5005
R9549 VSS.n4955 VSS.n4959 4.5005
R9550 VSS.n4956 VSS.n4960 4.57324
R9551 VSS.n4952 VSS.n4950 0.147342
R9552 VSS.n4953 VSS.n4954 0.0732424
R9553 VSS.n4954 VSS.n4955 0.147342
R9554 VSS.n4957 VSS.n4961 0.0721009
R9555 VSS.n4962 VSS.n4958 4.5005
R9556 VSS.n4963 VSS.n4959 4.5005
R9557 VSS.n4964 VSS.n4960 4.5005
R9558 VSS.n4950 VSS.n4961 4.57442
R9559 VSS.n4957 VSS.n4958 0.147342
R9560 VSS.n4958 VSS.n4959 0.147342
R9561 VSS.n4959 VSS.n4960 0.147342
R9562 VSS.n4961 VSS.n4962 2.39784
R9563 VSS.n4962 VSS.n4963 0.147342
R9564 VSS.n4963 VSS.n4964 0.147342
R9565 VSS.n4964 VSS.t158 3.13212
R9566 VSS.n4937 VSS.n4942 4.5005
R9567 VSS.n4939 VSS.n4943 4.5005
R9568 VSS.n4940 VSS.n4944 4.5005
R9569 VSS.n4941 VSS.n4945 4.57324
R9570 VSS.n4937 VSS.n4935 0.147342
R9571 VSS.n4938 VSS.n4939 0.0732424
R9572 VSS.n4939 VSS.n4940 0.147342
R9573 VSS.n4942 VSS.n4946 0.0721009
R9574 VSS.n4947 VSS.n4943 4.5005
R9575 VSS.n4948 VSS.n4944 4.5005
R9576 VSS.n4949 VSS.n4945 4.5005
R9577 VSS.n4935 VSS.n4946 4.57442
R9578 VSS.n4942 VSS.n4943 0.147342
R9579 VSS.n4943 VSS.n4944 0.147342
R9580 VSS.n4944 VSS.n4945 0.147342
R9581 VSS.n4946 VSS.n4947 2.39784
R9582 VSS.n4947 VSS.n4948 0.147342
R9583 VSS.n4948 VSS.n4949 0.147342
R9584 VSS.n4949 VSS.t263 3.13212
R9585 VSS.n4922 VSS.n4927 4.5005
R9586 VSS.n4924 VSS.n4928 4.5005
R9587 VSS.n4925 VSS.n4929 4.5005
R9588 VSS.n4926 VSS.n4930 4.57324
R9589 VSS.n4922 VSS.n4920 0.147342
R9590 VSS.n4923 VSS.n4924 0.0732424
R9591 VSS.n4924 VSS.n4925 0.147342
R9592 VSS.n4927 VSS.n4931 0.0721009
R9593 VSS.n4932 VSS.n4928 4.5005
R9594 VSS.n4933 VSS.n4929 4.5005
R9595 VSS.n4934 VSS.n4930 4.5005
R9596 VSS.n4920 VSS.n4931 4.57442
R9597 VSS.n4927 VSS.n4928 0.147342
R9598 VSS.n4928 VSS.n4929 0.147342
R9599 VSS.n4929 VSS.n4930 0.147342
R9600 VSS.n4931 VSS.n4932 2.39784
R9601 VSS.n4932 VSS.n4933 0.147342
R9602 VSS.n4933 VSS.n4934 0.147342
R9603 VSS.n4934 VSS.t95 3.13212
R9604 VSS.n4907 VSS.n4912 4.5005
R9605 VSS.n4909 VSS.n4913 4.5005
R9606 VSS.n4910 VSS.n4914 4.5005
R9607 VSS.n4911 VSS.n4915 4.57324
R9608 VSS.n4907 VSS.n4905 0.147342
R9609 VSS.n4908 VSS.n4909 0.0732424
R9610 VSS.n4909 VSS.n4910 0.147342
R9611 VSS.n4912 VSS.n4916 0.0721009
R9612 VSS.n4917 VSS.n4913 4.5005
R9613 VSS.n4918 VSS.n4914 4.5005
R9614 VSS.n4919 VSS.n4915 4.5005
R9615 VSS.n4905 VSS.n4916 4.57442
R9616 VSS.n4912 VSS.n4913 0.147342
R9617 VSS.n4913 VSS.n4914 0.147342
R9618 VSS.n4914 VSS.n4915 0.147342
R9619 VSS.n4916 VSS.n4917 2.39784
R9620 VSS.n4917 VSS.n4918 0.147342
R9621 VSS.n4918 VSS.n4919 0.147342
R9622 VSS.n4919 VSS.t483 3.13212
R9623 VSS.n4892 VSS.n4897 4.5005
R9624 VSS.n4894 VSS.n4898 4.5005
R9625 VSS.n4895 VSS.n4899 4.5005
R9626 VSS.n4896 VSS.n4900 4.57324
R9627 VSS.n4892 VSS.n4890 0.147342
R9628 VSS.n4893 VSS.n4894 0.0732424
R9629 VSS.n4894 VSS.n4895 0.147342
R9630 VSS.n4897 VSS.n4901 0.0721009
R9631 VSS.n4902 VSS.n4898 4.5005
R9632 VSS.n4903 VSS.n4899 4.5005
R9633 VSS.n4904 VSS.n4900 4.5005
R9634 VSS.n4890 VSS.n4901 4.57442
R9635 VSS.n4897 VSS.n4898 0.147342
R9636 VSS.n4898 VSS.n4899 0.147342
R9637 VSS.n4899 VSS.n4900 0.147342
R9638 VSS.n4901 VSS.n4902 2.39784
R9639 VSS.n4902 VSS.n4903 0.147342
R9640 VSS.n4903 VSS.n4904 0.147342
R9641 VSS.n4904 VSS.t63 3.13212
R9642 VSS.n4882 VSS.n4877 4.5005
R9643 VSS.n4883 VSS.n4879 4.5005
R9644 VSS.n4884 VSS.n4880 4.5005
R9645 VSS.n4885 VSS.n4881 4.57324
R9646 VSS.n4875 VSS.n4877 0.147342
R9647 VSS.n4878 VSS.n4879 0.0732424
R9648 VSS.n4879 VSS.n4880 0.147342
R9649 VSS.n4886 VSS.n4882 0.0722544
R9650 VSS.n4887 VSS.n4883 4.5005
R9651 VSS.n4888 VSS.n4884 4.5005
R9652 VSS.n4889 VSS.n4885 4.5005
R9653 VSS.n4886 VSS.n4875 4.57426
R9654 VSS.n4882 VSS.n4883 0.147342
R9655 VSS.n4883 VSS.n4884 0.147342
R9656 VSS.n4884 VSS.n4885 0.147342
R9657 VSS.n4887 VSS.n4886 2.37296
R9658 VSS.n4888 VSS.n4887 0.127318
R9659 VSS.n4889 VSS.n4888 0.127318
R9660 VSS.t0 VSS.n4889 2.73618
R9661 VSS.n4862 VSS.n4867 4.5005
R9662 VSS.n4864 VSS.n4868 4.5005
R9663 VSS.n4865 VSS.n4869 4.5005
R9664 VSS.n4866 VSS.n4870 4.57324
R9665 VSS.n4862 VSS.n4860 0.147342
R9666 VSS.n4863 VSS.n4864 0.0732424
R9667 VSS.n4864 VSS.n4865 0.147342
R9668 VSS.n4867 VSS.n4871 0.0721009
R9669 VSS.n4872 VSS.n4868 4.5005
R9670 VSS.n4873 VSS.n4869 4.5005
R9671 VSS.n4874 VSS.n4870 4.5005
R9672 VSS.n4860 VSS.n4871 4.57442
R9673 VSS.n4867 VSS.n4868 0.147342
R9674 VSS.n4868 VSS.n4869 0.147342
R9675 VSS.n4869 VSS.n4870 0.147342
R9676 VSS.n4871 VSS.n4872 2.39784
R9677 VSS.n4872 VSS.n4873 0.147342
R9678 VSS.n4873 VSS.n4874 0.147342
R9679 VSS.n4874 VSS.t34 3.13212
R9680 VSS.n4847 VSS.n4852 4.5005
R9681 VSS.n4849 VSS.n4853 4.5005
R9682 VSS.n4850 VSS.n4854 4.5005
R9683 VSS.n4851 VSS.n4855 4.57324
R9684 VSS.n4847 VSS.n4845 0.147342
R9685 VSS.n4848 VSS.n4849 0.0732424
R9686 VSS.n4849 VSS.n4850 0.147342
R9687 VSS.n4852 VSS.n4856 0.0721009
R9688 VSS.n4857 VSS.n4853 4.5005
R9689 VSS.n4858 VSS.n4854 4.5005
R9690 VSS.n4859 VSS.n4855 4.5005
R9691 VSS.n4845 VSS.n4856 4.57442
R9692 VSS.n4852 VSS.n4853 0.147342
R9693 VSS.n4853 VSS.n4854 0.147342
R9694 VSS.n4854 VSS.n4855 0.147342
R9695 VSS.n4856 VSS.n4857 2.39784
R9696 VSS.n4857 VSS.n4858 0.147342
R9697 VSS.n4858 VSS.n4859 0.147342
R9698 VSS.n4859 VSS.t210 3.13212
R9699 VSS.n4832 VSS.n4837 4.5005
R9700 VSS.n4834 VSS.n4838 4.5005
R9701 VSS.n4835 VSS.n4839 4.5005
R9702 VSS.n4836 VSS.n4840 4.57324
R9703 VSS.n4832 VSS.n4830 0.147342
R9704 VSS.n4833 VSS.n4834 0.0732424
R9705 VSS.n4834 VSS.n4835 0.147342
R9706 VSS.n4837 VSS.n4841 0.0721009
R9707 VSS.n4842 VSS.n4838 4.5005
R9708 VSS.n4843 VSS.n4839 4.5005
R9709 VSS.n4844 VSS.n4840 4.5005
R9710 VSS.n4830 VSS.n4841 4.57442
R9711 VSS.n4837 VSS.n4838 0.147342
R9712 VSS.n4838 VSS.n4839 0.147342
R9713 VSS.n4839 VSS.n4840 0.147342
R9714 VSS.n4841 VSS.n4842 2.39784
R9715 VSS.n4842 VSS.n4843 0.147342
R9716 VSS.n4843 VSS.n4844 0.147342
R9717 VSS.n4844 VSS.t236 3.13212
R9718 VSS.n4822 VSS.n4817 4.5005
R9719 VSS.n4823 VSS.n4819 4.5005
R9720 VSS.n4824 VSS.n4820 4.5005
R9721 VSS.n4825 VSS.n4821 4.57324
R9722 VSS.n4815 VSS.n4817 0.147342
R9723 VSS.n4818 VSS.n4819 0.0732424
R9724 VSS.n4819 VSS.n4820 0.147342
R9725 VSS.n4826 VSS.n4822 0.0722544
R9726 VSS.n4827 VSS.n4823 4.5005
R9727 VSS.n4828 VSS.n4824 4.5005
R9728 VSS.n4829 VSS.n4825 4.5005
R9729 VSS.n4826 VSS.n4815 4.57426
R9730 VSS.n4822 VSS.n4823 0.147342
R9731 VSS.n4823 VSS.n4824 0.147342
R9732 VSS.n4824 VSS.n4825 0.147342
R9733 VSS.n4827 VSS.n4826 2.37296
R9734 VSS.n4828 VSS.n4827 0.127318
R9735 VSS.n4829 VSS.n4828 0.127318
R9736 VSS.t0 VSS.n4829 2.73618
R9737 VSS.n4802 VSS.n4807 4.5005
R9738 VSS.n4804 VSS.n4808 4.5005
R9739 VSS.n4805 VSS.n4809 4.5005
R9740 VSS.n4806 VSS.n4810 4.57324
R9741 VSS.n4802 VSS.n4800 0.147342
R9742 VSS.n4803 VSS.n4804 0.0732424
R9743 VSS.n4804 VSS.n4805 0.147342
R9744 VSS.n4807 VSS.n4811 0.0721009
R9745 VSS.n4812 VSS.n4808 4.5005
R9746 VSS.n4813 VSS.n4809 4.5005
R9747 VSS.n4814 VSS.n4810 4.5005
R9748 VSS.n4800 VSS.n4811 4.57442
R9749 VSS.n4807 VSS.n4808 0.147342
R9750 VSS.n4808 VSS.n4809 0.147342
R9751 VSS.n4809 VSS.n4810 0.147342
R9752 VSS.n4811 VSS.n4812 2.39784
R9753 VSS.n4812 VSS.n4813 0.147342
R9754 VSS.n4813 VSS.n4814 0.147342
R9755 VSS.n4814 VSS.t140 3.13212
R9756 VSS.n4787 VSS.n4792 4.5005
R9757 VSS.n4789 VSS.n4793 4.5005
R9758 VSS.n4790 VSS.n4794 4.5005
R9759 VSS.n4791 VSS.n4795 4.57324
R9760 VSS.n4787 VSS.n4785 0.147342
R9761 VSS.n4788 VSS.n4789 0.0732424
R9762 VSS.n4789 VSS.n4790 0.147342
R9763 VSS.n4792 VSS.n4796 0.0721009
R9764 VSS.n4797 VSS.n4793 4.5005
R9765 VSS.n4798 VSS.n4794 4.5005
R9766 VSS.n4799 VSS.n4795 4.5005
R9767 VSS.n4785 VSS.n4796 4.57442
R9768 VSS.n4792 VSS.n4793 0.147342
R9769 VSS.n4793 VSS.n4794 0.147342
R9770 VSS.n4794 VSS.n4795 0.147342
R9771 VSS.n4796 VSS.n4797 2.39784
R9772 VSS.n4797 VSS.n4798 0.147342
R9773 VSS.n4798 VSS.n4799 0.147342
R9774 VSS.n4799 VSS.t135 3.13212
R9775 VSS.n2370 VSS.n2371 0.0722544
R9776 VSS.n2372 VSS.n2373 4.5005
R9777 VSS.n2374 VSS.n2375 4.5005
R9778 VSS.n2376 VSS.n2377 4.5005
R9779 VSS.n2372 VSS.n2370 2.37296
R9780 VSS.n2374 VSS.n2372 0.127318
R9781 VSS.n2376 VSS.n2374 0.127318
R9782 VSS.t5 VSS.n2376 2.73618
R9783 VSS.n2371 VSS.n2378 4.5005
R9784 VSS.n2373 VSS.n2379 4.5005
R9785 VSS.n2375 VSS.n2380 4.5005
R9786 VSS.n2377 VSS.n2381 4.5005
R9787 VSS.n2383 VSS.n2370 4.647
R9788 VSS.n2371 VSS.n2373 0.147342
R9789 VSS.n2373 VSS.n2375 0.147342
R9790 VSS.n2375 VSS.n2377 0.147342
R9791 VSS.n2383 VSS.n2384 2.21488
R9792 VSS.n2378 VSS.n2383 0.0732424
R9793 VSS.n2382 VSS.n2384 2.21488
R9794 VSS.n2382 VSS.n2380 0.0732424
R9795 VSS.n2381 VSS.n2384 4.5005
R9796 VSS.n2378 VSS.n2379 0.147342
R9797 VSS.n2379 VSS.n2382 0.0732424
R9798 VSS.n2380 VSS.n2381 0.147342
R9799 VSS.n2385 VSS.n2386 4.5005
R9800 VSS.n2388 VSS.n2387 0.0732424
R9801 VSS.n2386 VSS.n2388 2.21488
R9802 VSS.n2391 VSS.n2390 0.0732424
R9803 VSS.n2386 VSS.n2391 2.21488
R9804 VSS.n2400 VSS.n2401 4.5005
R9805 VSS.n2403 VSS.n2402 0.0732424
R9806 VSS.n2401 VSS.n2403 2.21488
R9807 VSS.n2406 VSS.n2405 0.0732424
R9808 VSS.n2401 VSS.n2406 2.21488
R9809 VSS.n2415 VSS.n2416 4.5005
R9810 VSS.n2417 VSS.n2418 0.0732424
R9811 VSS.n2418 VSS.n2416 2.21488
R9812 VSS.n2420 VSS.n2421 0.0732424
R9813 VSS.n2421 VSS.n2416 2.21488
R9814 VSS.n2430 VSS.n2431 4.5005
R9815 VSS.n2433 VSS.n2432 0.0732424
R9816 VSS.n2431 VSS.n2433 2.21488
R9817 VSS.n2436 VSS.n2435 0.0732424
R9818 VSS.n2431 VSS.n2436 2.21488
R9819 VSS.n2445 VSS.n2446 4.5005
R9820 VSS.n2448 VSS.n2447 0.0732424
R9821 VSS.n2446 VSS.n2448 2.21488
R9822 VSS.n2451 VSS.n2450 0.0732424
R9823 VSS.n2446 VSS.n2451 2.21488
R9824 VSS.n2460 VSS.n2461 4.5005
R9825 VSS.n2463 VSS.n2462 0.0732424
R9826 VSS.n2461 VSS.n2463 2.21488
R9827 VSS.n2466 VSS.n2465 0.0732424
R9828 VSS.n2461 VSS.n2466 2.21488
R9829 VSS.n2475 VSS.n2476 4.5005
R9830 VSS.n2477 VSS.n2478 0.0732424
R9831 VSS.n2478 VSS.n2476 2.21488
R9832 VSS.n2480 VSS.n2481 0.0732424
R9833 VSS.n2481 VSS.n2476 2.21488
R9834 VSS.n2490 VSS.n2491 4.5005
R9835 VSS.n2493 VSS.n2492 0.0732424
R9836 VSS.n2491 VSS.n2493 2.21488
R9837 VSS.n2496 VSS.n2495 0.0732424
R9838 VSS.n2491 VSS.n2496 2.21488
R9839 VSS.n2505 VSS.n2506 4.5005
R9840 VSS.n2508 VSS.n2507 0.0732424
R9841 VSS.n2506 VSS.n2508 2.21488
R9842 VSS.n2511 VSS.n2510 0.0732424
R9843 VSS.n2506 VSS.n2511 2.21488
R9844 VSS.n2520 VSS.n2521 4.5005
R9845 VSS.n2523 VSS.n2522 0.0732424
R9846 VSS.n2521 VSS.n2523 2.21488
R9847 VSS.n2526 VSS.n2525 0.0732424
R9848 VSS.n2521 VSS.n2526 2.21488
R9849 VSS.n2535 VSS.n2536 4.5005
R9850 VSS.n2538 VSS.n2537 0.0732424
R9851 VSS.n2536 VSS.n2538 2.21488
R9852 VSS.n2541 VSS.n2540 0.0732424
R9853 VSS.n2536 VSS.n2541 2.21488
R9854 VSS.n2550 VSS.n2551 4.5005
R9855 VSS.n2553 VSS.n2552 0.0732424
R9856 VSS.n2551 VSS.n2553 2.21488
R9857 VSS.n2556 VSS.n2555 0.0732424
R9858 VSS.n2551 VSS.n2556 2.21488
R9859 VSS.n2565 VSS.n2566 4.5005
R9860 VSS.n2568 VSS.n2567 0.0732424
R9861 VSS.n2566 VSS.n2568 2.21488
R9862 VSS.n2571 VSS.n2570 0.0732424
R9863 VSS.n2566 VSS.n2571 2.21488
R9864 VSS.n2580 VSS.n2581 4.5005
R9865 VSS.n2582 VSS.n2583 0.0732424
R9866 VSS.n2583 VSS.n2581 2.21488
R9867 VSS.n2585 VSS.n2586 0.0732424
R9868 VSS.n2586 VSS.n2581 2.21488
R9869 VSS.n2595 VSS.n2596 4.5005
R9870 VSS.n2598 VSS.n2597 0.0732424
R9871 VSS.n2596 VSS.n2598 2.21488
R9872 VSS.n2601 VSS.n2600 0.0732424
R9873 VSS.n2596 VSS.n2601 2.21488
R9874 VSS.n2610 VSS.n2611 4.5005
R9875 VSS.n2613 VSS.n2612 0.0732424
R9876 VSS.n2611 VSS.n2613 2.21488
R9877 VSS.n2616 VSS.n2615 0.0732424
R9878 VSS.n2611 VSS.n2616 2.21488
R9879 VSS.n2625 VSS.n2626 4.5005
R9880 VSS.n2628 VSS.n2627 0.0732424
R9881 VSS.n2626 VSS.n2628 2.21488
R9882 VSS.n2631 VSS.n2630 0.0732424
R9883 VSS.n2626 VSS.n2631 2.21488
R9884 VSS.n2640 VSS.n2641 4.5005
R9885 VSS.n2642 VSS.n2643 0.0732424
R9886 VSS.n2643 VSS.n2641 2.21488
R9887 VSS.n2645 VSS.n2646 0.0732424
R9888 VSS.n2646 VSS.n2641 2.21488
R9889 VSS.n2655 VSS.n2656 4.5005
R9890 VSS.n2658 VSS.n2657 0.0732424
R9891 VSS.n2656 VSS.n2658 2.21488
R9892 VSS.n2661 VSS.n2660 0.0732424
R9893 VSS.n2656 VSS.n2661 2.21488
R9894 VSS.n2670 VSS.n2671 4.5005
R9895 VSS.n2673 VSS.n2672 0.0732424
R9896 VSS.n2671 VSS.n2673 2.21488
R9897 VSS.n2676 VSS.n2675 0.0732424
R9898 VSS.n2671 VSS.n2676 2.21488
R9899 VSS.n2685 VSS.n2686 4.5005
R9900 VSS.n2688 VSS.n2687 0.0732424
R9901 VSS.n2686 VSS.n2688 2.21488
R9902 VSS.n2691 VSS.n2690 0.0732424
R9903 VSS.n2686 VSS.n2691 2.21488
R9904 VSS.n2700 VSS.n2701 4.5005
R9905 VSS.n2703 VSS.n2702 0.0732424
R9906 VSS.n2701 VSS.n2703 2.21488
R9907 VSS.n2706 VSS.n2705 0.0732424
R9908 VSS.n2701 VSS.n2706 2.21488
R9909 VSS.n2715 VSS.n2716 4.5005
R9910 VSS.n2717 VSS.n2718 0.0732424
R9911 VSS.n2718 VSS.n2716 2.21488
R9912 VSS.n2720 VSS.n2721 0.0732424
R9913 VSS.n2721 VSS.n2716 2.21488
R9914 VSS.n2730 VSS.n2731 4.5005
R9915 VSS.n2733 VSS.n2732 0.0732424
R9916 VSS.n2731 VSS.n2733 2.21488
R9917 VSS.n2736 VSS.n2735 0.0732424
R9918 VSS.n2731 VSS.n2736 2.21488
R9919 VSS.n2745 VSS.n2746 4.5005
R9920 VSS.n2748 VSS.n2747 0.0732424
R9921 VSS.n2746 VSS.n2748 2.21488
R9922 VSS.n2751 VSS.n2750 0.0732424
R9923 VSS.n2746 VSS.n2751 2.21488
R9924 VSS.n2760 VSS.n2761 4.5005
R9925 VSS.n2763 VSS.n2762 0.0732424
R9926 VSS.n2761 VSS.n2763 2.21488
R9927 VSS.n2766 VSS.n2765 0.0732424
R9928 VSS.n2761 VSS.n2766 2.21488
R9929 VSS.n2775 VSS.n2776 4.5005
R9930 VSS.n2777 VSS.n2778 0.0732424
R9931 VSS.n2778 VSS.n2776 2.21488
R9932 VSS.n2780 VSS.n2781 0.0732424
R9933 VSS.n2781 VSS.n2776 2.21488
R9934 VSS.n2790 VSS.n2791 4.5005
R9935 VSS.n2793 VSS.n2792 0.0732424
R9936 VSS.n2791 VSS.n2793 2.21488
R9937 VSS.n2796 VSS.n2795 0.0732424
R9938 VSS.n2791 VSS.n2796 2.21488
R9939 VSS.n2805 VSS.n2806 4.5005
R9940 VSS.n2808 VSS.n2807 0.0732424
R9941 VSS.n2806 VSS.n2808 2.21488
R9942 VSS.n2811 VSS.n2810 0.0732424
R9943 VSS.n2806 VSS.n2811 2.21488
R9944 VSS.n2820 VSS.n2821 4.5005
R9945 VSS.n2823 VSS.n2822 0.0732424
R9946 VSS.n2821 VSS.n2823 2.21488
R9947 VSS.n2826 VSS.n2825 0.0732424
R9948 VSS.n2821 VSS.n2826 2.21488
R9949 VSS.n2835 VSS.n2836 4.5005
R9950 VSS.n2838 VSS.n2837 0.0732424
R9951 VSS.n2836 VSS.n2838 2.21488
R9952 VSS.n2841 VSS.n2840 0.0732424
R9953 VSS.n2836 VSS.n2841 2.21488
R9954 VSS.n2850 VSS.n2851 4.5005
R9955 VSS.n2853 VSS.n2852 0.0732424
R9956 VSS.n2851 VSS.n2853 2.21488
R9957 VSS.n2856 VSS.n2855 0.0732424
R9958 VSS.n2851 VSS.n2856 2.21488
R9959 VSS.n2865 VSS.n2866 4.5005
R9960 VSS.n2868 VSS.n2867 0.0732424
R9961 VSS.n2866 VSS.n2868 2.21488
R9962 VSS.n2871 VSS.n2870 0.0732424
R9963 VSS.n2866 VSS.n2871 2.21488
R9964 VSS.n2880 VSS.n2881 4.5005
R9965 VSS.n2882 VSS.n2883 0.0732424
R9966 VSS.n2883 VSS.n2881 2.21488
R9967 VSS.n2885 VSS.n2886 0.0732424
R9968 VSS.n2886 VSS.n2881 2.21488
R9969 VSS.n2895 VSS.n2896 4.5005
R9970 VSS.n2898 VSS.n2897 0.0732424
R9971 VSS.n2896 VSS.n2898 2.21488
R9972 VSS.n2901 VSS.n2900 0.0732424
R9973 VSS.n2896 VSS.n2901 2.21488
R9974 VSS.n2910 VSS.n2911 4.5005
R9975 VSS.n2913 VSS.n2912 0.0732424
R9976 VSS.n2911 VSS.n2913 2.21488
R9977 VSS.n2916 VSS.n2915 0.0732424
R9978 VSS.n2911 VSS.n2916 2.21488
R9979 VSS.n2925 VSS.n2926 4.5005
R9980 VSS.n2928 VSS.n2927 0.0732424
R9981 VSS.n2926 VSS.n2928 2.21488
R9982 VSS.n2931 VSS.n2930 0.0732424
R9983 VSS.n2926 VSS.n2931 2.21488
R9984 VSS.n2940 VSS.n2941 4.5005
R9985 VSS.n2942 VSS.n2943 0.0732424
R9986 VSS.n2943 VSS.n2941 2.21488
R9987 VSS.n2945 VSS.n2946 0.0732424
R9988 VSS.n2946 VSS.n2941 2.21488
R9989 VSS.n2955 VSS.n2956 4.5005
R9990 VSS.n2958 VSS.n2957 0.0732424
R9991 VSS.n2956 VSS.n2958 2.21488
R9992 VSS.n2961 VSS.n2960 0.0732424
R9993 VSS.n2956 VSS.n2961 2.21488
R9994 VSS.n2970 VSS.n2971 4.5005
R9995 VSS.n2973 VSS.n2972 0.0732424
R9996 VSS.n2971 VSS.n2973 2.21488
R9997 VSS.n2976 VSS.n2975 0.0732424
R9998 VSS.n2971 VSS.n2976 2.21488
R9999 VSS.n2985 VSS.n2986 4.5005
R10000 VSS.n2988 VSS.n2987 0.0732424
R10001 VSS.n2986 VSS.n2988 2.21488
R10002 VSS.n2991 VSS.n2990 0.0732424
R10003 VSS.n2986 VSS.n2991 2.21488
R10004 VSS.n3000 VSS.n3001 4.5005
R10005 VSS.n3003 VSS.n3002 0.0732424
R10006 VSS.n3001 VSS.n3003 2.21488
R10007 VSS.n3006 VSS.n3005 0.0732424
R10008 VSS.n3001 VSS.n3006 2.21488
R10009 VSS.n3015 VSS.n3016 4.5005
R10010 VSS.n3017 VSS.n3018 0.0732424
R10011 VSS.n3018 VSS.n3016 2.21488
R10012 VSS.n3020 VSS.n3021 0.0732424
R10013 VSS.n3021 VSS.n3016 2.21488
R10014 VSS.n3030 VSS.n3031 4.5005
R10015 VSS.n3033 VSS.n3032 0.0732424
R10016 VSS.n3031 VSS.n3033 2.21488
R10017 VSS.n3036 VSS.n3035 0.0732424
R10018 VSS.n3031 VSS.n3036 2.21488
R10019 VSS.n3045 VSS.n3046 4.5005
R10020 VSS.n3048 VSS.n3047 0.0732424
R10021 VSS.n3046 VSS.n3048 2.21488
R10022 VSS.n3051 VSS.n3050 0.0732424
R10023 VSS.n3046 VSS.n3051 2.21488
R10024 VSS.n3060 VSS.n3061 4.5005
R10025 VSS.n3063 VSS.n3062 0.0732424
R10026 VSS.n3061 VSS.n3063 2.21488
R10027 VSS.n3066 VSS.n3065 0.0732424
R10028 VSS.n3061 VSS.n3066 2.21488
R10029 VSS.n3075 VSS.n3076 4.5005
R10030 VSS.n3077 VSS.n3078 0.0732424
R10031 VSS.n3078 VSS.n3076 2.21488
R10032 VSS.n3080 VSS.n3081 0.0732424
R10033 VSS.n3081 VSS.n3076 2.21488
R10034 VSS.n3090 VSS.n3091 4.5005
R10035 VSS.n3093 VSS.n3092 0.0732424
R10036 VSS.n3091 VSS.n3093 2.21488
R10037 VSS.n3096 VSS.n3095 0.0732424
R10038 VSS.n3091 VSS.n3096 2.21488
R10039 VSS.n3105 VSS.n3106 4.5005
R10040 VSS.n3108 VSS.n3107 0.0732424
R10041 VSS.n3106 VSS.n3108 2.21488
R10042 VSS.n3111 VSS.n3110 0.0732424
R10043 VSS.n3106 VSS.n3111 2.21488
R10044 VSS.n3120 VSS.n3121 4.5005
R10045 VSS.n3123 VSS.n3122 0.0732424
R10046 VSS.n3121 VSS.n3123 2.21488
R10047 VSS.n3126 VSS.n3125 0.0732424
R10048 VSS.n3121 VSS.n3126 2.21488
R10049 VSS.n3135 VSS.n3136 4.5005
R10050 VSS.n3138 VSS.n3137 0.0732424
R10051 VSS.n3136 VSS.n3138 2.21488
R10052 VSS.n3141 VSS.n3140 0.0732424
R10053 VSS.n3136 VSS.n3141 2.21488
R10054 VSS.n3150 VSS.n3151 4.5005
R10055 VSS.n3153 VSS.n3152 0.0732424
R10056 VSS.n3151 VSS.n3153 2.21488
R10057 VSS.n3156 VSS.n3155 0.0732424
R10058 VSS.n3151 VSS.n3156 2.21488
R10059 VSS.n3165 VSS.n3166 4.5005
R10060 VSS.n3168 VSS.n3167 0.0732424
R10061 VSS.n3166 VSS.n3168 2.21488
R10062 VSS.n3171 VSS.n3170 0.0732424
R10063 VSS.n3166 VSS.n3171 2.21488
R10064 VSS.n3180 VSS.n3181 4.5005
R10065 VSS.n3182 VSS.n3183 0.0732424
R10066 VSS.n3183 VSS.n3181 2.21488
R10067 VSS.n3185 VSS.n3186 0.0732424
R10068 VSS.n3186 VSS.n3181 2.21488
R10069 VSS.n3195 VSS.n3196 4.5005
R10070 VSS.n3198 VSS.n3197 0.0732424
R10071 VSS.n3196 VSS.n3198 2.21488
R10072 VSS.n3201 VSS.n3200 0.0732424
R10073 VSS.n3196 VSS.n3201 2.21488
R10074 VSS.n3210 VSS.n3211 4.5005
R10075 VSS.n3213 VSS.n3212 0.0732424
R10076 VSS.n3211 VSS.n3213 2.21488
R10077 VSS.n3216 VSS.n3215 0.0732424
R10078 VSS.n3211 VSS.n3216 2.21488
R10079 VSS.n3225 VSS.n3226 4.5005
R10080 VSS.n3228 VSS.n3227 0.0732424
R10081 VSS.n3226 VSS.n3228 2.21488
R10082 VSS.n3231 VSS.n3230 0.0732424
R10083 VSS.n3226 VSS.n3231 2.21488
R10084 VSS.n3240 VSS.n3241 4.5005
R10085 VSS.n3242 VSS.n3243 0.0732424
R10086 VSS.n3243 VSS.n3241 2.21488
R10087 VSS.n3245 VSS.n3246 0.0732424
R10088 VSS.n3246 VSS.n3241 2.21488
R10089 VSS.n3255 VSS.n3256 4.5005
R10090 VSS.n3258 VSS.n3257 0.0732424
R10091 VSS.n3256 VSS.n3258 2.21488
R10092 VSS.n3261 VSS.n3260 0.0732424
R10093 VSS.n3256 VSS.n3261 2.21488
R10094 VSS.n3270 VSS.n3271 4.5005
R10095 VSS.n3273 VSS.n3272 0.0732424
R10096 VSS.n3271 VSS.n3273 2.21488
R10097 VSS.n3276 VSS.n3275 0.0732424
R10098 VSS.n3271 VSS.n3276 2.21488
R10099 VSS.n3285 VSS.n3286 4.5005
R10100 VSS.n3288 VSS.n3287 0.0732424
R10101 VSS.n3286 VSS.n3288 2.21488
R10102 VSS.n3291 VSS.n3290 0.0732424
R10103 VSS.n3286 VSS.n3291 2.21488
R10104 VSS.n3300 VSS.n3301 4.5005
R10105 VSS.n3303 VSS.n3302 0.0732424
R10106 VSS.n3301 VSS.n3303 2.21488
R10107 VSS.n3306 VSS.n3305 0.0732424
R10108 VSS.n3301 VSS.n3306 2.21488
R10109 VSS.n3315 VSS.n3316 4.5005
R10110 VSS.n3317 VSS.n3318 0.0732424
R10111 VSS.n3318 VSS.n3316 2.21488
R10112 VSS.n3320 VSS.n3321 0.0732424
R10113 VSS.n3321 VSS.n3316 2.21488
R10114 VSS.n3330 VSS.n3331 4.5005
R10115 VSS.n3333 VSS.n3332 0.0732424
R10116 VSS.n3331 VSS.n3333 2.21488
R10117 VSS.n3336 VSS.n3335 0.0732424
R10118 VSS.n3331 VSS.n3336 2.21488
R10119 VSS.n3345 VSS.n3346 4.5005
R10120 VSS.n3348 VSS.n3347 0.0732424
R10121 VSS.n3346 VSS.n3348 2.21488
R10122 VSS.n3351 VSS.n3350 0.0732424
R10123 VSS.n3346 VSS.n3351 2.21488
R10124 VSS.n3360 VSS.n3361 4.5005
R10125 VSS.n3363 VSS.n3362 0.0732424
R10126 VSS.n3361 VSS.n3363 2.21488
R10127 VSS.n3366 VSS.n3365 0.0732424
R10128 VSS.n3361 VSS.n3366 2.21488
R10129 VSS.n3375 VSS.n3376 4.5005
R10130 VSS.n3377 VSS.n3378 0.0732424
R10131 VSS.n3378 VSS.n3376 2.21488
R10132 VSS.n3380 VSS.n3381 0.0732424
R10133 VSS.n3381 VSS.n3376 2.21488
R10134 VSS.n3390 VSS.n3391 4.5005
R10135 VSS.n3393 VSS.n3392 0.0732424
R10136 VSS.n3391 VSS.n3393 2.21488
R10137 VSS.n3396 VSS.n3395 0.0732424
R10138 VSS.n3391 VSS.n3396 2.21488
R10139 VSS.n3405 VSS.n3406 4.5005
R10140 VSS.n3408 VSS.n3407 0.0732424
R10141 VSS.n3406 VSS.n3408 2.21488
R10142 VSS.n3411 VSS.n3410 0.0732424
R10143 VSS.n3406 VSS.n3411 2.21488
R10144 VSS.n3420 VSS.n3421 4.5005
R10145 VSS.n3423 VSS.n3422 0.0732424
R10146 VSS.n3421 VSS.n3423 2.21488
R10147 VSS.n3426 VSS.n3425 0.0732424
R10148 VSS.n3421 VSS.n3426 2.21488
R10149 VSS.n3435 VSS.n3436 4.5005
R10150 VSS.n3438 VSS.n3437 0.0732424
R10151 VSS.n3436 VSS.n3438 2.21488
R10152 VSS.n3441 VSS.n3440 0.0732424
R10153 VSS.n3436 VSS.n3441 2.21488
R10154 VSS.n3450 VSS.n3451 4.5005
R10155 VSS.n3453 VSS.n3452 0.0732424
R10156 VSS.n3451 VSS.n3453 2.21488
R10157 VSS.n3456 VSS.n3455 0.0732424
R10158 VSS.n3451 VSS.n3456 2.21488
R10159 VSS.n3465 VSS.n3466 4.5005
R10160 VSS.n3468 VSS.n3467 0.0732424
R10161 VSS.n3466 VSS.n3468 2.21488
R10162 VSS.n3471 VSS.n3470 0.0732424
R10163 VSS.n3466 VSS.n3471 2.21488
R10164 VSS.n3480 VSS.n3481 4.5005
R10165 VSS.n3482 VSS.n3483 0.0732424
R10166 VSS.n3483 VSS.n3481 2.21488
R10167 VSS.n3485 VSS.n3486 0.0732424
R10168 VSS.n3486 VSS.n3481 2.21488
R10169 VSS.n3495 VSS.n3496 4.5005
R10170 VSS.n3498 VSS.n3497 0.0732424
R10171 VSS.n3496 VSS.n3498 2.21488
R10172 VSS.n3501 VSS.n3500 0.0732424
R10173 VSS.n3496 VSS.n3501 2.21488
R10174 VSS.n3510 VSS.n3511 4.5005
R10175 VSS.n3513 VSS.n3512 0.0732424
R10176 VSS.n3511 VSS.n3513 2.21488
R10177 VSS.n3516 VSS.n3515 0.0732424
R10178 VSS.n3511 VSS.n3516 2.21488
R10179 VSS.n3525 VSS.n3526 4.5005
R10180 VSS.n3528 VSS.n3527 0.0732424
R10181 VSS.n3526 VSS.n3528 2.21488
R10182 VSS.n3531 VSS.n3530 0.0732424
R10183 VSS.n3526 VSS.n3531 2.21488
R10184 VSS.n3540 VSS.n3541 4.5005
R10185 VSS.n3542 VSS.n3543 0.0732424
R10186 VSS.n3543 VSS.n3541 2.21488
R10187 VSS.n3545 VSS.n3546 0.0732424
R10188 VSS.n3546 VSS.n3541 2.21488
R10189 VSS.n3555 VSS.n3556 4.5005
R10190 VSS.n3558 VSS.n3557 0.0732424
R10191 VSS.n3556 VSS.n3558 2.21488
R10192 VSS.n3561 VSS.n3560 0.0732424
R10193 VSS.n3556 VSS.n3561 2.21488
R10194 VSS.n3570 VSS.n3571 4.5005
R10195 VSS.n3573 VSS.n3572 0.0732424
R10196 VSS.n3571 VSS.n3573 2.21488
R10197 VSS.n3576 VSS.n3575 0.0732424
R10198 VSS.n3571 VSS.n3576 2.21488
R10199 VSS.n3585 VSS.n3586 4.5005
R10200 VSS.n3588 VSS.n3587 0.0732424
R10201 VSS.n3586 VSS.n3588 2.21488
R10202 VSS.n3591 VSS.n3590 0.0732424
R10203 VSS.n3586 VSS.n3591 2.21488
R10204 VSS.n3600 VSS.n3601 4.5005
R10205 VSS.n3603 VSS.n3602 0.0732424
R10206 VSS.n3601 VSS.n3603 2.21488
R10207 VSS.n3606 VSS.n3605 0.0732424
R10208 VSS.n3601 VSS.n3606 2.21488
R10209 VSS.n3615 VSS.n3616 4.5005
R10210 VSS.n3617 VSS.n3618 0.0732424
R10211 VSS.n3618 VSS.n3616 2.21488
R10212 VSS.n3620 VSS.n3621 0.0732424
R10213 VSS.n3621 VSS.n3616 2.21488
R10214 VSS.n3630 VSS.n3631 4.5005
R10215 VSS.n3633 VSS.n3632 0.0732424
R10216 VSS.n3631 VSS.n3633 2.21488
R10217 VSS.n3636 VSS.n3635 0.0732424
R10218 VSS.n3631 VSS.n3636 2.21488
R10219 VSS.n3645 VSS.n3646 4.5005
R10220 VSS.n3648 VSS.n3647 0.0732424
R10221 VSS.n3646 VSS.n3648 2.21488
R10222 VSS.n3651 VSS.n3650 0.0732424
R10223 VSS.n3646 VSS.n3651 2.21488
R10224 VSS.n3660 VSS.n3661 4.5005
R10225 VSS.n3663 VSS.n3662 0.0732424
R10226 VSS.n3661 VSS.n3663 2.21488
R10227 VSS.n3666 VSS.n3665 0.0732424
R10228 VSS.n3661 VSS.n3666 2.21488
R10229 VSS.n3675 VSS.n3676 4.5005
R10230 VSS.n3677 VSS.n3678 0.0732424
R10231 VSS.n3678 VSS.n3676 2.21488
R10232 VSS.n3680 VSS.n3681 0.0732424
R10233 VSS.n3681 VSS.n3676 2.21488
R10234 VSS.n3690 VSS.n3691 4.5005
R10235 VSS.n3693 VSS.n3692 0.0732424
R10236 VSS.n3691 VSS.n3693 2.21488
R10237 VSS.n3696 VSS.n3695 0.0732424
R10238 VSS.n3691 VSS.n3696 2.21488
R10239 VSS.n3705 VSS.n3706 4.5005
R10240 VSS.n3708 VSS.n3707 0.0732424
R10241 VSS.n3706 VSS.n3708 2.21488
R10242 VSS.n3711 VSS.n3710 0.0732424
R10243 VSS.n3706 VSS.n3711 2.21488
R10244 VSS.n3720 VSS.n3721 4.5005
R10245 VSS.n3723 VSS.n3722 0.0732424
R10246 VSS.n3721 VSS.n3723 2.21488
R10247 VSS.n3726 VSS.n3725 0.0732424
R10248 VSS.n3721 VSS.n3726 2.21488
R10249 VSS.n3735 VSS.n3736 4.5005
R10250 VSS.n3738 VSS.n3737 0.0732424
R10251 VSS.n3736 VSS.n3738 2.21488
R10252 VSS.n3741 VSS.n3740 0.0732424
R10253 VSS.n3736 VSS.n3741 2.21488
R10254 VSS.n3750 VSS.n3751 4.5005
R10255 VSS.n3753 VSS.n3752 0.0732424
R10256 VSS.n3751 VSS.n3753 2.21488
R10257 VSS.n3756 VSS.n3755 0.0732424
R10258 VSS.n3751 VSS.n3756 2.21488
R10259 VSS.n3765 VSS.n3766 4.5005
R10260 VSS.n3768 VSS.n3767 0.0732424
R10261 VSS.n3766 VSS.n3768 2.21488
R10262 VSS.n3771 VSS.n3770 0.0732424
R10263 VSS.n3766 VSS.n3771 2.21488
R10264 VSS.n3780 VSS.n3781 4.5005
R10265 VSS.n3782 VSS.n3783 0.0732424
R10266 VSS.n3783 VSS.n3781 2.21488
R10267 VSS.n3785 VSS.n3786 0.0732424
R10268 VSS.n3786 VSS.n3781 2.21488
R10269 VSS.n3795 VSS.n3796 4.5005
R10270 VSS.n3798 VSS.n3797 0.0732424
R10271 VSS.n3796 VSS.n3798 2.21488
R10272 VSS.n3801 VSS.n3800 0.0732424
R10273 VSS.n3796 VSS.n3801 2.21488
R10274 VSS.n3810 VSS.n3811 4.5005
R10275 VSS.n3813 VSS.n3812 0.0732424
R10276 VSS.n3811 VSS.n3813 2.21488
R10277 VSS.n3816 VSS.n3815 0.0732424
R10278 VSS.n3811 VSS.n3816 2.21488
R10279 VSS.n3825 VSS.n3826 4.5005
R10280 VSS.n3828 VSS.n3827 0.0732424
R10281 VSS.n3826 VSS.n3828 2.21488
R10282 VSS.n3831 VSS.n3830 0.0732424
R10283 VSS.n3826 VSS.n3831 2.21488
R10284 VSS.n3840 VSS.n3841 4.5005
R10285 VSS.n3842 VSS.n3843 0.0732424
R10286 VSS.n3843 VSS.n3841 2.21488
R10287 VSS.n3845 VSS.n3846 0.0732424
R10288 VSS.n3846 VSS.n3841 2.21488
R10289 VSS.n3855 VSS.n3856 4.5005
R10290 VSS.n3858 VSS.n3857 0.0732424
R10291 VSS.n3856 VSS.n3858 2.21488
R10292 VSS.n3861 VSS.n3860 0.0732424
R10293 VSS.n3856 VSS.n3861 2.21488
R10294 VSS.n3870 VSS.n3871 4.5005
R10295 VSS.n3873 VSS.n3872 0.0732424
R10296 VSS.n3871 VSS.n3873 2.21488
R10297 VSS.n3876 VSS.n3875 0.0732424
R10298 VSS.n3871 VSS.n3876 2.21488
R10299 VSS.n3885 VSS.n3886 4.5005
R10300 VSS.n3888 VSS.n3887 0.0732424
R10301 VSS.n3886 VSS.n3888 2.21488
R10302 VSS.n3891 VSS.n3890 0.0732424
R10303 VSS.n3886 VSS.n3891 2.21488
R10304 VSS.n3900 VSS.n3901 4.5005
R10305 VSS.n3903 VSS.n3902 0.0732424
R10306 VSS.n3901 VSS.n3903 2.21488
R10307 VSS.n3906 VSS.n3905 0.0732424
R10308 VSS.n3901 VSS.n3906 2.21488
R10309 VSS.n3915 VSS.n3916 4.5005
R10310 VSS.n3917 VSS.n3918 0.0732424
R10311 VSS.n3918 VSS.n3916 2.21488
R10312 VSS.n3920 VSS.n3921 0.0732424
R10313 VSS.n3921 VSS.n3916 2.21488
R10314 VSS.n3930 VSS.n3931 4.5005
R10315 VSS.n3933 VSS.n3932 0.0732424
R10316 VSS.n3931 VSS.n3933 2.21488
R10317 VSS.n3936 VSS.n3935 0.0732424
R10318 VSS.n3931 VSS.n3936 2.21488
R10319 VSS.n3945 VSS.n3946 4.5005
R10320 VSS.n3948 VSS.n3947 0.0732424
R10321 VSS.n3946 VSS.n3948 2.21488
R10322 VSS.n3951 VSS.n3950 0.0732424
R10323 VSS.n3946 VSS.n3951 2.21488
R10324 VSS.n3960 VSS.n3961 4.5005
R10325 VSS.n3963 VSS.n3962 0.0732424
R10326 VSS.n3961 VSS.n3963 2.21488
R10327 VSS.n3966 VSS.n3965 0.0732424
R10328 VSS.n3961 VSS.n3966 2.21488
R10329 VSS.n3975 VSS.n3976 4.5005
R10330 VSS.n3977 VSS.n3978 0.0732424
R10331 VSS.n3978 VSS.n3976 2.21488
R10332 VSS.n3980 VSS.n3981 0.0732424
R10333 VSS.n3981 VSS.n3976 2.21488
R10334 VSS.n3990 VSS.n3991 4.5005
R10335 VSS.n3993 VSS.n3992 0.0732424
R10336 VSS.n3991 VSS.n3993 2.21488
R10337 VSS.n3996 VSS.n3995 0.0732424
R10338 VSS.n3991 VSS.n3996 2.21488
R10339 VSS.n4005 VSS.n4006 4.5005
R10340 VSS.n4008 VSS.n4007 0.0732424
R10341 VSS.n4006 VSS.n4008 2.21488
R10342 VSS.n4011 VSS.n4010 0.0732424
R10343 VSS.n4006 VSS.n4011 2.21488
R10344 VSS.n4020 VSS.n4021 4.5005
R10345 VSS.n4023 VSS.n4022 0.0732424
R10346 VSS.n4021 VSS.n4023 2.21488
R10347 VSS.n4026 VSS.n4025 0.0732424
R10348 VSS.n4021 VSS.n4026 2.21488
R10349 VSS.n4035 VSS.n4036 4.5005
R10350 VSS.n4038 VSS.n4037 0.0732424
R10351 VSS.n4036 VSS.n4038 2.21488
R10352 VSS.n4041 VSS.n4040 0.0732424
R10353 VSS.n4036 VSS.n4041 2.21488
R10354 VSS.n4050 VSS.n4051 4.5005
R10355 VSS.n4053 VSS.n4052 0.0732424
R10356 VSS.n4051 VSS.n4053 2.21488
R10357 VSS.n4056 VSS.n4055 0.0732424
R10358 VSS.n4051 VSS.n4056 2.21488
R10359 VSS.n4065 VSS.n4066 4.5005
R10360 VSS.n4068 VSS.n4067 0.0732424
R10361 VSS.n4066 VSS.n4068 2.21488
R10362 VSS.n4071 VSS.n4070 0.0732424
R10363 VSS.n4066 VSS.n4071 2.21488
R10364 VSS.n4080 VSS.n4081 4.5005
R10365 VSS.n4082 VSS.n4083 0.0732424
R10366 VSS.n4083 VSS.n4081 2.21488
R10367 VSS.n4085 VSS.n4086 0.0732424
R10368 VSS.n4086 VSS.n4081 2.21488
R10369 VSS.n4095 VSS.n4096 4.5005
R10370 VSS.n4098 VSS.n4097 0.0732424
R10371 VSS.n4096 VSS.n4098 2.21488
R10372 VSS.n4101 VSS.n4100 0.0732424
R10373 VSS.n4096 VSS.n4101 2.21488
R10374 VSS.n4110 VSS.n4111 4.5005
R10375 VSS.n4113 VSS.n4112 0.0732424
R10376 VSS.n4111 VSS.n4113 2.21488
R10377 VSS.n4116 VSS.n4115 0.0732424
R10378 VSS.n4111 VSS.n4116 2.21488
R10379 VSS.n4125 VSS.n4126 4.5005
R10380 VSS.n4128 VSS.n4127 0.0732424
R10381 VSS.n4126 VSS.n4128 2.21488
R10382 VSS.n4131 VSS.n4130 0.0732424
R10383 VSS.n4126 VSS.n4131 2.21488
R10384 VSS.n4140 VSS.n4141 4.5005
R10385 VSS.n4142 VSS.n4143 0.0732424
R10386 VSS.n4143 VSS.n4141 2.21488
R10387 VSS.n4145 VSS.n4146 0.0732424
R10388 VSS.n4146 VSS.n4141 2.21488
R10389 VSS.n4155 VSS.n4156 4.5005
R10390 VSS.n4158 VSS.n4157 0.0732424
R10391 VSS.n4156 VSS.n4158 2.21488
R10392 VSS.n4161 VSS.n4160 0.0732424
R10393 VSS.n4156 VSS.n4161 2.21488
R10394 VSS.n4170 VSS.n4171 4.5005
R10395 VSS.n4173 VSS.n4172 0.0732424
R10396 VSS.n4171 VSS.n4173 2.21488
R10397 VSS.n4176 VSS.n4175 0.0732424
R10398 VSS.n4171 VSS.n4176 2.21488
R10399 VSS.n4185 VSS.n4186 4.5005
R10400 VSS.n4188 VSS.n4187 0.0732424
R10401 VSS.n4186 VSS.n4188 2.21488
R10402 VSS.n4191 VSS.n4190 0.0732424
R10403 VSS.n4186 VSS.n4191 2.21488
R10404 VSS.n4200 VSS.n4201 4.5005
R10405 VSS.n4203 VSS.n4202 0.0732424
R10406 VSS.n4201 VSS.n4203 2.21488
R10407 VSS.n4206 VSS.n4205 0.0732424
R10408 VSS.n4201 VSS.n4206 2.21488
R10409 VSS.n4215 VSS.n4216 4.5005
R10410 VSS.n4217 VSS.n4218 0.0732424
R10411 VSS.n4218 VSS.n4216 2.21488
R10412 VSS.n4220 VSS.n4221 0.0732424
R10413 VSS.n4221 VSS.n4216 2.21488
R10414 VSS.n4230 VSS.n4231 4.5005
R10415 VSS.n4233 VSS.n4232 0.0732424
R10416 VSS.n4231 VSS.n4233 2.21488
R10417 VSS.n4236 VSS.n4235 0.0732424
R10418 VSS.n4231 VSS.n4236 2.21488
R10419 VSS.n4245 VSS.n4246 4.5005
R10420 VSS.n4248 VSS.n4247 0.0732424
R10421 VSS.n4246 VSS.n4248 2.21488
R10422 VSS.n4251 VSS.n4250 0.0732424
R10423 VSS.n4246 VSS.n4251 2.21488
R10424 VSS.n4260 VSS.n4261 4.5005
R10425 VSS.n4263 VSS.n4262 0.0732424
R10426 VSS.n4261 VSS.n4263 2.21488
R10427 VSS.n4266 VSS.n4265 0.0732424
R10428 VSS.n4261 VSS.n4266 2.21488
R10429 VSS.n4275 VSS.n4276 4.5005
R10430 VSS.n4277 VSS.n4278 0.0732424
R10431 VSS.n4278 VSS.n4276 2.21488
R10432 VSS.n4280 VSS.n4281 0.0732424
R10433 VSS.n4281 VSS.n4276 2.21488
R10434 VSS.n4290 VSS.n4291 4.5005
R10435 VSS.n4293 VSS.n4292 0.0732424
R10436 VSS.n4291 VSS.n4293 2.21488
R10437 VSS.n4296 VSS.n4295 0.0732424
R10438 VSS.n4291 VSS.n4296 2.21488
R10439 VSS.n4305 VSS.n4306 4.5005
R10440 VSS.n4308 VSS.n4307 0.0732424
R10441 VSS.n4306 VSS.n4308 2.21488
R10442 VSS.n4311 VSS.n4310 0.0732424
R10443 VSS.n4306 VSS.n4311 2.21488
R10444 VSS.n4320 VSS.n4321 4.5005
R10445 VSS.n4323 VSS.n4322 0.0732424
R10446 VSS.n4321 VSS.n4323 2.21488
R10447 VSS.n4326 VSS.n4325 0.0732424
R10448 VSS.n4321 VSS.n4326 2.21488
R10449 VSS.n4335 VSS.n4336 4.5005
R10450 VSS.n4338 VSS.n4337 0.0732424
R10451 VSS.n4336 VSS.n4338 2.21488
R10452 VSS.n4341 VSS.n4340 0.0732424
R10453 VSS.n4336 VSS.n4341 2.21488
R10454 VSS.n4350 VSS.n4351 4.5005
R10455 VSS.n4353 VSS.n4352 0.0732424
R10456 VSS.n4351 VSS.n4353 2.21488
R10457 VSS.n4356 VSS.n4355 0.0732424
R10458 VSS.n4351 VSS.n4356 2.21488
R10459 VSS.n4365 VSS.n4366 4.5005
R10460 VSS.n4368 VSS.n4367 0.0732424
R10461 VSS.n4366 VSS.n4368 2.21488
R10462 VSS.n4371 VSS.n4370 0.0732424
R10463 VSS.n4366 VSS.n4371 2.21488
R10464 VSS.n4380 VSS.n4381 4.5005
R10465 VSS.n4382 VSS.n4383 0.0732424
R10466 VSS.n4383 VSS.n4381 2.21488
R10467 VSS.n4385 VSS.n4386 0.0732424
R10468 VSS.n4386 VSS.n4381 2.21488
R10469 VSS.n4395 VSS.n4396 4.5005
R10470 VSS.n4398 VSS.n4397 0.0732424
R10471 VSS.n4396 VSS.n4398 2.21488
R10472 VSS.n4401 VSS.n4400 0.0732424
R10473 VSS.n4396 VSS.n4401 2.21488
R10474 VSS.n4410 VSS.n4411 4.5005
R10475 VSS.n4413 VSS.n4412 0.0732424
R10476 VSS.n4411 VSS.n4413 2.21488
R10477 VSS.n4416 VSS.n4415 0.0732424
R10478 VSS.n4411 VSS.n4416 2.21488
R10479 VSS.n4425 VSS.n4426 4.5005
R10480 VSS.n4428 VSS.n4427 0.0732424
R10481 VSS.n4426 VSS.n4428 2.21488
R10482 VSS.n4431 VSS.n4430 0.0732424
R10483 VSS.n4426 VSS.n4431 2.21488
R10484 VSS.n4440 VSS.n4441 4.5005
R10485 VSS.n4442 VSS.n4443 0.0732424
R10486 VSS.n4443 VSS.n4441 2.21488
R10487 VSS.n4445 VSS.n4446 0.0732424
R10488 VSS.n4446 VSS.n4441 2.21488
R10489 VSS.n4455 VSS.n4456 4.5005
R10490 VSS.n4458 VSS.n4457 0.0732424
R10491 VSS.n4456 VSS.n4458 2.21488
R10492 VSS.n4461 VSS.n4460 0.0732424
R10493 VSS.n4456 VSS.n4461 2.21488
R10494 VSS.n4470 VSS.n4471 4.5005
R10495 VSS.n4473 VSS.n4472 0.0732424
R10496 VSS.n4471 VSS.n4473 2.21488
R10497 VSS.n4476 VSS.n4475 0.0732424
R10498 VSS.n4471 VSS.n4476 2.21488
R10499 VSS.n4485 VSS.n4486 4.5005
R10500 VSS.n4488 VSS.n4487 0.0732424
R10501 VSS.n4486 VSS.n4488 2.21488
R10502 VSS.n4491 VSS.n4490 0.0732424
R10503 VSS.n4486 VSS.n4491 2.21488
R10504 VSS.n4500 VSS.n4501 4.5005
R10505 VSS.n4503 VSS.n4502 0.0732424
R10506 VSS.n4501 VSS.n4503 2.21488
R10507 VSS.n4506 VSS.n4505 0.0732424
R10508 VSS.n4501 VSS.n4506 2.21488
R10509 VSS.n4515 VSS.n4516 4.5005
R10510 VSS.n4517 VSS.n4518 0.0732424
R10511 VSS.n4518 VSS.n4516 2.21488
R10512 VSS.n4520 VSS.n4521 0.0732424
R10513 VSS.n4521 VSS.n4516 2.21488
R10514 VSS.n4530 VSS.n4531 4.5005
R10515 VSS.n4533 VSS.n4532 0.0732424
R10516 VSS.n4531 VSS.n4533 2.21488
R10517 VSS.n4536 VSS.n4535 0.0732424
R10518 VSS.n4531 VSS.n4536 2.21488
R10519 VSS.n4545 VSS.n4546 4.5005
R10520 VSS.n4548 VSS.n4547 0.0732424
R10521 VSS.n4546 VSS.n4548 2.21488
R10522 VSS.n4551 VSS.n4550 0.0732424
R10523 VSS.n4546 VSS.n4551 2.21488
R10524 VSS.n4560 VSS.n4561 4.5005
R10525 VSS.n4563 VSS.n4562 0.0732424
R10526 VSS.n4561 VSS.n4563 2.21488
R10527 VSS.n4566 VSS.n4565 0.0732424
R10528 VSS.n4561 VSS.n4566 2.21488
R10529 VSS.n4575 VSS.n4576 4.5005
R10530 VSS.n4577 VSS.n4578 0.0732424
R10531 VSS.n4578 VSS.n4576 2.21488
R10532 VSS.n4580 VSS.n4581 0.0732424
R10533 VSS.n4581 VSS.n4576 2.21488
R10534 VSS.n4590 VSS.n4591 4.5005
R10535 VSS.n4593 VSS.n4592 0.0732424
R10536 VSS.n4591 VSS.n4593 2.21488
R10537 VSS.n4596 VSS.n4595 0.0732424
R10538 VSS.n4591 VSS.n4596 2.21488
R10539 VSS.n4605 VSS.n4606 4.5005
R10540 VSS.n4608 VSS.n4607 0.0732424
R10541 VSS.n4606 VSS.n4608 2.21488
R10542 VSS.n4611 VSS.n4610 0.0732424
R10543 VSS.n4606 VSS.n4611 2.21488
R10544 VSS.n4620 VSS.n4621 4.5005
R10545 VSS.n4623 VSS.n4622 0.0732424
R10546 VSS.n4621 VSS.n4623 2.21488
R10547 VSS.n4626 VSS.n4625 0.0732424
R10548 VSS.n4621 VSS.n4626 2.21488
R10549 VSS.n4635 VSS.n4636 4.5005
R10550 VSS.n4638 VSS.n4637 0.0732424
R10551 VSS.n4636 VSS.n4638 2.21488
R10552 VSS.n4641 VSS.n4640 0.0732424
R10553 VSS.n4636 VSS.n4641 2.21488
R10554 VSS.n4650 VSS.n4651 4.5005
R10555 VSS.n4653 VSS.n4652 0.0732424
R10556 VSS.n4651 VSS.n4653 2.21488
R10557 VSS.n4656 VSS.n4655 0.0732424
R10558 VSS.n4651 VSS.n4656 2.21488
R10559 VSS.n4665 VSS.n4666 4.5005
R10560 VSS.n4668 VSS.n4667 0.0732424
R10561 VSS.n4666 VSS.n4668 2.21488
R10562 VSS.n4671 VSS.n4670 0.0732424
R10563 VSS.n4666 VSS.n4671 2.21488
R10564 VSS.n4680 VSS.n4681 4.5005
R10565 VSS.n4682 VSS.n4683 0.0732424
R10566 VSS.n4683 VSS.n4681 2.21488
R10567 VSS.n4685 VSS.n4686 0.0732424
R10568 VSS.n4686 VSS.n4681 2.21488
R10569 VSS.n4695 VSS.n4696 4.5005
R10570 VSS.n4698 VSS.n4697 0.0732424
R10571 VSS.n4696 VSS.n4698 2.21488
R10572 VSS.n4701 VSS.n4700 0.0732424
R10573 VSS.n4696 VSS.n4701 2.21488
R10574 VSS.n4710 VSS.n4711 4.5005
R10575 VSS.n4713 VSS.n4712 0.0732424
R10576 VSS.n4711 VSS.n4713 2.21488
R10577 VSS.n4716 VSS.n4715 0.0732424
R10578 VSS.n4711 VSS.n4716 2.21488
R10579 VSS.n4725 VSS.n4726 4.5005
R10580 VSS.n4728 VSS.n4727 0.0732424
R10581 VSS.n4726 VSS.n4728 2.21488
R10582 VSS.n4731 VSS.n4730 0.0732424
R10583 VSS.n4726 VSS.n4731 2.21488
R10584 VSS.n4740 VSS.n4741 4.5005
R10585 VSS.n4743 VSS.n4742 0.0732424
R10586 VSS.n4741 VSS.n4743 2.21488
R10587 VSS.n4746 VSS.n4745 0.0732424
R10588 VSS.n4741 VSS.n4746 2.21488
R10589 VSS.n4755 VSS.n4756 4.5005
R10590 VSS.n4758 VSS.n4757 0.0732424
R10591 VSS.n4756 VSS.n4758 2.21488
R10592 VSS.n4761 VSS.n4760 0.0732424
R10593 VSS.n4756 VSS.n4761 2.21488
R10594 VSS.n4741 VSS.n4756 0.0584021
R10595 VSS.n2384 VSS.n4741 0.0596608
R10596 VSS.n2384 VSS.n4726 0.0244161
R10597 VSS.n4726 VSS.n4711 0.0585594
R10598 VSS.n4711 VSS.n4696 0.0584021
R10599 VSS.n4681 VSS.n4696 0.0596608
R10600 VSS.n4681 VSS.n4666 0.0244161
R10601 VSS.n4666 VSS.n4651 0.0585594
R10602 VSS.n4651 VSS.n4636 0.0584021
R10603 VSS.n4636 VSS 0.16272
R10604 VSS VSS.n4621 0.143052
R10605 VSS.n4606 VSS.n4621 0.0584021
R10606 VSS.n4591 VSS.n4606 0.0584021
R10607 VSS.n4576 VSS.n4591 0.0244161
R10608 VSS.n4576 VSS.n4561 0.0598182
R10609 VSS.n4561 VSS.n4546 0.0584021
R10610 VSS.n4531 VSS.n4546 0.0584021
R10611 VSS.n4516 VSS.n4531 0.0244161
R10612 VSS.n4516 VSS.n4501 0.0598182
R10613 VSS.n4501 VSS.n4486 0.0584021
R10614 VSS.n4486 VSS.n4471 0.0231573
R10615 VSS.n4456 VSS.n4471 0.0584021
R10616 VSS.n4441 VSS.n4456 0.0596608
R10617 VSS.n4441 VSS.n4426 0.0244161
R10618 VSS.n4426 VSS.n4411 0.0585594
R10619 VSS.n4411 VSS.n4396 0.0584021
R10620 VSS.n4381 VSS.n4396 0.0596608
R10621 VSS.n4381 VSS.n4366 0.0244161
R10622 VSS.n4366 VSS.n4351 0.0585594
R10623 VSS.n4351 VSS.n4336 0.0584021
R10624 VSS.n4336 VSS 0.16272
R10625 VSS VSS.n4321 0.143052
R10626 VSS.n4306 VSS.n4321 0.0584021
R10627 VSS.n4291 VSS.n4306 0.0584021
R10628 VSS.n4276 VSS.n4291 0.0244161
R10629 VSS.n4276 VSS.n4261 0.0598182
R10630 VSS.n4261 VSS.n4246 0.0584021
R10631 VSS.n4231 VSS.n4246 0.0584021
R10632 VSS.n4216 VSS.n4231 0.0244161
R10633 VSS.n4216 VSS.n4201 0.0598182
R10634 VSS.n4201 VSS.n4186 0.0584021
R10635 VSS.n4186 VSS.n4171 0.0231573
R10636 VSS.n4156 VSS.n4171 0.0584021
R10637 VSS.n4141 VSS.n4156 0.0596608
R10638 VSS.n4141 VSS.n4126 0.0244161
R10639 VSS.n4126 VSS.n4111 0.0585594
R10640 VSS.n4111 VSS.n4096 0.0584021
R10641 VSS.n4081 VSS.n4096 0.0596608
R10642 VSS.n4081 VSS.n4066 0.0244161
R10643 VSS.n4066 VSS.n4051 0.0585594
R10644 VSS.n4051 VSS.n4036 0.0584021
R10645 VSS.n4036 VSS 0.16272
R10646 VSS VSS.n4021 0.143052
R10647 VSS.n4006 VSS.n4021 0.0584021
R10648 VSS.n3991 VSS.n4006 0.0584021
R10649 VSS.n3976 VSS.n3991 0.0244161
R10650 VSS.n3976 VSS.n3961 0.0598182
R10651 VSS.n3961 VSS.n3946 0.0584021
R10652 VSS.n3931 VSS.n3946 0.0584021
R10653 VSS.n3916 VSS.n3931 0.0244161
R10654 VSS.n3916 VSS.n3901 0.0598182
R10655 VSS.n3901 VSS.n3886 0.0584021
R10656 VSS.n3886 VSS.n3871 0.0231573
R10657 VSS.n3856 VSS.n3871 0.0584021
R10658 VSS.n3841 VSS.n3856 0.0596608
R10659 VSS.n3841 VSS.n3826 0.0244161
R10660 VSS.n3826 VSS.n3811 0.0585594
R10661 VSS.n3811 VSS.n3796 0.0584021
R10662 VSS.n3781 VSS.n3796 0.0596608
R10663 VSS.n3781 VSS.n3766 0.0244161
R10664 VSS.n3766 VSS.n3751 0.0585594
R10665 VSS.n3751 VSS.n3736 0.0584021
R10666 VSS.n3736 VSS 0.16272
R10667 VSS VSS.n3721 0.143052
R10668 VSS.n3706 VSS.n3721 0.0584021
R10669 VSS.n3691 VSS.n3706 0.0584021
R10670 VSS.n3676 VSS.n3691 0.0244161
R10671 VSS.n3676 VSS.n3661 0.0598182
R10672 VSS.n3661 VSS.n3646 0.0584021
R10673 VSS.n3631 VSS.n3646 0.0584021
R10674 VSS.n3616 VSS.n3631 0.0244161
R10675 VSS.n3616 VSS.n3601 0.0598182
R10676 VSS.n3601 VSS.n3586 0.0584021
R10677 VSS.n3586 VSS.n3571 0.0231573
R10678 VSS.n3556 VSS.n3571 0.0584021
R10679 VSS.n3541 VSS.n3556 0.0596608
R10680 VSS.n3541 VSS.n3526 0.0244161
R10681 VSS.n3526 VSS.n3511 0.0585594
R10682 VSS.n3511 VSS.n3496 0.0584021
R10683 VSS.n3481 VSS.n3496 0.0596608
R10684 VSS.n3481 VSS.n3466 0.0244161
R10685 VSS.n3466 VSS.n3451 0.0585594
R10686 VSS.n3451 VSS.n3436 0.0584021
R10687 VSS.n3436 VSS 0.16272
R10688 VSS VSS.n3421 0.143052
R10689 VSS.n3406 VSS.n3421 0.0584021
R10690 VSS.n3391 VSS.n3406 0.0584021
R10691 VSS.n3376 VSS.n3391 0.0244161
R10692 VSS.n3376 VSS.n3361 0.0598182
R10693 VSS.n3361 VSS.n3346 0.0584021
R10694 VSS.n3331 VSS.n3346 0.0584021
R10695 VSS.n3316 VSS.n3331 0.0244161
R10696 VSS.n3316 VSS.n3301 0.0598182
R10697 VSS.n3301 VSS.n3286 0.0584021
R10698 VSS.n3286 VSS.n3271 0.0231573
R10699 VSS.n3256 VSS.n3271 0.0584021
R10700 VSS.n3241 VSS.n3256 0.0596608
R10701 VSS.n3241 VSS.n3226 0.0244161
R10702 VSS.n3226 VSS.n3211 0.0585594
R10703 VSS.n3211 VSS.n3196 0.0584021
R10704 VSS.n3181 VSS.n3196 0.0596608
R10705 VSS.n3181 VSS.n3166 0.0244161
R10706 VSS.n3166 VSS.n3151 0.0585594
R10707 VSS.n3151 VSS.n3136 0.0584021
R10708 VSS.n3136 VSS 0.16272
R10709 VSS VSS.n3121 0.143052
R10710 VSS.n3106 VSS.n3121 0.0584021
R10711 VSS.n3091 VSS.n3106 0.0584021
R10712 VSS.n3076 VSS.n3091 0.0244161
R10713 VSS.n3076 VSS.n3061 0.0598182
R10714 VSS.n3061 VSS.n3046 0.0584021
R10715 VSS.n3031 VSS.n3046 0.0584021
R10716 VSS.n3016 VSS.n3031 0.0244161
R10717 VSS.n3016 VSS.n3001 0.0598182
R10718 VSS.n3001 VSS.n2986 0.0584021
R10719 VSS.n2986 VSS.n2971 0.0231573
R10720 VSS.n2956 VSS.n2971 0.0584021
R10721 VSS.n2941 VSS.n2956 0.0596608
R10722 VSS.n2941 VSS.n2926 0.0244161
R10723 VSS.n2926 VSS.n2911 0.0585594
R10724 VSS.n2911 VSS.n2896 0.0584021
R10725 VSS.n2881 VSS.n2896 0.0596608
R10726 VSS.n2881 VSS.n2866 0.0244161
R10727 VSS.n2866 VSS.n2851 0.0585594
R10728 VSS.n2851 VSS.n2836 0.0584021
R10729 VSS.n2836 VSS 0.16272
R10730 VSS VSS.n2821 0.143052
R10731 VSS.n2806 VSS.n2821 0.0584021
R10732 VSS.n2791 VSS.n2806 0.0584021
R10733 VSS.n2776 VSS.n2791 0.0244161
R10734 VSS.n2776 VSS.n2761 0.0598182
R10735 VSS.n2761 VSS.n2746 0.0584021
R10736 VSS.n2731 VSS.n2746 0.0584021
R10737 VSS.n2716 VSS.n2731 0.0244161
R10738 VSS.n2716 VSS.n2701 0.0598182
R10739 VSS.n2701 VSS.n2686 0.0584021
R10740 VSS.n2686 VSS.n2671 0.0231573
R10741 VSS.n2656 VSS.n2671 0.0584021
R10742 VSS.n2641 VSS.n2656 0.0596608
R10743 VSS.n2641 VSS.n2626 0.0244161
R10744 VSS.n2626 VSS.n2611 0.0585594
R10745 VSS.n2611 VSS.n2596 0.0584021
R10746 VSS.n2581 VSS.n2596 0.0596608
R10747 VSS.n2581 VSS.n2566 0.0244161
R10748 VSS.n2566 VSS.n2551 0.0585594
R10749 VSS.n2551 VSS.n2536 0.0584021
R10750 VSS.n2536 VSS 0.16272
R10751 VSS VSS.n2521 0.143052
R10752 VSS.n2506 VSS.n2521 0.0584021
R10753 VSS.n2491 VSS.n2506 0.0584021
R10754 VSS.n2476 VSS.n2491 0.0244161
R10755 VSS.n2476 VSS.n2461 0.0598182
R10756 VSS.n2461 VSS.n2446 0.0584021
R10757 VSS.n2431 VSS.n2446 0.0584021
R10758 VSS.n2416 VSS.n2431 0.0244161
R10759 VSS.n2416 VSS.n2401 0.0598182
R10760 VSS.n2401 VSS.n2386 0.0584021
R10761 VSS.n4757 VSS.n4762 4.5005
R10762 VSS.n4759 VSS.n4763 4.5005
R10763 VSS.n4760 VSS.n4764 4.5005
R10764 VSS.n4761 VSS.n4765 4.57324
R10765 VSS.n4757 VSS.n4755 0.147342
R10766 VSS.n4758 VSS.n4759 0.0732424
R10767 VSS.n4759 VSS.n4760 0.147342
R10768 VSS.n4762 VSS.n4766 0.0721009
R10769 VSS.n4767 VSS.n4763 4.5005
R10770 VSS.n4768 VSS.n4764 4.5005
R10771 VSS.n4769 VSS.n4765 4.5005
R10772 VSS.n4755 VSS.n4766 4.57442
R10773 VSS.n4762 VSS.n4763 0.147342
R10774 VSS.n4763 VSS.n4764 0.147342
R10775 VSS.n4764 VSS.n4765 0.147342
R10776 VSS.n4766 VSS.n4767 2.39784
R10777 VSS.n4767 VSS.n4768 0.147342
R10778 VSS.n4768 VSS.n4769 0.147342
R10779 VSS.n4769 VSS.t247 3.13212
R10780 VSS.n4742 VSS.n4747 4.5005
R10781 VSS.n4744 VSS.n4748 4.5005
R10782 VSS.n4745 VSS.n4749 4.5005
R10783 VSS.n4746 VSS.n4750 4.57324
R10784 VSS.n4742 VSS.n4740 0.147342
R10785 VSS.n4743 VSS.n4744 0.0732424
R10786 VSS.n4744 VSS.n4745 0.147342
R10787 VSS.n4747 VSS.n4751 0.0721009
R10788 VSS.n4752 VSS.n4748 4.5005
R10789 VSS.n4753 VSS.n4749 4.5005
R10790 VSS.n4754 VSS.n4750 4.5005
R10791 VSS.n4740 VSS.n4751 4.57442
R10792 VSS.n4747 VSS.n4748 0.147342
R10793 VSS.n4748 VSS.n4749 0.147342
R10794 VSS.n4749 VSS.n4750 0.147342
R10795 VSS.n4751 VSS.n4752 2.39784
R10796 VSS.n4752 VSS.n4753 0.147342
R10797 VSS.n4753 VSS.n4754 0.147342
R10798 VSS.n4754 VSS.t250 3.13212
R10799 VSS.n4727 VSS.n4732 4.5005
R10800 VSS.n4729 VSS.n4733 4.5005
R10801 VSS.n4730 VSS.n4734 4.5005
R10802 VSS.n4731 VSS.n4735 4.57324
R10803 VSS.n4727 VSS.n4725 0.147342
R10804 VSS.n4728 VSS.n4729 0.0732424
R10805 VSS.n4729 VSS.n4730 0.147342
R10806 VSS.n4732 VSS.n4736 0.0721009
R10807 VSS.n4737 VSS.n4733 4.5005
R10808 VSS.n4738 VSS.n4734 4.5005
R10809 VSS.n4739 VSS.n4735 4.5005
R10810 VSS.n4725 VSS.n4736 4.57442
R10811 VSS.n4732 VSS.n4733 0.147342
R10812 VSS.n4733 VSS.n4734 0.147342
R10813 VSS.n4734 VSS.n4735 0.147342
R10814 VSS.n4736 VSS.n4737 2.39784
R10815 VSS.n4737 VSS.n4738 0.147342
R10816 VSS.n4738 VSS.n4739 0.147342
R10817 VSS.n4739 VSS.t403 3.13212
R10818 VSS.n4712 VSS.n4717 4.5005
R10819 VSS.n4714 VSS.n4718 4.5005
R10820 VSS.n4715 VSS.n4719 4.5005
R10821 VSS.n4716 VSS.n4720 4.57324
R10822 VSS.n4712 VSS.n4710 0.147342
R10823 VSS.n4713 VSS.n4714 0.0732424
R10824 VSS.n4714 VSS.n4715 0.147342
R10825 VSS.n4717 VSS.n4721 0.0721009
R10826 VSS.n4722 VSS.n4718 4.5005
R10827 VSS.n4723 VSS.n4719 4.5005
R10828 VSS.n4724 VSS.n4720 4.5005
R10829 VSS.n4710 VSS.n4721 4.57442
R10830 VSS.n4717 VSS.n4718 0.147342
R10831 VSS.n4718 VSS.n4719 0.147342
R10832 VSS.n4719 VSS.n4720 0.147342
R10833 VSS.n4721 VSS.n4722 2.39784
R10834 VSS.n4722 VSS.n4723 0.147342
R10835 VSS.n4723 VSS.n4724 0.147342
R10836 VSS.n4724 VSS.t85 3.13212
R10837 VSS.n4697 VSS.n4702 4.5005
R10838 VSS.n4699 VSS.n4703 4.5005
R10839 VSS.n4700 VSS.n4704 4.5005
R10840 VSS.n4701 VSS.n4705 4.57324
R10841 VSS.n4697 VSS.n4695 0.147342
R10842 VSS.n4698 VSS.n4699 0.0732424
R10843 VSS.n4699 VSS.n4700 0.147342
R10844 VSS.n4702 VSS.n4706 0.0721009
R10845 VSS.n4707 VSS.n4703 4.5005
R10846 VSS.n4708 VSS.n4704 4.5005
R10847 VSS.n4709 VSS.n4705 4.5005
R10848 VSS.n4695 VSS.n4706 4.57442
R10849 VSS.n4702 VSS.n4703 0.147342
R10850 VSS.n4703 VSS.n4704 0.147342
R10851 VSS.n4704 VSS.n4705 0.147342
R10852 VSS.n4706 VSS.n4707 2.39784
R10853 VSS.n4707 VSS.n4708 0.147342
R10854 VSS.n4708 VSS.n4709 0.147342
R10855 VSS.n4709 VSS.t517 3.13212
R10856 VSS.n4687 VSS.n4682 4.5005
R10857 VSS.n4688 VSS.n4684 4.5005
R10858 VSS.n4689 VSS.n4685 4.5005
R10859 VSS.n4690 VSS.n4686 4.57324
R10860 VSS.n4680 VSS.n4682 0.147342
R10861 VSS.n4683 VSS.n4684 0.0732424
R10862 VSS.n4684 VSS.n4685 0.147342
R10863 VSS.n4691 VSS.n4687 0.0722544
R10864 VSS.n4692 VSS.n4688 4.5005
R10865 VSS.n4693 VSS.n4689 4.5005
R10866 VSS.n4694 VSS.n4690 4.5005
R10867 VSS.n4691 VSS.n4680 4.57426
R10868 VSS.n4687 VSS.n4688 0.147342
R10869 VSS.n4688 VSS.n4689 0.147342
R10870 VSS.n4689 VSS.n4690 0.147342
R10871 VSS.n4692 VSS.n4691 2.37296
R10872 VSS.n4693 VSS.n4692 0.127318
R10873 VSS.n4694 VSS.n4693 0.127318
R10874 VSS.t5 VSS.n4694 2.73618
R10875 VSS.n4667 VSS.n4672 4.5005
R10876 VSS.n4669 VSS.n4673 4.5005
R10877 VSS.n4670 VSS.n4674 4.5005
R10878 VSS.n4671 VSS.n4675 4.57324
R10879 VSS.n4667 VSS.n4665 0.147342
R10880 VSS.n4668 VSS.n4669 0.0732424
R10881 VSS.n4669 VSS.n4670 0.147342
R10882 VSS.n4672 VSS.n4676 0.0721009
R10883 VSS.n4677 VSS.n4673 4.5005
R10884 VSS.n4678 VSS.n4674 4.5005
R10885 VSS.n4679 VSS.n4675 4.5005
R10886 VSS.n4665 VSS.n4676 4.57442
R10887 VSS.n4672 VSS.n4673 0.147342
R10888 VSS.n4673 VSS.n4674 0.147342
R10889 VSS.n4674 VSS.n4675 0.147342
R10890 VSS.n4676 VSS.n4677 2.39784
R10891 VSS.n4677 VSS.n4678 0.147342
R10892 VSS.n4678 VSS.n4679 0.147342
R10893 VSS.n4679 VSS.t619 3.13212
R10894 VSS.n4652 VSS.n4657 4.5005
R10895 VSS.n4654 VSS.n4658 4.5005
R10896 VSS.n4655 VSS.n4659 4.5005
R10897 VSS.n4656 VSS.n4660 4.57324
R10898 VSS.n4652 VSS.n4650 0.147342
R10899 VSS.n4653 VSS.n4654 0.0732424
R10900 VSS.n4654 VSS.n4655 0.147342
R10901 VSS.n4657 VSS.n4661 0.0721009
R10902 VSS.n4662 VSS.n4658 4.5005
R10903 VSS.n4663 VSS.n4659 4.5005
R10904 VSS.n4664 VSS.n4660 4.5005
R10905 VSS.n4650 VSS.n4661 4.57442
R10906 VSS.n4657 VSS.n4658 0.147342
R10907 VSS.n4658 VSS.n4659 0.147342
R10908 VSS.n4659 VSS.n4660 0.147342
R10909 VSS.n4661 VSS.n4662 2.39784
R10910 VSS.n4662 VSS.n4663 0.147342
R10911 VSS.n4663 VSS.n4664 0.147342
R10912 VSS.n4664 VSS.t184 3.13212
R10913 VSS.n4637 VSS.n4642 4.5005
R10914 VSS.n4639 VSS.n4643 4.5005
R10915 VSS.n4640 VSS.n4644 4.5005
R10916 VSS.n4641 VSS.n4645 4.57324
R10917 VSS.n4637 VSS.n4635 0.147342
R10918 VSS.n4638 VSS.n4639 0.0732424
R10919 VSS.n4639 VSS.n4640 0.147342
R10920 VSS.n4642 VSS.n4646 0.0721009
R10921 VSS.n4647 VSS.n4643 4.5005
R10922 VSS.n4648 VSS.n4644 4.5005
R10923 VSS.n4649 VSS.n4645 4.5005
R10924 VSS.n4635 VSS.n4646 4.57442
R10925 VSS.n4642 VSS.n4643 0.147342
R10926 VSS.n4643 VSS.n4644 0.147342
R10927 VSS.n4644 VSS.n4645 0.147342
R10928 VSS.n4646 VSS.n4647 2.39784
R10929 VSS.n4647 VSS.n4648 0.147342
R10930 VSS.n4648 VSS.n4649 0.147342
R10931 VSS.n4649 VSS.t107 3.13212
R10932 VSS.n4622 VSS.n4627 4.5005
R10933 VSS.n4624 VSS.n4628 4.5005
R10934 VSS.n4625 VSS.n4629 4.5005
R10935 VSS.n4626 VSS.n4630 4.57324
R10936 VSS.n4622 VSS.n4620 0.147342
R10937 VSS.n4623 VSS.n4624 0.0732424
R10938 VSS.n4624 VSS.n4625 0.147342
R10939 VSS.n4627 VSS.n4631 0.0721009
R10940 VSS.n4632 VSS.n4628 4.5005
R10941 VSS.n4633 VSS.n4629 4.5005
R10942 VSS.n4634 VSS.n4630 4.5005
R10943 VSS.n4620 VSS.n4631 4.57442
R10944 VSS.n4627 VSS.n4628 0.147342
R10945 VSS.n4628 VSS.n4629 0.147342
R10946 VSS.n4629 VSS.n4630 0.147342
R10947 VSS.n4631 VSS.n4632 2.39784
R10948 VSS.n4632 VSS.n4633 0.147342
R10949 VSS.n4633 VSS.n4634 0.147342
R10950 VSS.n4634 VSS.t13 3.13212
R10951 VSS.n4607 VSS.n4612 4.5005
R10952 VSS.n4609 VSS.n4613 4.5005
R10953 VSS.n4610 VSS.n4614 4.5005
R10954 VSS.n4611 VSS.n4615 4.57324
R10955 VSS.n4607 VSS.n4605 0.147342
R10956 VSS.n4608 VSS.n4609 0.0732424
R10957 VSS.n4609 VSS.n4610 0.147342
R10958 VSS.n4612 VSS.n4616 0.0721009
R10959 VSS.n4617 VSS.n4613 4.5005
R10960 VSS.n4618 VSS.n4614 4.5005
R10961 VSS.n4619 VSS.n4615 4.5005
R10962 VSS.n4605 VSS.n4616 4.57442
R10963 VSS.n4612 VSS.n4613 0.147342
R10964 VSS.n4613 VSS.n4614 0.147342
R10965 VSS.n4614 VSS.n4615 0.147342
R10966 VSS.n4616 VSS.n4617 2.39784
R10967 VSS.n4617 VSS.n4618 0.147342
R10968 VSS.n4618 VSS.n4619 0.147342
R10969 VSS.n4619 VSS.t603 3.13212
R10970 VSS.n4592 VSS.n4597 4.5005
R10971 VSS.n4594 VSS.n4598 4.5005
R10972 VSS.n4595 VSS.n4599 4.5005
R10973 VSS.n4596 VSS.n4600 4.57324
R10974 VSS.n4592 VSS.n4590 0.147342
R10975 VSS.n4593 VSS.n4594 0.0732424
R10976 VSS.n4594 VSS.n4595 0.147342
R10977 VSS.n4597 VSS.n4601 0.0721009
R10978 VSS.n4602 VSS.n4598 4.5005
R10979 VSS.n4603 VSS.n4599 4.5005
R10980 VSS.n4604 VSS.n4600 4.5005
R10981 VSS.n4590 VSS.n4601 4.57442
R10982 VSS.n4597 VSS.n4598 0.147342
R10983 VSS.n4598 VSS.n4599 0.147342
R10984 VSS.n4599 VSS.n4600 0.147342
R10985 VSS.n4601 VSS.n4602 2.39784
R10986 VSS.n4602 VSS.n4603 0.147342
R10987 VSS.n4603 VSS.n4604 0.147342
R10988 VSS.n4604 VSS.t495 3.13212
R10989 VSS.n4582 VSS.n4577 4.5005
R10990 VSS.n4583 VSS.n4579 4.5005
R10991 VSS.n4584 VSS.n4580 4.5005
R10992 VSS.n4585 VSS.n4581 4.57324
R10993 VSS.n4575 VSS.n4577 0.147342
R10994 VSS.n4578 VSS.n4579 0.0732424
R10995 VSS.n4579 VSS.n4580 0.147342
R10996 VSS.n4586 VSS.n4582 0.0722544
R10997 VSS.n4587 VSS.n4583 4.5005
R10998 VSS.n4588 VSS.n4584 4.5005
R10999 VSS.n4589 VSS.n4585 4.5005
R11000 VSS.n4586 VSS.n4575 4.57426
R11001 VSS.n4582 VSS.n4583 0.147342
R11002 VSS.n4583 VSS.n4584 0.147342
R11003 VSS.n4584 VSS.n4585 0.147342
R11004 VSS.n4587 VSS.n4586 2.37296
R11005 VSS.n4588 VSS.n4587 0.127318
R11006 VSS.n4589 VSS.n4588 0.127318
R11007 VSS.t5 VSS.n4589 2.73618
R11008 VSS.n4562 VSS.n4567 4.5005
R11009 VSS.n4564 VSS.n4568 4.5005
R11010 VSS.n4565 VSS.n4569 4.5005
R11011 VSS.n4566 VSS.n4570 4.57324
R11012 VSS.n4562 VSS.n4560 0.147342
R11013 VSS.n4563 VSS.n4564 0.0732424
R11014 VSS.n4564 VSS.n4565 0.147342
R11015 VSS.n4567 VSS.n4571 0.0721009
R11016 VSS.n4572 VSS.n4568 4.5005
R11017 VSS.n4573 VSS.n4569 4.5005
R11018 VSS.n4574 VSS.n4570 4.5005
R11019 VSS.n4560 VSS.n4571 4.57442
R11020 VSS.n4567 VSS.n4568 0.147342
R11021 VSS.n4568 VSS.n4569 0.147342
R11022 VSS.n4569 VSS.n4570 0.147342
R11023 VSS.n4571 VSS.n4572 2.39784
R11024 VSS.n4572 VSS.n4573 0.147342
R11025 VSS.n4573 VSS.n4574 0.147342
R11026 VSS.n4574 VSS.t347 3.13212
R11027 VSS.n4547 VSS.n4552 4.5005
R11028 VSS.n4549 VSS.n4553 4.5005
R11029 VSS.n4550 VSS.n4554 4.5005
R11030 VSS.n4551 VSS.n4555 4.57324
R11031 VSS.n4547 VSS.n4545 0.147342
R11032 VSS.n4548 VSS.n4549 0.0732424
R11033 VSS.n4549 VSS.n4550 0.147342
R11034 VSS.n4552 VSS.n4556 0.0721009
R11035 VSS.n4557 VSS.n4553 4.5005
R11036 VSS.n4558 VSS.n4554 4.5005
R11037 VSS.n4559 VSS.n4555 4.5005
R11038 VSS.n4545 VSS.n4556 4.57442
R11039 VSS.n4552 VSS.n4553 0.147342
R11040 VSS.n4553 VSS.n4554 0.147342
R11041 VSS.n4554 VSS.n4555 0.147342
R11042 VSS.n4556 VSS.n4557 2.39784
R11043 VSS.n4557 VSS.n4558 0.147342
R11044 VSS.n4558 VSS.n4559 0.147342
R11045 VSS.n4559 VSS.t36 3.13212
R11046 VSS.n4532 VSS.n4537 4.5005
R11047 VSS.n4534 VSS.n4538 4.5005
R11048 VSS.n4535 VSS.n4539 4.5005
R11049 VSS.n4536 VSS.n4540 4.57324
R11050 VSS.n4532 VSS.n4530 0.147342
R11051 VSS.n4533 VSS.n4534 0.0732424
R11052 VSS.n4534 VSS.n4535 0.147342
R11053 VSS.n4537 VSS.n4541 0.0721009
R11054 VSS.n4542 VSS.n4538 4.5005
R11055 VSS.n4543 VSS.n4539 4.5005
R11056 VSS.n4544 VSS.n4540 4.5005
R11057 VSS.n4530 VSS.n4541 4.57442
R11058 VSS.n4537 VSS.n4538 0.147342
R11059 VSS.n4538 VSS.n4539 0.147342
R11060 VSS.n4539 VSS.n4540 0.147342
R11061 VSS.n4541 VSS.n4542 2.39784
R11062 VSS.n4542 VSS.n4543 0.147342
R11063 VSS.n4543 VSS.n4544 0.147342
R11064 VSS.n4544 VSS.t14 3.13212
R11065 VSS.n4522 VSS.n4517 4.5005
R11066 VSS.n4523 VSS.n4519 4.5005
R11067 VSS.n4524 VSS.n4520 4.5005
R11068 VSS.n4525 VSS.n4521 4.57324
R11069 VSS.n4515 VSS.n4517 0.147342
R11070 VSS.n4518 VSS.n4519 0.0732424
R11071 VSS.n4519 VSS.n4520 0.147342
R11072 VSS.n4526 VSS.n4522 0.0722544
R11073 VSS.n4527 VSS.n4523 4.5005
R11074 VSS.n4528 VSS.n4524 4.5005
R11075 VSS.n4529 VSS.n4525 4.5005
R11076 VSS.n4526 VSS.n4515 4.57426
R11077 VSS.n4522 VSS.n4523 0.147342
R11078 VSS.n4523 VSS.n4524 0.147342
R11079 VSS.n4524 VSS.n4525 0.147342
R11080 VSS.n4527 VSS.n4526 2.37296
R11081 VSS.n4528 VSS.n4527 0.127318
R11082 VSS.n4529 VSS.n4528 0.127318
R11083 VSS.t5 VSS.n4529 2.73618
R11084 VSS.n4502 VSS.n4507 4.5005
R11085 VSS.n4504 VSS.n4508 4.5005
R11086 VSS.n4505 VSS.n4509 4.5005
R11087 VSS.n4506 VSS.n4510 4.57324
R11088 VSS.n4502 VSS.n4500 0.147342
R11089 VSS.n4503 VSS.n4504 0.0732424
R11090 VSS.n4504 VSS.n4505 0.147342
R11091 VSS.n4507 VSS.n4511 0.0721009
R11092 VSS.n4512 VSS.n4508 4.5005
R11093 VSS.n4513 VSS.n4509 4.5005
R11094 VSS.n4514 VSS.n4510 4.5005
R11095 VSS.n4500 VSS.n4511 4.57442
R11096 VSS.n4507 VSS.n4508 0.147342
R11097 VSS.n4508 VSS.n4509 0.147342
R11098 VSS.n4509 VSS.n4510 0.147342
R11099 VSS.n4511 VSS.n4512 2.39784
R11100 VSS.n4512 VSS.n4513 0.147342
R11101 VSS.n4513 VSS.n4514 0.147342
R11102 VSS.n4514 VSS.t230 3.13212
R11103 VSS.n4487 VSS.n4492 4.5005
R11104 VSS.n4489 VSS.n4493 4.5005
R11105 VSS.n4490 VSS.n4494 4.5005
R11106 VSS.n4491 VSS.n4495 4.57324
R11107 VSS.n4487 VSS.n4485 0.147342
R11108 VSS.n4488 VSS.n4489 0.0732424
R11109 VSS.n4489 VSS.n4490 0.147342
R11110 VSS.n4492 VSS.n4496 0.0721009
R11111 VSS.n4497 VSS.n4493 4.5005
R11112 VSS.n4498 VSS.n4494 4.5005
R11113 VSS.n4499 VSS.n4495 4.5005
R11114 VSS.n4485 VSS.n4496 4.57442
R11115 VSS.n4492 VSS.n4493 0.147342
R11116 VSS.n4493 VSS.n4494 0.147342
R11117 VSS.n4494 VSS.n4495 0.147342
R11118 VSS.n4496 VSS.n4497 2.39784
R11119 VSS.n4497 VSS.n4498 0.147342
R11120 VSS.n4498 VSS.n4499 0.147342
R11121 VSS.n4499 VSS.t467 3.13212
R11122 VSS.n4472 VSS.n4477 4.5005
R11123 VSS.n4474 VSS.n4478 4.5005
R11124 VSS.n4475 VSS.n4479 4.5005
R11125 VSS.n4476 VSS.n4480 4.57324
R11126 VSS.n4472 VSS.n4470 0.147342
R11127 VSS.n4473 VSS.n4474 0.0732424
R11128 VSS.n4474 VSS.n4475 0.147342
R11129 VSS.n4477 VSS.n4481 0.0721009
R11130 VSS.n4482 VSS.n4478 4.5005
R11131 VSS.n4483 VSS.n4479 4.5005
R11132 VSS.n4484 VSS.n4480 4.5005
R11133 VSS.n4470 VSS.n4481 4.57442
R11134 VSS.n4477 VSS.n4478 0.147342
R11135 VSS.n4478 VSS.n4479 0.147342
R11136 VSS.n4479 VSS.n4480 0.147342
R11137 VSS.n4481 VSS.n4482 2.39784
R11138 VSS.n4482 VSS.n4483 0.147342
R11139 VSS.n4483 VSS.n4484 0.147342
R11140 VSS.n4484 VSS.t246 3.13212
R11141 VSS.n4457 VSS.n4462 4.5005
R11142 VSS.n4459 VSS.n4463 4.5005
R11143 VSS.n4460 VSS.n4464 4.5005
R11144 VSS.n4461 VSS.n4465 4.57324
R11145 VSS.n4457 VSS.n4455 0.147342
R11146 VSS.n4458 VSS.n4459 0.0732424
R11147 VSS.n4459 VSS.n4460 0.147342
R11148 VSS.n4462 VSS.n4466 0.0721009
R11149 VSS.n4467 VSS.n4463 4.5005
R11150 VSS.n4468 VSS.n4464 4.5005
R11151 VSS.n4469 VSS.n4465 4.5005
R11152 VSS.n4455 VSS.n4466 4.57442
R11153 VSS.n4462 VSS.n4463 0.147342
R11154 VSS.n4463 VSS.n4464 0.147342
R11155 VSS.n4464 VSS.n4465 0.147342
R11156 VSS.n4466 VSS.n4467 2.39784
R11157 VSS.n4467 VSS.n4468 0.147342
R11158 VSS.n4468 VSS.n4469 0.147342
R11159 VSS.n4469 VSS.t251 3.13212
R11160 VSS.n4447 VSS.n4442 4.5005
R11161 VSS.n4448 VSS.n4444 4.5005
R11162 VSS.n4449 VSS.n4445 4.5005
R11163 VSS.n4450 VSS.n4446 4.57324
R11164 VSS.n4440 VSS.n4442 0.147342
R11165 VSS.n4443 VSS.n4444 0.0732424
R11166 VSS.n4444 VSS.n4445 0.147342
R11167 VSS.n4451 VSS.n4447 0.0722544
R11168 VSS.n4452 VSS.n4448 4.5005
R11169 VSS.n4453 VSS.n4449 4.5005
R11170 VSS.n4454 VSS.n4450 4.5005
R11171 VSS.n4451 VSS.n4440 4.57426
R11172 VSS.n4447 VSS.n4448 0.147342
R11173 VSS.n4448 VSS.n4449 0.147342
R11174 VSS.n4449 VSS.n4450 0.147342
R11175 VSS.n4452 VSS.n4451 2.37296
R11176 VSS.n4453 VSS.n4452 0.127318
R11177 VSS.n4454 VSS.n4453 0.127318
R11178 VSS.t5 VSS.n4454 2.73618
R11179 VSS.n4427 VSS.n4432 4.5005
R11180 VSS.n4429 VSS.n4433 4.5005
R11181 VSS.n4430 VSS.n4434 4.5005
R11182 VSS.n4431 VSS.n4435 4.57324
R11183 VSS.n4427 VSS.n4425 0.147342
R11184 VSS.n4428 VSS.n4429 0.0732424
R11185 VSS.n4429 VSS.n4430 0.147342
R11186 VSS.n4432 VSS.n4436 0.0721009
R11187 VSS.n4437 VSS.n4433 4.5005
R11188 VSS.n4438 VSS.n4434 4.5005
R11189 VSS.n4439 VSS.n4435 4.5005
R11190 VSS.n4425 VSS.n4436 4.57442
R11191 VSS.n4432 VSS.n4433 0.147342
R11192 VSS.n4433 VSS.n4434 0.147342
R11193 VSS.n4434 VSS.n4435 0.147342
R11194 VSS.n4436 VSS.n4437 2.39784
R11195 VSS.n4437 VSS.n4438 0.147342
R11196 VSS.n4438 VSS.n4439 0.147342
R11197 VSS.n4439 VSS.t415 3.13212
R11198 VSS.n4412 VSS.n4417 4.5005
R11199 VSS.n4414 VSS.n4418 4.5005
R11200 VSS.n4415 VSS.n4419 4.5005
R11201 VSS.n4416 VSS.n4420 4.57324
R11202 VSS.n4412 VSS.n4410 0.147342
R11203 VSS.n4413 VSS.n4414 0.0732424
R11204 VSS.n4414 VSS.n4415 0.147342
R11205 VSS.n4417 VSS.n4421 0.0721009
R11206 VSS.n4422 VSS.n4418 4.5005
R11207 VSS.n4423 VSS.n4419 4.5005
R11208 VSS.n4424 VSS.n4420 4.5005
R11209 VSS.n4410 VSS.n4421 4.57442
R11210 VSS.n4417 VSS.n4418 0.147342
R11211 VSS.n4418 VSS.n4419 0.147342
R11212 VSS.n4419 VSS.n4420 0.147342
R11213 VSS.n4421 VSS.n4422 2.39784
R11214 VSS.n4422 VSS.n4423 0.147342
R11215 VSS.n4423 VSS.n4424 0.147342
R11216 VSS.n4424 VSS.t92 3.13212
R11217 VSS.n4397 VSS.n4402 4.5005
R11218 VSS.n4399 VSS.n4403 4.5005
R11219 VSS.n4400 VSS.n4404 4.5005
R11220 VSS.n4401 VSS.n4405 4.57324
R11221 VSS.n4397 VSS.n4395 0.147342
R11222 VSS.n4398 VSS.n4399 0.0732424
R11223 VSS.n4399 VSS.n4400 0.147342
R11224 VSS.n4402 VSS.n4406 0.0721009
R11225 VSS.n4407 VSS.n4403 4.5005
R11226 VSS.n4408 VSS.n4404 4.5005
R11227 VSS.n4409 VSS.n4405 4.5005
R11228 VSS.n4395 VSS.n4406 4.57442
R11229 VSS.n4402 VSS.n4403 0.147342
R11230 VSS.n4403 VSS.n4404 0.147342
R11231 VSS.n4404 VSS.n4405 0.147342
R11232 VSS.n4406 VSS.n4407 2.39784
R11233 VSS.n4407 VSS.n4408 0.147342
R11234 VSS.n4408 VSS.n4409 0.147342
R11235 VSS.n4409 VSS.t122 3.13212
R11236 VSS.n4387 VSS.n4382 4.5005
R11237 VSS.n4388 VSS.n4384 4.5005
R11238 VSS.n4389 VSS.n4385 4.5005
R11239 VSS.n4390 VSS.n4386 4.57324
R11240 VSS.n4380 VSS.n4382 0.147342
R11241 VSS.n4383 VSS.n4384 0.0732424
R11242 VSS.n4384 VSS.n4385 0.147342
R11243 VSS.n4391 VSS.n4387 0.0722544
R11244 VSS.n4392 VSS.n4388 4.5005
R11245 VSS.n4393 VSS.n4389 4.5005
R11246 VSS.n4394 VSS.n4390 4.5005
R11247 VSS.n4391 VSS.n4380 4.57426
R11248 VSS.n4387 VSS.n4388 0.147342
R11249 VSS.n4388 VSS.n4389 0.147342
R11250 VSS.n4389 VSS.n4390 0.147342
R11251 VSS.n4392 VSS.n4391 2.37296
R11252 VSS.n4393 VSS.n4392 0.127318
R11253 VSS.n4394 VSS.n4393 0.127318
R11254 VSS.t5 VSS.n4394 2.73618
R11255 VSS.n4367 VSS.n4372 4.5005
R11256 VSS.n4369 VSS.n4373 4.5005
R11257 VSS.n4370 VSS.n4374 4.5005
R11258 VSS.n4371 VSS.n4375 4.57324
R11259 VSS.n4367 VSS.n4365 0.147342
R11260 VSS.n4368 VSS.n4369 0.0732424
R11261 VSS.n4369 VSS.n4370 0.147342
R11262 VSS.n4372 VSS.n4376 0.0721009
R11263 VSS.n4377 VSS.n4373 4.5005
R11264 VSS.n4378 VSS.n4374 4.5005
R11265 VSS.n4379 VSS.n4375 4.5005
R11266 VSS.n4365 VSS.n4376 4.57442
R11267 VSS.n4372 VSS.n4373 0.147342
R11268 VSS.n4373 VSS.n4374 0.147342
R11269 VSS.n4374 VSS.n4375 0.147342
R11270 VSS.n4376 VSS.n4377 2.39784
R11271 VSS.n4377 VSS.n4378 0.147342
R11272 VSS.n4378 VSS.n4379 0.147342
R11273 VSS.n4379 VSS.t73 3.13212
R11274 VSS.n4352 VSS.n4357 4.5005
R11275 VSS.n4354 VSS.n4358 4.5005
R11276 VSS.n4355 VSS.n4359 4.5005
R11277 VSS.n4356 VSS.n4360 4.57324
R11278 VSS.n4352 VSS.n4350 0.147342
R11279 VSS.n4353 VSS.n4354 0.0732424
R11280 VSS.n4354 VSS.n4355 0.147342
R11281 VSS.n4357 VSS.n4361 0.0721009
R11282 VSS.n4362 VSS.n4358 4.5005
R11283 VSS.n4363 VSS.n4359 4.5005
R11284 VSS.n4364 VSS.n4360 4.5005
R11285 VSS.n4350 VSS.n4361 4.57442
R11286 VSS.n4357 VSS.n4358 0.147342
R11287 VSS.n4358 VSS.n4359 0.147342
R11288 VSS.n4359 VSS.n4360 0.147342
R11289 VSS.n4361 VSS.n4362 2.39784
R11290 VSS.n4362 VSS.n4363 0.147342
R11291 VSS.n4363 VSS.n4364 0.147342
R11292 VSS.n4364 VSS.t189 3.13212
R11293 VSS.n4337 VSS.n4342 4.5005
R11294 VSS.n4339 VSS.n4343 4.5005
R11295 VSS.n4340 VSS.n4344 4.5005
R11296 VSS.n4341 VSS.n4345 4.57324
R11297 VSS.n4337 VSS.n4335 0.147342
R11298 VSS.n4338 VSS.n4339 0.0732424
R11299 VSS.n4339 VSS.n4340 0.147342
R11300 VSS.n4342 VSS.n4346 0.0721009
R11301 VSS.n4347 VSS.n4343 4.5005
R11302 VSS.n4348 VSS.n4344 4.5005
R11303 VSS.n4349 VSS.n4345 4.5005
R11304 VSS.n4335 VSS.n4346 4.57442
R11305 VSS.n4342 VSS.n4343 0.147342
R11306 VSS.n4343 VSS.n4344 0.147342
R11307 VSS.n4344 VSS.n4345 0.147342
R11308 VSS.n4346 VSS.n4347 2.39784
R11309 VSS.n4347 VSS.n4348 0.147342
R11310 VSS.n4348 VSS.n4349 0.147342
R11311 VSS.n4349 VSS.t147 3.13212
R11312 VSS.n4322 VSS.n4327 4.5005
R11313 VSS.n4324 VSS.n4328 4.5005
R11314 VSS.n4325 VSS.n4329 4.5005
R11315 VSS.n4326 VSS.n4330 4.57324
R11316 VSS.n4322 VSS.n4320 0.147342
R11317 VSS.n4323 VSS.n4324 0.0732424
R11318 VSS.n4324 VSS.n4325 0.147342
R11319 VSS.n4327 VSS.n4331 0.0721009
R11320 VSS.n4332 VSS.n4328 4.5005
R11321 VSS.n4333 VSS.n4329 4.5005
R11322 VSS.n4334 VSS.n4330 4.5005
R11323 VSS.n4320 VSS.n4331 4.57442
R11324 VSS.n4327 VSS.n4328 0.147342
R11325 VSS.n4328 VSS.n4329 0.147342
R11326 VSS.n4329 VSS.n4330 0.147342
R11327 VSS.n4331 VSS.n4332 2.39784
R11328 VSS.n4332 VSS.n4333 0.147342
R11329 VSS.n4333 VSS.n4334 0.147342
R11330 VSS.n4334 VSS.t10 3.13212
R11331 VSS.n4307 VSS.n4312 4.5005
R11332 VSS.n4309 VSS.n4313 4.5005
R11333 VSS.n4310 VSS.n4314 4.5005
R11334 VSS.n4311 VSS.n4315 4.57324
R11335 VSS.n4307 VSS.n4305 0.147342
R11336 VSS.n4308 VSS.n4309 0.0732424
R11337 VSS.n4309 VSS.n4310 0.147342
R11338 VSS.n4312 VSS.n4316 0.0721009
R11339 VSS.n4317 VSS.n4313 4.5005
R11340 VSS.n4318 VSS.n4314 4.5005
R11341 VSS.n4319 VSS.n4315 4.5005
R11342 VSS.n4305 VSS.n4316 4.57442
R11343 VSS.n4312 VSS.n4313 0.147342
R11344 VSS.n4313 VSS.n4314 0.147342
R11345 VSS.n4314 VSS.n4315 0.147342
R11346 VSS.n4316 VSS.n4317 2.39784
R11347 VSS.n4317 VSS.n4318 0.147342
R11348 VSS.n4318 VSS.n4319 0.147342
R11349 VSS.n4319 VSS.t196 3.13212
R11350 VSS.n4292 VSS.n4297 4.5005
R11351 VSS.n4294 VSS.n4298 4.5005
R11352 VSS.n4295 VSS.n4299 4.5005
R11353 VSS.n4296 VSS.n4300 4.57324
R11354 VSS.n4292 VSS.n4290 0.147342
R11355 VSS.n4293 VSS.n4294 0.0732424
R11356 VSS.n4294 VSS.n4295 0.147342
R11357 VSS.n4297 VSS.n4301 0.0721009
R11358 VSS.n4302 VSS.n4298 4.5005
R11359 VSS.n4303 VSS.n4299 4.5005
R11360 VSS.n4304 VSS.n4300 4.5005
R11361 VSS.n4290 VSS.n4301 4.57442
R11362 VSS.n4297 VSS.n4298 0.147342
R11363 VSS.n4298 VSS.n4299 0.147342
R11364 VSS.n4299 VSS.n4300 0.147342
R11365 VSS.n4301 VSS.n4302 2.39784
R11366 VSS.n4302 VSS.n4303 0.147342
R11367 VSS.n4303 VSS.n4304 0.147342
R11368 VSS.n4304 VSS.t170 3.13212
R11369 VSS.n4282 VSS.n4277 4.5005
R11370 VSS.n4283 VSS.n4279 4.5005
R11371 VSS.n4284 VSS.n4280 4.5005
R11372 VSS.n4285 VSS.n4281 4.57324
R11373 VSS.n4275 VSS.n4277 0.147342
R11374 VSS.n4278 VSS.n4279 0.0732424
R11375 VSS.n4279 VSS.n4280 0.147342
R11376 VSS.n4286 VSS.n4282 0.0722544
R11377 VSS.n4287 VSS.n4283 4.5005
R11378 VSS.n4288 VSS.n4284 4.5005
R11379 VSS.n4289 VSS.n4285 4.5005
R11380 VSS.n4286 VSS.n4275 4.57426
R11381 VSS.n4282 VSS.n4283 0.147342
R11382 VSS.n4283 VSS.n4284 0.147342
R11383 VSS.n4284 VSS.n4285 0.147342
R11384 VSS.n4287 VSS.n4286 2.37296
R11385 VSS.n4288 VSS.n4287 0.127318
R11386 VSS.n4289 VSS.n4288 0.127318
R11387 VSS.t5 VSS.n4289 2.73618
R11388 VSS.n4262 VSS.n4267 4.5005
R11389 VSS.n4264 VSS.n4268 4.5005
R11390 VSS.n4265 VSS.n4269 4.5005
R11391 VSS.n4266 VSS.n4270 4.57324
R11392 VSS.n4262 VSS.n4260 0.147342
R11393 VSS.n4263 VSS.n4264 0.0732424
R11394 VSS.n4264 VSS.n4265 0.147342
R11395 VSS.n4267 VSS.n4271 0.0721009
R11396 VSS.n4272 VSS.n4268 4.5005
R11397 VSS.n4273 VSS.n4269 4.5005
R11398 VSS.n4274 VSS.n4270 4.5005
R11399 VSS.n4260 VSS.n4271 4.57442
R11400 VSS.n4267 VSS.n4268 0.147342
R11401 VSS.n4268 VSS.n4269 0.147342
R11402 VSS.n4269 VSS.n4270 0.147342
R11403 VSS.n4271 VSS.n4272 2.39784
R11404 VSS.n4272 VSS.n4273 0.147342
R11405 VSS.n4273 VSS.n4274 0.147342
R11406 VSS.n4274 VSS.t362 3.13212
R11407 VSS.n4247 VSS.n4252 4.5005
R11408 VSS.n4249 VSS.n4253 4.5005
R11409 VSS.n4250 VSS.n4254 4.5005
R11410 VSS.n4251 VSS.n4255 4.57324
R11411 VSS.n4247 VSS.n4245 0.147342
R11412 VSS.n4248 VSS.n4249 0.0732424
R11413 VSS.n4249 VSS.n4250 0.147342
R11414 VSS.n4252 VSS.n4256 0.0721009
R11415 VSS.n4257 VSS.n4253 4.5005
R11416 VSS.n4258 VSS.n4254 4.5005
R11417 VSS.n4259 VSS.n4255 4.5005
R11418 VSS.n4245 VSS.n4256 4.57442
R11419 VSS.n4252 VSS.n4253 0.147342
R11420 VSS.n4253 VSS.n4254 0.147342
R11421 VSS.n4254 VSS.n4255 0.147342
R11422 VSS.n4256 VSS.n4257 2.39784
R11423 VSS.n4257 VSS.n4258 0.147342
R11424 VSS.n4258 VSS.n4259 0.147342
R11425 VSS.n4259 VSS.t127 3.13212
R11426 VSS.n4232 VSS.n4237 4.5005
R11427 VSS.n4234 VSS.n4238 4.5005
R11428 VSS.n4235 VSS.n4239 4.5005
R11429 VSS.n4236 VSS.n4240 4.57324
R11430 VSS.n4232 VSS.n4230 0.147342
R11431 VSS.n4233 VSS.n4234 0.0732424
R11432 VSS.n4234 VSS.n4235 0.147342
R11433 VSS.n4237 VSS.n4241 0.0721009
R11434 VSS.n4242 VSS.n4238 4.5005
R11435 VSS.n4243 VSS.n4239 4.5005
R11436 VSS.n4244 VSS.n4240 4.5005
R11437 VSS.n4230 VSS.n4241 4.57442
R11438 VSS.n4237 VSS.n4238 0.147342
R11439 VSS.n4238 VSS.n4239 0.147342
R11440 VSS.n4239 VSS.n4240 0.147342
R11441 VSS.n4241 VSS.n4242 2.39784
R11442 VSS.n4242 VSS.n4243 0.147342
R11443 VSS.n4243 VSS.n4244 0.147342
R11444 VSS.n4244 VSS.t16 3.13212
R11445 VSS.n4222 VSS.n4217 4.5005
R11446 VSS.n4223 VSS.n4219 4.5005
R11447 VSS.n4224 VSS.n4220 4.5005
R11448 VSS.n4225 VSS.n4221 4.57324
R11449 VSS.n4215 VSS.n4217 0.147342
R11450 VSS.n4218 VSS.n4219 0.0732424
R11451 VSS.n4219 VSS.n4220 0.147342
R11452 VSS.n4226 VSS.n4222 0.0722544
R11453 VSS.n4227 VSS.n4223 4.5005
R11454 VSS.n4228 VSS.n4224 4.5005
R11455 VSS.n4229 VSS.n4225 4.5005
R11456 VSS.n4226 VSS.n4215 4.57426
R11457 VSS.n4222 VSS.n4223 0.147342
R11458 VSS.n4223 VSS.n4224 0.147342
R11459 VSS.n4224 VSS.n4225 0.147342
R11460 VSS.n4227 VSS.n4226 2.37296
R11461 VSS.n4228 VSS.n4227 0.127318
R11462 VSS.n4229 VSS.n4228 0.127318
R11463 VSS.t5 VSS.n4229 2.73618
R11464 VSS.n4202 VSS.n4207 4.5005
R11465 VSS.n4204 VSS.n4208 4.5005
R11466 VSS.n4205 VSS.n4209 4.5005
R11467 VSS.n4206 VSS.n4210 4.57324
R11468 VSS.n4202 VSS.n4200 0.147342
R11469 VSS.n4203 VSS.n4204 0.0732424
R11470 VSS.n4204 VSS.n4205 0.147342
R11471 VSS.n4207 VSS.n4211 0.0721009
R11472 VSS.n4212 VSS.n4208 4.5005
R11473 VSS.n4213 VSS.n4209 4.5005
R11474 VSS.n4214 VSS.n4210 4.5005
R11475 VSS.n4200 VSS.n4211 4.57442
R11476 VSS.n4207 VSS.n4208 0.147342
R11477 VSS.n4208 VSS.n4209 0.147342
R11478 VSS.n4209 VSS.n4210 0.147342
R11479 VSS.n4211 VSS.n4212 2.39784
R11480 VSS.n4212 VSS.n4213 0.147342
R11481 VSS.n4213 VSS.n4214 0.147342
R11482 VSS.n4214 VSS.t331 3.13212
R11483 VSS.n4187 VSS.n4192 4.5005
R11484 VSS.n4189 VSS.n4193 4.5005
R11485 VSS.n4190 VSS.n4194 4.5005
R11486 VSS.n4191 VSS.n4195 4.57324
R11487 VSS.n4187 VSS.n4185 0.147342
R11488 VSS.n4188 VSS.n4189 0.0732424
R11489 VSS.n4189 VSS.n4190 0.147342
R11490 VSS.n4192 VSS.n4196 0.0721009
R11491 VSS.n4197 VSS.n4193 4.5005
R11492 VSS.n4198 VSS.n4194 4.5005
R11493 VSS.n4199 VSS.n4195 4.5005
R11494 VSS.n4185 VSS.n4196 4.57442
R11495 VSS.n4192 VSS.n4193 0.147342
R11496 VSS.n4193 VSS.n4194 0.147342
R11497 VSS.n4194 VSS.n4195 0.147342
R11498 VSS.n4196 VSS.n4197 2.39784
R11499 VSS.n4197 VSS.n4198 0.147342
R11500 VSS.n4198 VSS.n4199 0.147342
R11501 VSS.n4199 VSS.t259 3.13212
R11502 VSS.n4172 VSS.n4177 4.5005
R11503 VSS.n4174 VSS.n4178 4.5005
R11504 VSS.n4175 VSS.n4179 4.5005
R11505 VSS.n4176 VSS.n4180 4.57324
R11506 VSS.n4172 VSS.n4170 0.147342
R11507 VSS.n4173 VSS.n4174 0.0732424
R11508 VSS.n4174 VSS.n4175 0.147342
R11509 VSS.n4177 VSS.n4181 0.0721009
R11510 VSS.n4182 VSS.n4178 4.5005
R11511 VSS.n4183 VSS.n4179 4.5005
R11512 VSS.n4184 VSS.n4180 4.5005
R11513 VSS.n4170 VSS.n4181 4.57442
R11514 VSS.n4177 VSS.n4178 0.147342
R11515 VSS.n4178 VSS.n4179 0.147342
R11516 VSS.n4179 VSS.n4180 0.147342
R11517 VSS.n4181 VSS.n4182 2.39784
R11518 VSS.n4182 VSS.n4183 0.147342
R11519 VSS.n4183 VSS.n4184 0.147342
R11520 VSS.n4184 VSS.t244 3.13212
R11521 VSS.n4157 VSS.n4162 4.5005
R11522 VSS.n4159 VSS.n4163 4.5005
R11523 VSS.n4160 VSS.n4164 4.5005
R11524 VSS.n4161 VSS.n4165 4.57324
R11525 VSS.n4157 VSS.n4155 0.147342
R11526 VSS.n4158 VSS.n4159 0.0732424
R11527 VSS.n4159 VSS.n4160 0.147342
R11528 VSS.n4162 VSS.n4166 0.0721009
R11529 VSS.n4167 VSS.n4163 4.5005
R11530 VSS.n4168 VSS.n4164 4.5005
R11531 VSS.n4169 VSS.n4165 4.5005
R11532 VSS.n4155 VSS.n4166 4.57442
R11533 VSS.n4162 VSS.n4163 0.147342
R11534 VSS.n4163 VSS.n4164 0.147342
R11535 VSS.n4164 VSS.n4165 0.147342
R11536 VSS.n4166 VSS.n4167 2.39784
R11537 VSS.n4167 VSS.n4168 0.147342
R11538 VSS.n4168 VSS.n4169 0.147342
R11539 VSS.n4169 VSS.t254 3.13212
R11540 VSS.n4147 VSS.n4142 4.5005
R11541 VSS.n4148 VSS.n4144 4.5005
R11542 VSS.n4149 VSS.n4145 4.5005
R11543 VSS.n4150 VSS.n4146 4.57324
R11544 VSS.n4140 VSS.n4142 0.147342
R11545 VSS.n4143 VSS.n4144 0.0732424
R11546 VSS.n4144 VSS.n4145 0.147342
R11547 VSS.n4151 VSS.n4147 0.0722544
R11548 VSS.n4152 VSS.n4148 4.5005
R11549 VSS.n4153 VSS.n4149 4.5005
R11550 VSS.n4154 VSS.n4150 4.5005
R11551 VSS.n4151 VSS.n4140 4.57426
R11552 VSS.n4147 VSS.n4148 0.147342
R11553 VSS.n4148 VSS.n4149 0.147342
R11554 VSS.n4149 VSS.n4150 0.147342
R11555 VSS.n4152 VSS.n4151 2.37296
R11556 VSS.n4153 VSS.n4152 0.127318
R11557 VSS.n4154 VSS.n4153 0.127318
R11558 VSS.t5 VSS.n4154 2.73618
R11559 VSS.n4127 VSS.n4132 4.5005
R11560 VSS.n4129 VSS.n4133 4.5005
R11561 VSS.n4130 VSS.n4134 4.5005
R11562 VSS.n4131 VSS.n4135 4.57324
R11563 VSS.n4127 VSS.n4125 0.147342
R11564 VSS.n4128 VSS.n4129 0.0732424
R11565 VSS.n4129 VSS.n4130 0.147342
R11566 VSS.n4132 VSS.n4136 0.0721009
R11567 VSS.n4137 VSS.n4133 4.5005
R11568 VSS.n4138 VSS.n4134 4.5005
R11569 VSS.n4139 VSS.n4135 4.5005
R11570 VSS.n4125 VSS.n4136 4.57442
R11571 VSS.n4132 VSS.n4133 0.147342
R11572 VSS.n4133 VSS.n4134 0.147342
R11573 VSS.n4134 VSS.n4135 0.147342
R11574 VSS.n4136 VSS.n4137 2.39784
R11575 VSS.n4137 VSS.n4138 0.147342
R11576 VSS.n4138 VSS.n4139 0.147342
R11577 VSS.n4139 VSS.t298 3.13212
R11578 VSS.n4112 VSS.n4117 4.5005
R11579 VSS.n4114 VSS.n4118 4.5005
R11580 VSS.n4115 VSS.n4119 4.5005
R11581 VSS.n4116 VSS.n4120 4.57324
R11582 VSS.n4112 VSS.n4110 0.147342
R11583 VSS.n4113 VSS.n4114 0.0732424
R11584 VSS.n4114 VSS.n4115 0.147342
R11585 VSS.n4117 VSS.n4121 0.0721009
R11586 VSS.n4122 VSS.n4118 4.5005
R11587 VSS.n4123 VSS.n4119 4.5005
R11588 VSS.n4124 VSS.n4120 4.5005
R11589 VSS.n4110 VSS.n4121 4.57442
R11590 VSS.n4117 VSS.n4118 0.147342
R11591 VSS.n4118 VSS.n4119 0.147342
R11592 VSS.n4119 VSS.n4120 0.147342
R11593 VSS.n4121 VSS.n4122 2.39784
R11594 VSS.n4122 VSS.n4123 0.147342
R11595 VSS.n4123 VSS.n4124 0.147342
R11596 VSS.n4124 VSS.t88 3.13212
R11597 VSS.n4097 VSS.n4102 4.5005
R11598 VSS.n4099 VSS.n4103 4.5005
R11599 VSS.n4100 VSS.n4104 4.5005
R11600 VSS.n4101 VSS.n4105 4.57324
R11601 VSS.n4097 VSS.n4095 0.147342
R11602 VSS.n4098 VSS.n4099 0.0732424
R11603 VSS.n4099 VSS.n4100 0.147342
R11604 VSS.n4102 VSS.n4106 0.0721009
R11605 VSS.n4107 VSS.n4103 4.5005
R11606 VSS.n4108 VSS.n4104 4.5005
R11607 VSS.n4109 VSS.n4105 4.5005
R11608 VSS.n4095 VSS.n4106 4.57442
R11609 VSS.n4102 VSS.n4103 0.147342
R11610 VSS.n4103 VSS.n4104 0.147342
R11611 VSS.n4104 VSS.n4105 0.147342
R11612 VSS.n4106 VSS.n4107 2.39784
R11613 VSS.n4107 VSS.n4108 0.147342
R11614 VSS.n4108 VSS.n4109 0.147342
R11615 VSS.n4109 VSS.t519 3.13212
R11616 VSS.n4087 VSS.n4082 4.5005
R11617 VSS.n4088 VSS.n4084 4.5005
R11618 VSS.n4089 VSS.n4085 4.5005
R11619 VSS.n4090 VSS.n4086 4.57324
R11620 VSS.n4080 VSS.n4082 0.147342
R11621 VSS.n4083 VSS.n4084 0.0732424
R11622 VSS.n4084 VSS.n4085 0.147342
R11623 VSS.n4091 VSS.n4087 0.0722544
R11624 VSS.n4092 VSS.n4088 4.5005
R11625 VSS.n4093 VSS.n4089 4.5005
R11626 VSS.n4094 VSS.n4090 4.5005
R11627 VSS.n4091 VSS.n4080 4.57426
R11628 VSS.n4087 VSS.n4088 0.147342
R11629 VSS.n4088 VSS.n4089 0.147342
R11630 VSS.n4089 VSS.n4090 0.147342
R11631 VSS.n4092 VSS.n4091 2.37296
R11632 VSS.n4093 VSS.n4092 0.127318
R11633 VSS.n4094 VSS.n4093 0.127318
R11634 VSS.t5 VSS.n4094 2.73618
R11635 VSS.n4067 VSS.n4072 4.5005
R11636 VSS.n4069 VSS.n4073 4.5005
R11637 VSS.n4070 VSS.n4074 4.5005
R11638 VSS.n4071 VSS.n4075 4.57324
R11639 VSS.n4067 VSS.n4065 0.147342
R11640 VSS.n4068 VSS.n4069 0.0732424
R11641 VSS.n4069 VSS.n4070 0.147342
R11642 VSS.n4072 VSS.n4076 0.0721009
R11643 VSS.n4077 VSS.n4073 4.5005
R11644 VSS.n4078 VSS.n4074 4.5005
R11645 VSS.n4079 VSS.n4075 4.5005
R11646 VSS.n4065 VSS.n4076 4.57442
R11647 VSS.n4072 VSS.n4073 0.147342
R11648 VSS.n4073 VSS.n4074 0.147342
R11649 VSS.n4074 VSS.n4075 0.147342
R11650 VSS.n4076 VSS.n4077 2.39784
R11651 VSS.n4077 VSS.n4078 0.147342
R11652 VSS.n4078 VSS.n4079 0.147342
R11653 VSS.n4079 VSS.t71 3.13212
R11654 VSS.n4052 VSS.n4057 4.5005
R11655 VSS.n4054 VSS.n4058 4.5005
R11656 VSS.n4055 VSS.n4059 4.5005
R11657 VSS.n4056 VSS.n4060 4.57324
R11658 VSS.n4052 VSS.n4050 0.147342
R11659 VSS.n4053 VSS.n4054 0.0732424
R11660 VSS.n4054 VSS.n4055 0.147342
R11661 VSS.n4057 VSS.n4061 0.0721009
R11662 VSS.n4062 VSS.n4058 4.5005
R11663 VSS.n4063 VSS.n4059 4.5005
R11664 VSS.n4064 VSS.n4060 4.5005
R11665 VSS.n4050 VSS.n4061 4.57442
R11666 VSS.n4057 VSS.n4058 0.147342
R11667 VSS.n4058 VSS.n4059 0.147342
R11668 VSS.n4059 VSS.n4060 0.147342
R11669 VSS.n4061 VSS.n4062 2.39784
R11670 VSS.n4062 VSS.n4063 0.147342
R11671 VSS.n4063 VSS.n4064 0.147342
R11672 VSS.n4064 VSS.t186 3.13212
R11673 VSS.n4037 VSS.n4042 4.5005
R11674 VSS.n4039 VSS.n4043 4.5005
R11675 VSS.n4040 VSS.n4044 4.5005
R11676 VSS.n4041 VSS.n4045 4.57324
R11677 VSS.n4037 VSS.n4035 0.147342
R11678 VSS.n4038 VSS.n4039 0.0732424
R11679 VSS.n4039 VSS.n4040 0.147342
R11680 VSS.n4042 VSS.n4046 0.0721009
R11681 VSS.n4047 VSS.n4043 4.5005
R11682 VSS.n4048 VSS.n4044 4.5005
R11683 VSS.n4049 VSS.n4045 4.5005
R11684 VSS.n4035 VSS.n4046 4.57442
R11685 VSS.n4042 VSS.n4043 0.147342
R11686 VSS.n4043 VSS.n4044 0.147342
R11687 VSS.n4044 VSS.n4045 0.147342
R11688 VSS.n4046 VSS.n4047 2.39784
R11689 VSS.n4047 VSS.n4048 0.147342
R11690 VSS.n4048 VSS.n4049 0.147342
R11691 VSS.n4049 VSS.t108 3.13212
R11692 VSS.n4022 VSS.n4027 4.5005
R11693 VSS.n4024 VSS.n4028 4.5005
R11694 VSS.n4025 VSS.n4029 4.5005
R11695 VSS.n4026 VSS.n4030 4.57324
R11696 VSS.n4022 VSS.n4020 0.147342
R11697 VSS.n4023 VSS.n4024 0.0732424
R11698 VSS.n4024 VSS.n4025 0.147342
R11699 VSS.n4027 VSS.n4031 0.0721009
R11700 VSS.n4032 VSS.n4028 4.5005
R11701 VSS.n4033 VSS.n4029 4.5005
R11702 VSS.n4034 VSS.n4030 4.5005
R11703 VSS.n4020 VSS.n4031 4.57442
R11704 VSS.n4027 VSS.n4028 0.147342
R11705 VSS.n4028 VSS.n4029 0.147342
R11706 VSS.n4029 VSS.n4030 0.147342
R11707 VSS.n4031 VSS.n4032 2.39784
R11708 VSS.n4032 VSS.n4033 0.147342
R11709 VSS.n4033 VSS.n4034 0.147342
R11710 VSS.n4034 VSS.t12 3.13212
R11711 VSS.n4007 VSS.n4012 4.5005
R11712 VSS.n4009 VSS.n4013 4.5005
R11713 VSS.n4010 VSS.n4014 4.5005
R11714 VSS.n4011 VSS.n4015 4.57324
R11715 VSS.n4007 VSS.n4005 0.147342
R11716 VSS.n4008 VSS.n4009 0.0732424
R11717 VSS.n4009 VSS.n4010 0.147342
R11718 VSS.n4012 VSS.n4016 0.0721009
R11719 VSS.n4017 VSS.n4013 4.5005
R11720 VSS.n4018 VSS.n4014 4.5005
R11721 VSS.n4019 VSS.n4015 4.5005
R11722 VSS.n4005 VSS.n4016 4.57442
R11723 VSS.n4012 VSS.n4013 0.147342
R11724 VSS.n4013 VSS.n4014 0.147342
R11725 VSS.n4014 VSS.n4015 0.147342
R11726 VSS.n4016 VSS.n4017 2.39784
R11727 VSS.n4017 VSS.n4018 0.147342
R11728 VSS.n4018 VSS.n4019 0.147342
R11729 VSS.n4019 VSS.t194 3.13212
R11730 VSS.n3992 VSS.n3997 4.5005
R11731 VSS.n3994 VSS.n3998 4.5005
R11732 VSS.n3995 VSS.n3999 4.5005
R11733 VSS.n3996 VSS.n4000 4.57324
R11734 VSS.n3992 VSS.n3990 0.147342
R11735 VSS.n3993 VSS.n3994 0.0732424
R11736 VSS.n3994 VSS.n3995 0.147342
R11737 VSS.n3997 VSS.n4001 0.0721009
R11738 VSS.n4002 VSS.n3998 4.5005
R11739 VSS.n4003 VSS.n3999 4.5005
R11740 VSS.n4004 VSS.n4000 4.5005
R11741 VSS.n3990 VSS.n4001 4.57442
R11742 VSS.n3997 VSS.n3998 0.147342
R11743 VSS.n3998 VSS.n3999 0.147342
R11744 VSS.n3999 VSS.n4000 0.147342
R11745 VSS.n4001 VSS.n4002 2.39784
R11746 VSS.n4002 VSS.n4003 0.147342
R11747 VSS.n4003 VSS.n4004 0.147342
R11748 VSS.n4004 VSS.t168 3.13212
R11749 VSS.n3982 VSS.n3977 4.5005
R11750 VSS.n3983 VSS.n3979 4.5005
R11751 VSS.n3984 VSS.n3980 4.5005
R11752 VSS.n3985 VSS.n3981 4.57324
R11753 VSS.n3975 VSS.n3977 0.147342
R11754 VSS.n3978 VSS.n3979 0.0732424
R11755 VSS.n3979 VSS.n3980 0.147342
R11756 VSS.n3986 VSS.n3982 0.0722544
R11757 VSS.n3987 VSS.n3983 4.5005
R11758 VSS.n3988 VSS.n3984 4.5005
R11759 VSS.n3989 VSS.n3985 4.5005
R11760 VSS.n3986 VSS.n3975 4.57426
R11761 VSS.n3982 VSS.n3983 0.147342
R11762 VSS.n3983 VSS.n3984 0.147342
R11763 VSS.n3984 VSS.n3985 0.147342
R11764 VSS.n3987 VSS.n3986 2.37296
R11765 VSS.n3988 VSS.n3987 0.127318
R11766 VSS.n3989 VSS.n3988 0.127318
R11767 VSS.t5 VSS.n3989 2.73618
R11768 VSS.n3962 VSS.n3967 4.5005
R11769 VSS.n3964 VSS.n3968 4.5005
R11770 VSS.n3965 VSS.n3969 4.5005
R11771 VSS.n3966 VSS.n3970 4.57324
R11772 VSS.n3962 VSS.n3960 0.147342
R11773 VSS.n3963 VSS.n3964 0.0732424
R11774 VSS.n3964 VSS.n3965 0.147342
R11775 VSS.n3967 VSS.n3971 0.0721009
R11776 VSS.n3972 VSS.n3968 4.5005
R11777 VSS.n3973 VSS.n3969 4.5005
R11778 VSS.n3974 VSS.n3970 4.5005
R11779 VSS.n3960 VSS.n3971 4.57442
R11780 VSS.n3967 VSS.n3968 0.147342
R11781 VSS.n3968 VSS.n3969 0.147342
R11782 VSS.n3969 VSS.n3970 0.147342
R11783 VSS.n3971 VSS.n3972 2.39784
R11784 VSS.n3972 VSS.n3973 0.147342
R11785 VSS.n3973 VSS.n3974 0.147342
R11786 VSS.n3974 VSS.t364 3.13212
R11787 VSS.n3947 VSS.n3952 4.5005
R11788 VSS.n3949 VSS.n3953 4.5005
R11789 VSS.n3950 VSS.n3954 4.5005
R11790 VSS.n3951 VSS.n3955 4.57324
R11791 VSS.n3947 VSS.n3945 0.147342
R11792 VSS.n3948 VSS.n3949 0.0732424
R11793 VSS.n3949 VSS.n3950 0.147342
R11794 VSS.n3952 VSS.n3956 0.0721009
R11795 VSS.n3957 VSS.n3953 4.5005
R11796 VSS.n3958 VSS.n3954 4.5005
R11797 VSS.n3959 VSS.n3955 4.5005
R11798 VSS.n3945 VSS.n3956 4.57442
R11799 VSS.n3952 VSS.n3953 0.147342
R11800 VSS.n3953 VSS.n3954 0.147342
R11801 VSS.n3954 VSS.n3955 0.147342
R11802 VSS.n3956 VSS.n3957 2.39784
R11803 VSS.n3957 VSS.n3958 0.147342
R11804 VSS.n3958 VSS.n3959 0.147342
R11805 VSS.n3959 VSS.t325 3.13212
R11806 VSS.n3932 VSS.n3937 4.5005
R11807 VSS.n3934 VSS.n3938 4.5005
R11808 VSS.n3935 VSS.n3939 4.5005
R11809 VSS.n3936 VSS.n3940 4.57324
R11810 VSS.n3932 VSS.n3930 0.147342
R11811 VSS.n3933 VSS.n3934 0.0732424
R11812 VSS.n3934 VSS.n3935 0.147342
R11813 VSS.n3937 VSS.n3941 0.0721009
R11814 VSS.n3942 VSS.n3938 4.5005
R11815 VSS.n3943 VSS.n3939 4.5005
R11816 VSS.n3944 VSS.n3940 4.5005
R11817 VSS.n3930 VSS.n3941 4.57442
R11818 VSS.n3937 VSS.n3938 0.147342
R11819 VSS.n3938 VSS.n3939 0.147342
R11820 VSS.n3939 VSS.n3940 0.147342
R11821 VSS.n3941 VSS.n3942 2.39784
R11822 VSS.n3942 VSS.n3943 0.147342
R11823 VSS.n3943 VSS.n3944 0.147342
R11824 VSS.n3944 VSS.t18 3.13212
R11825 VSS.n3922 VSS.n3917 4.5005
R11826 VSS.n3923 VSS.n3919 4.5005
R11827 VSS.n3924 VSS.n3920 4.5005
R11828 VSS.n3925 VSS.n3921 4.57324
R11829 VSS.n3915 VSS.n3917 0.147342
R11830 VSS.n3918 VSS.n3919 0.0732424
R11831 VSS.n3919 VSS.n3920 0.147342
R11832 VSS.n3926 VSS.n3922 0.0722544
R11833 VSS.n3927 VSS.n3923 4.5005
R11834 VSS.n3928 VSS.n3924 4.5005
R11835 VSS.n3929 VSS.n3925 4.5005
R11836 VSS.n3926 VSS.n3915 4.57426
R11837 VSS.n3922 VSS.n3923 0.147342
R11838 VSS.n3923 VSS.n3924 0.147342
R11839 VSS.n3924 VSS.n3925 0.147342
R11840 VSS.n3927 VSS.n3926 2.37296
R11841 VSS.n3928 VSS.n3927 0.127318
R11842 VSS.n3929 VSS.n3928 0.127318
R11843 VSS.t5 VSS.n3929 2.73618
R11844 VSS.n3902 VSS.n3907 4.5005
R11845 VSS.n3904 VSS.n3908 4.5005
R11846 VSS.n3905 VSS.n3909 4.5005
R11847 VSS.n3906 VSS.n3910 4.57324
R11848 VSS.n3902 VSS.n3900 0.147342
R11849 VSS.n3903 VSS.n3904 0.0732424
R11850 VSS.n3904 VSS.n3905 0.147342
R11851 VSS.n3907 VSS.n3911 0.0721009
R11852 VSS.n3912 VSS.n3908 4.5005
R11853 VSS.n3913 VSS.n3909 4.5005
R11854 VSS.n3914 VSS.n3910 4.5005
R11855 VSS.n3900 VSS.n3911 4.57442
R11856 VSS.n3907 VSS.n3908 0.147342
R11857 VSS.n3908 VSS.n3909 0.147342
R11858 VSS.n3909 VSS.n3910 0.147342
R11859 VSS.n3911 VSS.n3912 2.39784
R11860 VSS.n3912 VSS.n3913 0.147342
R11861 VSS.n3913 VSS.n3914 0.147342
R11862 VSS.n3914 VSS.t229 3.13212
R11863 VSS.n3887 VSS.n3892 4.5005
R11864 VSS.n3889 VSS.n3893 4.5005
R11865 VSS.n3890 VSS.n3894 4.5005
R11866 VSS.n3891 VSS.n3895 4.57324
R11867 VSS.n3887 VSS.n3885 0.147342
R11868 VSS.n3888 VSS.n3889 0.0732424
R11869 VSS.n3889 VSS.n3890 0.147342
R11870 VSS.n3892 VSS.n3896 0.0721009
R11871 VSS.n3897 VSS.n3893 4.5005
R11872 VSS.n3898 VSS.n3894 4.5005
R11873 VSS.n3899 VSS.n3895 4.5005
R11874 VSS.n3885 VSS.n3896 4.57442
R11875 VSS.n3892 VSS.n3893 0.147342
R11876 VSS.n3893 VSS.n3894 0.147342
R11877 VSS.n3894 VSS.n3895 0.147342
R11878 VSS.n3896 VSS.n3897 2.39784
R11879 VSS.n3897 VSS.n3898 0.147342
R11880 VSS.n3898 VSS.n3899 0.147342
R11881 VSS.n3899 VSS.t491 3.13212
R11882 VSS.n3872 VSS.n3877 4.5005
R11883 VSS.n3874 VSS.n3878 4.5005
R11884 VSS.n3875 VSS.n3879 4.5005
R11885 VSS.n3876 VSS.n3880 4.57324
R11886 VSS.n3872 VSS.n3870 0.147342
R11887 VSS.n3873 VSS.n3874 0.0732424
R11888 VSS.n3874 VSS.n3875 0.147342
R11889 VSS.n3877 VSS.n3881 0.0721009
R11890 VSS.n3882 VSS.n3878 4.5005
R11891 VSS.n3883 VSS.n3879 4.5005
R11892 VSS.n3884 VSS.n3880 4.5005
R11893 VSS.n3870 VSS.n3881 4.57442
R11894 VSS.n3877 VSS.n3878 0.147342
R11895 VSS.n3878 VSS.n3879 0.147342
R11896 VSS.n3879 VSS.n3880 0.147342
R11897 VSS.n3881 VSS.n3882 2.39784
R11898 VSS.n3882 VSS.n3883 0.147342
R11899 VSS.n3883 VSS.n3884 0.147342
R11900 VSS.n3884 VSS.t242 3.13212
R11901 VSS.n3857 VSS.n3862 4.5005
R11902 VSS.n3859 VSS.n3863 4.5005
R11903 VSS.n3860 VSS.n3864 4.5005
R11904 VSS.n3861 VSS.n3865 4.57324
R11905 VSS.n3857 VSS.n3855 0.147342
R11906 VSS.n3858 VSS.n3859 0.0732424
R11907 VSS.n3859 VSS.n3860 0.147342
R11908 VSS.n3862 VSS.n3866 0.0721009
R11909 VSS.n3867 VSS.n3863 4.5005
R11910 VSS.n3868 VSS.n3864 4.5005
R11911 VSS.n3869 VSS.n3865 4.5005
R11912 VSS.n3855 VSS.n3866 4.57442
R11913 VSS.n3862 VSS.n3863 0.147342
R11914 VSS.n3863 VSS.n3864 0.147342
R11915 VSS.n3864 VSS.n3865 0.147342
R11916 VSS.n3866 VSS.n3867 2.39784
R11917 VSS.n3867 VSS.n3868 0.147342
R11918 VSS.n3868 VSS.n3869 0.147342
R11919 VSS.n3869 VSS.t346 3.13212
R11920 VSS.n3847 VSS.n3842 4.5005
R11921 VSS.n3848 VSS.n3844 4.5005
R11922 VSS.n3849 VSS.n3845 4.5005
R11923 VSS.n3850 VSS.n3846 4.57324
R11924 VSS.n3840 VSS.n3842 0.147342
R11925 VSS.n3843 VSS.n3844 0.0732424
R11926 VSS.n3844 VSS.n3845 0.147342
R11927 VSS.n3851 VSS.n3847 0.0722544
R11928 VSS.n3852 VSS.n3848 4.5005
R11929 VSS.n3853 VSS.n3849 4.5005
R11930 VSS.n3854 VSS.n3850 4.5005
R11931 VSS.n3851 VSS.n3840 4.57426
R11932 VSS.n3847 VSS.n3848 0.147342
R11933 VSS.n3848 VSS.n3849 0.147342
R11934 VSS.n3849 VSS.n3850 0.147342
R11935 VSS.n3852 VSS.n3851 2.37296
R11936 VSS.n3853 VSS.n3852 0.127318
R11937 VSS.n3854 VSS.n3853 0.127318
R11938 VSS.t5 VSS.n3854 2.73618
R11939 VSS.n3827 VSS.n3832 4.5005
R11940 VSS.n3829 VSS.n3833 4.5005
R11941 VSS.n3830 VSS.n3834 4.5005
R11942 VSS.n3831 VSS.n3835 4.57324
R11943 VSS.n3827 VSS.n3825 0.147342
R11944 VSS.n3828 VSS.n3829 0.0732424
R11945 VSS.n3829 VSS.n3830 0.147342
R11946 VSS.n3832 VSS.n3836 0.0721009
R11947 VSS.n3837 VSS.n3833 4.5005
R11948 VSS.n3838 VSS.n3834 4.5005
R11949 VSS.n3839 VSS.n3835 4.5005
R11950 VSS.n3825 VSS.n3836 4.57442
R11951 VSS.n3832 VSS.n3833 0.147342
R11952 VSS.n3833 VSS.n3834 0.147342
R11953 VSS.n3834 VSS.n3835 0.147342
R11954 VSS.n3836 VSS.n3837 2.39784
R11955 VSS.n3837 VSS.n3838 0.147342
R11956 VSS.n3838 VSS.n3839 0.147342
R11957 VSS.n3839 VSS.t427 3.13212
R11958 VSS.n3812 VSS.n3817 4.5005
R11959 VSS.n3814 VSS.n3818 4.5005
R11960 VSS.n3815 VSS.n3819 4.5005
R11961 VSS.n3816 VSS.n3820 4.57324
R11962 VSS.n3812 VSS.n3810 0.147342
R11963 VSS.n3813 VSS.n3814 0.0732424
R11964 VSS.n3814 VSS.n3815 0.147342
R11965 VSS.n3817 VSS.n3821 0.0721009
R11966 VSS.n3822 VSS.n3818 4.5005
R11967 VSS.n3823 VSS.n3819 4.5005
R11968 VSS.n3824 VSS.n3820 4.5005
R11969 VSS.n3810 VSS.n3821 4.57442
R11970 VSS.n3817 VSS.n3818 0.147342
R11971 VSS.n3818 VSS.n3819 0.147342
R11972 VSS.n3819 VSS.n3820 0.147342
R11973 VSS.n3821 VSS.n3822 2.39784
R11974 VSS.n3822 VSS.n3823 0.147342
R11975 VSS.n3823 VSS.n3824 0.147342
R11976 VSS.n3824 VSS.t90 3.13212
R11977 VSS.n3797 VSS.n3802 4.5005
R11978 VSS.n3799 VSS.n3803 4.5005
R11979 VSS.n3800 VSS.n3804 4.5005
R11980 VSS.n3801 VSS.n3805 4.57324
R11981 VSS.n3797 VSS.n3795 0.147342
R11982 VSS.n3798 VSS.n3799 0.0732424
R11983 VSS.n3799 VSS.n3800 0.147342
R11984 VSS.n3802 VSS.n3806 0.0721009
R11985 VSS.n3807 VSS.n3803 4.5005
R11986 VSS.n3808 VSS.n3804 4.5005
R11987 VSS.n3809 VSS.n3805 4.5005
R11988 VSS.n3795 VSS.n3806 4.57442
R11989 VSS.n3802 VSS.n3803 0.147342
R11990 VSS.n3803 VSS.n3804 0.147342
R11991 VSS.n3804 VSS.n3805 0.147342
R11992 VSS.n3806 VSS.n3807 2.39784
R11993 VSS.n3807 VSS.n3808 0.147342
R11994 VSS.n3808 VSS.n3809 0.147342
R11995 VSS.n3809 VSS.t119 3.13212
R11996 VSS.n3787 VSS.n3782 4.5005
R11997 VSS.n3788 VSS.n3784 4.5005
R11998 VSS.n3789 VSS.n3785 4.5005
R11999 VSS.n3790 VSS.n3786 4.57324
R12000 VSS.n3780 VSS.n3782 0.147342
R12001 VSS.n3783 VSS.n3784 0.0732424
R12002 VSS.n3784 VSS.n3785 0.147342
R12003 VSS.n3791 VSS.n3787 0.0722544
R12004 VSS.n3792 VSS.n3788 4.5005
R12005 VSS.n3793 VSS.n3789 4.5005
R12006 VSS.n3794 VSS.n3790 4.5005
R12007 VSS.n3791 VSS.n3780 4.57426
R12008 VSS.n3787 VSS.n3788 0.147342
R12009 VSS.n3788 VSS.n3789 0.147342
R12010 VSS.n3789 VSS.n3790 0.147342
R12011 VSS.n3792 VSS.n3791 2.37296
R12012 VSS.n3793 VSS.n3792 0.127318
R12013 VSS.n3794 VSS.n3793 0.127318
R12014 VSS.t5 VSS.n3794 2.73618
R12015 VSS.n3767 VSS.n3772 4.5005
R12016 VSS.n3769 VSS.n3773 4.5005
R12017 VSS.n3770 VSS.n3774 4.5005
R12018 VSS.n3771 VSS.n3775 4.57324
R12019 VSS.n3767 VSS.n3765 0.147342
R12020 VSS.n3768 VSS.n3769 0.0732424
R12021 VSS.n3769 VSS.n3770 0.147342
R12022 VSS.n3772 VSS.n3776 0.0721009
R12023 VSS.n3777 VSS.n3773 4.5005
R12024 VSS.n3778 VSS.n3774 4.5005
R12025 VSS.n3779 VSS.n3775 4.5005
R12026 VSS.n3765 VSS.n3776 4.57442
R12027 VSS.n3772 VSS.n3773 0.147342
R12028 VSS.n3773 VSS.n3774 0.147342
R12029 VSS.n3774 VSS.n3775 0.147342
R12030 VSS.n3776 VSS.n3777 2.39784
R12031 VSS.n3777 VSS.n3778 0.147342
R12032 VSS.n3778 VSS.n3779 0.147342
R12033 VSS.n3779 VSS.t75 3.13212
R12034 VSS.n3752 VSS.n3757 4.5005
R12035 VSS.n3754 VSS.n3758 4.5005
R12036 VSS.n3755 VSS.n3759 4.5005
R12037 VSS.n3756 VSS.n3760 4.57324
R12038 VSS.n3752 VSS.n3750 0.147342
R12039 VSS.n3753 VSS.n3754 0.0732424
R12040 VSS.n3754 VSS.n3755 0.147342
R12041 VSS.n3757 VSS.n3761 0.0721009
R12042 VSS.n3762 VSS.n3758 4.5005
R12043 VSS.n3763 VSS.n3759 4.5005
R12044 VSS.n3764 VSS.n3760 4.5005
R12045 VSS.n3750 VSS.n3761 4.57442
R12046 VSS.n3757 VSS.n3758 0.147342
R12047 VSS.n3758 VSS.n3759 0.147342
R12048 VSS.n3759 VSS.n3760 0.147342
R12049 VSS.n3761 VSS.n3762 2.39784
R12050 VSS.n3762 VSS.n3763 0.147342
R12051 VSS.n3763 VSS.n3764 0.147342
R12052 VSS.n3764 VSS.t187 3.13212
R12053 VSS.n3737 VSS.n3742 4.5005
R12054 VSS.n3739 VSS.n3743 4.5005
R12055 VSS.n3740 VSS.n3744 4.5005
R12056 VSS.n3741 VSS.n3745 4.57324
R12057 VSS.n3737 VSS.n3735 0.147342
R12058 VSS.n3738 VSS.n3739 0.0732424
R12059 VSS.n3739 VSS.n3740 0.147342
R12060 VSS.n3742 VSS.n3746 0.0721009
R12061 VSS.n3747 VSS.n3743 4.5005
R12062 VSS.n3748 VSS.n3744 4.5005
R12063 VSS.n3749 VSS.n3745 4.5005
R12064 VSS.n3735 VSS.n3746 4.57442
R12065 VSS.n3742 VSS.n3743 0.147342
R12066 VSS.n3743 VSS.n3744 0.147342
R12067 VSS.n3744 VSS.n3745 0.147342
R12068 VSS.n3746 VSS.n3747 2.39784
R12069 VSS.n3747 VSS.n3748 0.147342
R12070 VSS.n3748 VSS.n3749 0.147342
R12071 VSS.n3749 VSS.t109 3.13212
R12072 VSS.n3722 VSS.n3727 4.5005
R12073 VSS.n3724 VSS.n3728 4.5005
R12074 VSS.n3725 VSS.n3729 4.5005
R12075 VSS.n3726 VSS.n3730 4.57324
R12076 VSS.n3722 VSS.n3720 0.147342
R12077 VSS.n3723 VSS.n3724 0.0732424
R12078 VSS.n3724 VSS.n3725 0.147342
R12079 VSS.n3727 VSS.n3731 0.0721009
R12080 VSS.n3732 VSS.n3728 4.5005
R12081 VSS.n3733 VSS.n3729 4.5005
R12082 VSS.n3734 VSS.n3730 4.5005
R12083 VSS.n3720 VSS.n3731 4.57442
R12084 VSS.n3727 VSS.n3728 0.147342
R12085 VSS.n3728 VSS.n3729 0.147342
R12086 VSS.n3729 VSS.n3730 0.147342
R12087 VSS.n3731 VSS.n3732 2.39784
R12088 VSS.n3732 VSS.n3733 0.147342
R12089 VSS.n3733 VSS.n3734 0.147342
R12090 VSS.n3734 VSS.t7 3.13212
R12091 VSS.n3707 VSS.n3712 4.5005
R12092 VSS.n3709 VSS.n3713 4.5005
R12093 VSS.n3710 VSS.n3714 4.5005
R12094 VSS.n3711 VSS.n3715 4.57324
R12095 VSS.n3707 VSS.n3705 0.147342
R12096 VSS.n3708 VSS.n3709 0.0732424
R12097 VSS.n3709 VSS.n3710 0.147342
R12098 VSS.n3712 VSS.n3716 0.0721009
R12099 VSS.n3717 VSS.n3713 4.5005
R12100 VSS.n3718 VSS.n3714 4.5005
R12101 VSS.n3719 VSS.n3715 4.5005
R12102 VSS.n3705 VSS.n3716 4.57442
R12103 VSS.n3712 VSS.n3713 0.147342
R12104 VSS.n3713 VSS.n3714 0.147342
R12105 VSS.n3714 VSS.n3715 0.147342
R12106 VSS.n3716 VSS.n3717 2.39784
R12107 VSS.n3717 VSS.n3718 0.147342
R12108 VSS.n3718 VSS.n3719 0.147342
R12109 VSS.n3719 VSS.t191 3.13212
R12110 VSS.n3692 VSS.n3697 4.5005
R12111 VSS.n3694 VSS.n3698 4.5005
R12112 VSS.n3695 VSS.n3699 4.5005
R12113 VSS.n3696 VSS.n3700 4.57324
R12114 VSS.n3692 VSS.n3690 0.147342
R12115 VSS.n3693 VSS.n3694 0.0732424
R12116 VSS.n3694 VSS.n3695 0.147342
R12117 VSS.n3697 VSS.n3701 0.0721009
R12118 VSS.n3702 VSS.n3698 4.5005
R12119 VSS.n3703 VSS.n3699 4.5005
R12120 VSS.n3704 VSS.n3700 4.5005
R12121 VSS.n3690 VSS.n3701 4.57442
R12122 VSS.n3697 VSS.n3698 0.147342
R12123 VSS.n3698 VSS.n3699 0.147342
R12124 VSS.n3699 VSS.n3700 0.147342
R12125 VSS.n3701 VSS.n3702 2.39784
R12126 VSS.n3702 VSS.n3703 0.147342
R12127 VSS.n3703 VSS.n3704 0.147342
R12128 VSS.n3704 VSS.t496 3.13212
R12129 VSS.n3682 VSS.n3677 4.5005
R12130 VSS.n3683 VSS.n3679 4.5005
R12131 VSS.n3684 VSS.n3680 4.5005
R12132 VSS.n3685 VSS.n3681 4.57324
R12133 VSS.n3675 VSS.n3677 0.147342
R12134 VSS.n3678 VSS.n3679 0.0732424
R12135 VSS.n3679 VSS.n3680 0.147342
R12136 VSS.n3686 VSS.n3682 0.0722544
R12137 VSS.n3687 VSS.n3683 4.5005
R12138 VSS.n3688 VSS.n3684 4.5005
R12139 VSS.n3689 VSS.n3685 4.5005
R12140 VSS.n3686 VSS.n3675 4.57426
R12141 VSS.n3682 VSS.n3683 0.147342
R12142 VSS.n3683 VSS.n3684 0.147342
R12143 VSS.n3684 VSS.n3685 0.147342
R12144 VSS.n3687 VSS.n3686 2.37296
R12145 VSS.n3688 VSS.n3687 0.127318
R12146 VSS.n3689 VSS.n3688 0.127318
R12147 VSS.t5 VSS.n3689 2.73618
R12148 VSS.n3662 VSS.n3667 4.5005
R12149 VSS.n3664 VSS.n3668 4.5005
R12150 VSS.n3665 VSS.n3669 4.5005
R12151 VSS.n3666 VSS.n3670 4.57324
R12152 VSS.n3662 VSS.n3660 0.147342
R12153 VSS.n3663 VSS.n3664 0.0732424
R12154 VSS.n3664 VSS.n3665 0.147342
R12155 VSS.n3667 VSS.n3671 0.0721009
R12156 VSS.n3672 VSS.n3668 4.5005
R12157 VSS.n3673 VSS.n3669 4.5005
R12158 VSS.n3674 VSS.n3670 4.5005
R12159 VSS.n3660 VSS.n3671 4.57442
R12160 VSS.n3667 VSS.n3668 0.147342
R12161 VSS.n3668 VSS.n3669 0.147342
R12162 VSS.n3669 VSS.n3670 0.147342
R12163 VSS.n3671 VSS.n3672 2.39784
R12164 VSS.n3672 VSS.n3673 0.147342
R12165 VSS.n3673 VSS.n3674 0.147342
R12166 VSS.n3674 VSS.t348 3.13212
R12167 VSS.n3647 VSS.n3652 4.5005
R12168 VSS.n3649 VSS.n3653 4.5005
R12169 VSS.n3650 VSS.n3654 4.5005
R12170 VSS.n3651 VSS.n3655 4.57324
R12171 VSS.n3647 VSS.n3645 0.147342
R12172 VSS.n3648 VSS.n3649 0.0732424
R12173 VSS.n3649 VSS.n3650 0.147342
R12174 VSS.n3652 VSS.n3656 0.0721009
R12175 VSS.n3657 VSS.n3653 4.5005
R12176 VSS.n3658 VSS.n3654 4.5005
R12177 VSS.n3659 VSS.n3655 4.5005
R12178 VSS.n3645 VSS.n3656 4.57442
R12179 VSS.n3652 VSS.n3653 0.147342
R12180 VSS.n3653 VSS.n3654 0.147342
R12181 VSS.n3654 VSS.n3655 0.147342
R12182 VSS.n3656 VSS.n3657 2.39784
R12183 VSS.n3657 VSS.n3658 0.147342
R12184 VSS.n3658 VSS.n3659 0.147342
R12185 VSS.n3659 VSS.t326 3.13212
R12186 VSS.n3632 VSS.n3637 4.5005
R12187 VSS.n3634 VSS.n3638 4.5005
R12188 VSS.n3635 VSS.n3639 4.5005
R12189 VSS.n3636 VSS.n3640 4.57324
R12190 VSS.n3632 VSS.n3630 0.147342
R12191 VSS.n3633 VSS.n3634 0.0732424
R12192 VSS.n3634 VSS.n3635 0.147342
R12193 VSS.n3637 VSS.n3641 0.0721009
R12194 VSS.n3642 VSS.n3638 4.5005
R12195 VSS.n3643 VSS.n3639 4.5005
R12196 VSS.n3644 VSS.n3640 4.5005
R12197 VSS.n3630 VSS.n3641 4.57442
R12198 VSS.n3637 VSS.n3638 0.147342
R12199 VSS.n3638 VSS.n3639 0.147342
R12200 VSS.n3639 VSS.n3640 0.147342
R12201 VSS.n3641 VSS.n3642 2.39784
R12202 VSS.n3642 VSS.n3643 0.147342
R12203 VSS.n3643 VSS.n3644 0.147342
R12204 VSS.n3644 VSS.t30 3.13212
R12205 VSS.n3622 VSS.n3617 4.5005
R12206 VSS.n3623 VSS.n3619 4.5005
R12207 VSS.n3624 VSS.n3620 4.5005
R12208 VSS.n3625 VSS.n3621 4.57324
R12209 VSS.n3615 VSS.n3617 0.147342
R12210 VSS.n3618 VSS.n3619 0.0732424
R12211 VSS.n3619 VSS.n3620 0.147342
R12212 VSS.n3626 VSS.n3622 0.0722544
R12213 VSS.n3627 VSS.n3623 4.5005
R12214 VSS.n3628 VSS.n3624 4.5005
R12215 VSS.n3629 VSS.n3625 4.5005
R12216 VSS.n3626 VSS.n3615 4.57426
R12217 VSS.n3622 VSS.n3623 0.147342
R12218 VSS.n3623 VSS.n3624 0.147342
R12219 VSS.n3624 VSS.n3625 0.147342
R12220 VSS.n3627 VSS.n3626 2.37296
R12221 VSS.n3628 VSS.n3627 0.127318
R12222 VSS.n3629 VSS.n3628 0.127318
R12223 VSS.t5 VSS.n3629 2.73618
R12224 VSS.n3602 VSS.n3607 4.5005
R12225 VSS.n3604 VSS.n3608 4.5005
R12226 VSS.n3605 VSS.n3609 4.5005
R12227 VSS.n3606 VSS.n3610 4.57324
R12228 VSS.n3602 VSS.n3600 0.147342
R12229 VSS.n3603 VSS.n3604 0.0732424
R12230 VSS.n3604 VSS.n3605 0.147342
R12231 VSS.n3607 VSS.n3611 0.0721009
R12232 VSS.n3612 VSS.n3608 4.5005
R12233 VSS.n3613 VSS.n3609 4.5005
R12234 VSS.n3614 VSS.n3610 4.5005
R12235 VSS.n3600 VSS.n3611 4.57442
R12236 VSS.n3607 VSS.n3608 0.147342
R12237 VSS.n3608 VSS.n3609 0.147342
R12238 VSS.n3609 VSS.n3610 0.147342
R12239 VSS.n3611 VSS.n3612 2.39784
R12240 VSS.n3612 VSS.n3613 0.147342
R12241 VSS.n3613 VSS.n3614 0.147342
R12242 VSS.n3614 VSS.t233 3.13212
R12243 VSS.n3587 VSS.n3592 4.5005
R12244 VSS.n3589 VSS.n3593 4.5005
R12245 VSS.n3590 VSS.n3594 4.5005
R12246 VSS.n3591 VSS.n3595 4.57324
R12247 VSS.n3587 VSS.n3585 0.147342
R12248 VSS.n3588 VSS.n3589 0.0732424
R12249 VSS.n3589 VSS.n3590 0.147342
R12250 VSS.n3592 VSS.n3596 0.0721009
R12251 VSS.n3597 VSS.n3593 4.5005
R12252 VSS.n3598 VSS.n3594 4.5005
R12253 VSS.n3599 VSS.n3595 4.5005
R12254 VSS.n3585 VSS.n3596 4.57442
R12255 VSS.n3592 VSS.n3593 0.147342
R12256 VSS.n3593 VSS.n3594 0.147342
R12257 VSS.n3594 VSS.n3595 0.147342
R12258 VSS.n3596 VSS.n3597 2.39784
R12259 VSS.n3597 VSS.n3598 0.147342
R12260 VSS.n3598 VSS.n3599 0.147342
R12261 VSS.n3599 VSS.t468 3.13212
R12262 VSS.n3572 VSS.n3577 4.5005
R12263 VSS.n3574 VSS.n3578 4.5005
R12264 VSS.n3575 VSS.n3579 4.5005
R12265 VSS.n3576 VSS.n3580 4.57324
R12266 VSS.n3572 VSS.n3570 0.147342
R12267 VSS.n3573 VSS.n3574 0.0732424
R12268 VSS.n3574 VSS.n3575 0.147342
R12269 VSS.n3577 VSS.n3581 0.0721009
R12270 VSS.n3582 VSS.n3578 4.5005
R12271 VSS.n3583 VSS.n3579 4.5005
R12272 VSS.n3584 VSS.n3580 4.5005
R12273 VSS.n3570 VSS.n3581 4.57442
R12274 VSS.n3577 VSS.n3578 0.147342
R12275 VSS.n3578 VSS.n3579 0.147342
R12276 VSS.n3579 VSS.n3580 0.147342
R12277 VSS.n3581 VSS.n3582 2.39784
R12278 VSS.n3582 VSS.n3583 0.147342
R12279 VSS.n3583 VSS.n3584 0.147342
R12280 VSS.n3584 VSS.t245 3.13212
R12281 VSS.n3557 VSS.n3562 4.5005
R12282 VSS.n3559 VSS.n3563 4.5005
R12283 VSS.n3560 VSS.n3564 4.5005
R12284 VSS.n3561 VSS.n3565 4.57324
R12285 VSS.n3557 VSS.n3555 0.147342
R12286 VSS.n3558 VSS.n3559 0.0732424
R12287 VSS.n3559 VSS.n3560 0.147342
R12288 VSS.n3562 VSS.n3566 0.0721009
R12289 VSS.n3567 VSS.n3563 4.5005
R12290 VSS.n3568 VSS.n3564 4.5005
R12291 VSS.n3569 VSS.n3565 4.5005
R12292 VSS.n3555 VSS.n3566 4.57442
R12293 VSS.n3562 VSS.n3563 0.147342
R12294 VSS.n3563 VSS.n3564 0.147342
R12295 VSS.n3564 VSS.n3565 0.147342
R12296 VSS.n3566 VSS.n3567 2.39784
R12297 VSS.n3567 VSS.n3568 0.147342
R12298 VSS.n3568 VSS.n3569 0.147342
R12299 VSS.n3569 VSS.t249 3.13212
R12300 VSS.n3547 VSS.n3542 4.5005
R12301 VSS.n3548 VSS.n3544 4.5005
R12302 VSS.n3549 VSS.n3545 4.5005
R12303 VSS.n3550 VSS.n3546 4.57324
R12304 VSS.n3540 VSS.n3542 0.147342
R12305 VSS.n3543 VSS.n3544 0.0732424
R12306 VSS.n3544 VSS.n3545 0.147342
R12307 VSS.n3551 VSS.n3547 0.0722544
R12308 VSS.n3552 VSS.n3548 4.5005
R12309 VSS.n3553 VSS.n3549 4.5005
R12310 VSS.n3554 VSS.n3550 4.5005
R12311 VSS.n3551 VSS.n3540 4.57426
R12312 VSS.n3547 VSS.n3548 0.147342
R12313 VSS.n3548 VSS.n3549 0.147342
R12314 VSS.n3549 VSS.n3550 0.147342
R12315 VSS.n3552 VSS.n3551 2.37296
R12316 VSS.n3553 VSS.n3552 0.127318
R12317 VSS.n3554 VSS.n3553 0.127318
R12318 VSS.t5 VSS.n3554 2.73618
R12319 VSS.n3527 VSS.n3532 4.5005
R12320 VSS.n3529 VSS.n3533 4.5005
R12321 VSS.n3530 VSS.n3534 4.5005
R12322 VSS.n3531 VSS.n3535 4.57324
R12323 VSS.n3527 VSS.n3525 0.147342
R12324 VSS.n3528 VSS.n3529 0.0732424
R12325 VSS.n3529 VSS.n3530 0.147342
R12326 VSS.n3532 VSS.n3536 0.0721009
R12327 VSS.n3537 VSS.n3533 4.5005
R12328 VSS.n3538 VSS.n3534 4.5005
R12329 VSS.n3539 VSS.n3535 4.5005
R12330 VSS.n3525 VSS.n3536 4.57442
R12331 VSS.n3532 VSS.n3533 0.147342
R12332 VSS.n3533 VSS.n3534 0.147342
R12333 VSS.n3534 VSS.n3535 0.147342
R12334 VSS.n3536 VSS.n3537 2.39784
R12335 VSS.n3537 VSS.n3538 0.147342
R12336 VSS.n3538 VSS.n3539 0.147342
R12337 VSS.n3539 VSS.t414 3.13212
R12338 VSS.n3512 VSS.n3517 4.5005
R12339 VSS.n3514 VSS.n3518 4.5005
R12340 VSS.n3515 VSS.n3519 4.5005
R12341 VSS.n3516 VSS.n3520 4.57324
R12342 VSS.n3512 VSS.n3510 0.147342
R12343 VSS.n3513 VSS.n3514 0.0732424
R12344 VSS.n3514 VSS.n3515 0.147342
R12345 VSS.n3517 VSS.n3521 0.0721009
R12346 VSS.n3522 VSS.n3518 4.5005
R12347 VSS.n3523 VSS.n3519 4.5005
R12348 VSS.n3524 VSS.n3520 4.5005
R12349 VSS.n3510 VSS.n3521 4.57442
R12350 VSS.n3517 VSS.n3518 0.147342
R12351 VSS.n3518 VSS.n3519 0.147342
R12352 VSS.n3519 VSS.n3520 0.147342
R12353 VSS.n3521 VSS.n3522 2.39784
R12354 VSS.n3522 VSS.n3523 0.147342
R12355 VSS.n3523 VSS.n3524 0.147342
R12356 VSS.n3524 VSS.t86 3.13212
R12357 VSS.n3497 VSS.n3502 4.5005
R12358 VSS.n3499 VSS.n3503 4.5005
R12359 VSS.n3500 VSS.n3504 4.5005
R12360 VSS.n3501 VSS.n3505 4.57324
R12361 VSS.n3497 VSS.n3495 0.147342
R12362 VSS.n3498 VSS.n3499 0.0732424
R12363 VSS.n3499 VSS.n3500 0.147342
R12364 VSS.n3502 VSS.n3506 0.0721009
R12365 VSS.n3507 VSS.n3503 4.5005
R12366 VSS.n3508 VSS.n3504 4.5005
R12367 VSS.n3509 VSS.n3505 4.5005
R12368 VSS.n3495 VSS.n3506 4.57442
R12369 VSS.n3502 VSS.n3503 0.147342
R12370 VSS.n3503 VSS.n3504 0.147342
R12371 VSS.n3504 VSS.n3505 0.147342
R12372 VSS.n3506 VSS.n3507 2.39784
R12373 VSS.n3507 VSS.n3508 0.147342
R12374 VSS.n3508 VSS.n3509 0.147342
R12375 VSS.n3509 VSS.t120 3.13212
R12376 VSS.n3487 VSS.n3482 4.5005
R12377 VSS.n3488 VSS.n3484 4.5005
R12378 VSS.n3489 VSS.n3485 4.5005
R12379 VSS.n3490 VSS.n3486 4.57324
R12380 VSS.n3480 VSS.n3482 0.147342
R12381 VSS.n3483 VSS.n3484 0.0732424
R12382 VSS.n3484 VSS.n3485 0.147342
R12383 VSS.n3491 VSS.n3487 0.0722544
R12384 VSS.n3492 VSS.n3488 4.5005
R12385 VSS.n3493 VSS.n3489 4.5005
R12386 VSS.n3494 VSS.n3490 4.5005
R12387 VSS.n3491 VSS.n3480 4.57426
R12388 VSS.n3487 VSS.n3488 0.147342
R12389 VSS.n3488 VSS.n3489 0.147342
R12390 VSS.n3489 VSS.n3490 0.147342
R12391 VSS.n3492 VSS.n3491 2.37296
R12392 VSS.n3493 VSS.n3492 0.127318
R12393 VSS.n3494 VSS.n3493 0.127318
R12394 VSS.t5 VSS.n3494 2.73618
R12395 VSS.n3467 VSS.n3472 4.5005
R12396 VSS.n3469 VSS.n3473 4.5005
R12397 VSS.n3470 VSS.n3474 4.5005
R12398 VSS.n3471 VSS.n3475 4.57324
R12399 VSS.n3467 VSS.n3465 0.147342
R12400 VSS.n3468 VSS.n3469 0.0732424
R12401 VSS.n3469 VSS.n3470 0.147342
R12402 VSS.n3472 VSS.n3476 0.0721009
R12403 VSS.n3477 VSS.n3473 4.5005
R12404 VSS.n3478 VSS.n3474 4.5005
R12405 VSS.n3479 VSS.n3475 4.5005
R12406 VSS.n3465 VSS.n3476 4.57442
R12407 VSS.n3472 VSS.n3473 0.147342
R12408 VSS.n3473 VSS.n3474 0.147342
R12409 VSS.n3474 VSS.n3475 0.147342
R12410 VSS.n3476 VSS.n3477 2.39784
R12411 VSS.n3477 VSS.n3478 0.147342
R12412 VSS.n3478 VSS.n3479 0.147342
R12413 VSS.n3479 VSS.t70 3.13212
R12414 VSS.n3452 VSS.n3457 4.5005
R12415 VSS.n3454 VSS.n3458 4.5005
R12416 VSS.n3455 VSS.n3459 4.5005
R12417 VSS.n3456 VSS.n3460 4.57324
R12418 VSS.n3452 VSS.n3450 0.147342
R12419 VSS.n3453 VSS.n3454 0.0732424
R12420 VSS.n3454 VSS.n3455 0.147342
R12421 VSS.n3457 VSS.n3461 0.0721009
R12422 VSS.n3462 VSS.n3458 4.5005
R12423 VSS.n3463 VSS.n3459 4.5005
R12424 VSS.n3464 VSS.n3460 4.5005
R12425 VSS.n3450 VSS.n3461 4.57442
R12426 VSS.n3457 VSS.n3458 0.147342
R12427 VSS.n3458 VSS.n3459 0.147342
R12428 VSS.n3459 VSS.n3460 0.147342
R12429 VSS.n3461 VSS.n3462 2.39784
R12430 VSS.n3462 VSS.n3463 0.147342
R12431 VSS.n3463 VSS.n3464 0.147342
R12432 VSS.n3464 VSS.t188 3.13212
R12433 VSS.n3437 VSS.n3442 4.5005
R12434 VSS.n3439 VSS.n3443 4.5005
R12435 VSS.n3440 VSS.n3444 4.5005
R12436 VSS.n3441 VSS.n3445 4.57324
R12437 VSS.n3437 VSS.n3435 0.147342
R12438 VSS.n3438 VSS.n3439 0.0732424
R12439 VSS.n3439 VSS.n3440 0.147342
R12440 VSS.n3442 VSS.n3446 0.0721009
R12441 VSS.n3447 VSS.n3443 4.5005
R12442 VSS.n3448 VSS.n3444 4.5005
R12443 VSS.n3449 VSS.n3445 4.5005
R12444 VSS.n3435 VSS.n3446 4.57442
R12445 VSS.n3442 VSS.n3443 0.147342
R12446 VSS.n3443 VSS.n3444 0.147342
R12447 VSS.n3444 VSS.n3445 0.147342
R12448 VSS.n3446 VSS.n3447 2.39784
R12449 VSS.n3447 VSS.n3448 0.147342
R12450 VSS.n3448 VSS.n3449 0.147342
R12451 VSS.n3449 VSS.t146 3.13212
R12452 VSS.n3422 VSS.n3427 4.5005
R12453 VSS.n3424 VSS.n3428 4.5005
R12454 VSS.n3425 VSS.n3429 4.5005
R12455 VSS.n3426 VSS.n3430 4.57324
R12456 VSS.n3422 VSS.n3420 0.147342
R12457 VSS.n3423 VSS.n3424 0.0732424
R12458 VSS.n3424 VSS.n3425 0.147342
R12459 VSS.n3427 VSS.n3431 0.0721009
R12460 VSS.n3432 VSS.n3428 4.5005
R12461 VSS.n3433 VSS.n3429 4.5005
R12462 VSS.n3434 VSS.n3430 4.5005
R12463 VSS.n3420 VSS.n3431 4.57442
R12464 VSS.n3427 VSS.n3428 0.147342
R12465 VSS.n3428 VSS.n3429 0.147342
R12466 VSS.n3429 VSS.n3430 0.147342
R12467 VSS.n3431 VSS.n3432 2.39784
R12468 VSS.n3432 VSS.n3433 0.147342
R12469 VSS.n3433 VSS.n3434 0.147342
R12470 VSS.n3434 VSS.t8 3.13212
R12471 VSS.n3407 VSS.n3412 4.5005
R12472 VSS.n3409 VSS.n3413 4.5005
R12473 VSS.n3410 VSS.n3414 4.5005
R12474 VSS.n3411 VSS.n3415 4.57324
R12475 VSS.n3407 VSS.n3405 0.147342
R12476 VSS.n3408 VSS.n3409 0.0732424
R12477 VSS.n3409 VSS.n3410 0.147342
R12478 VSS.n3412 VSS.n3416 0.0721009
R12479 VSS.n3417 VSS.n3413 4.5005
R12480 VSS.n3418 VSS.n3414 4.5005
R12481 VSS.n3419 VSS.n3415 4.5005
R12482 VSS.n3405 VSS.n3416 4.57442
R12483 VSS.n3412 VSS.n3413 0.147342
R12484 VSS.n3413 VSS.n3414 0.147342
R12485 VSS.n3414 VSS.n3415 0.147342
R12486 VSS.n3416 VSS.n3417 2.39784
R12487 VSS.n3417 VSS.n3418 0.147342
R12488 VSS.n3418 VSS.n3419 0.147342
R12489 VSS.n3419 VSS.t192 3.13212
R12490 VSS.n3392 VSS.n3397 4.5005
R12491 VSS.n3394 VSS.n3398 4.5005
R12492 VSS.n3395 VSS.n3399 4.5005
R12493 VSS.n3396 VSS.n3400 4.57324
R12494 VSS.n3392 VSS.n3390 0.147342
R12495 VSS.n3393 VSS.n3394 0.0732424
R12496 VSS.n3394 VSS.n3395 0.147342
R12497 VSS.n3397 VSS.n3401 0.0721009
R12498 VSS.n3402 VSS.n3398 4.5005
R12499 VSS.n3403 VSS.n3399 4.5005
R12500 VSS.n3404 VSS.n3400 4.5005
R12501 VSS.n3390 VSS.n3401 4.57442
R12502 VSS.n3397 VSS.n3398 0.147342
R12503 VSS.n3398 VSS.n3399 0.147342
R12504 VSS.n3399 VSS.n3400 0.147342
R12505 VSS.n3401 VSS.n3402 2.39784
R12506 VSS.n3402 VSS.n3403 0.147342
R12507 VSS.n3403 VSS.n3404 0.147342
R12508 VSS.n3404 VSS.t166 3.13212
R12509 VSS.n3382 VSS.n3377 4.5005
R12510 VSS.n3383 VSS.n3379 4.5005
R12511 VSS.n3384 VSS.n3380 4.5005
R12512 VSS.n3385 VSS.n3381 4.57324
R12513 VSS.n3375 VSS.n3377 0.147342
R12514 VSS.n3378 VSS.n3379 0.0732424
R12515 VSS.n3379 VSS.n3380 0.147342
R12516 VSS.n3386 VSS.n3382 0.0722544
R12517 VSS.n3387 VSS.n3383 4.5005
R12518 VSS.n3388 VSS.n3384 4.5005
R12519 VSS.n3389 VSS.n3385 4.5005
R12520 VSS.n3386 VSS.n3375 4.57426
R12521 VSS.n3382 VSS.n3383 0.147342
R12522 VSS.n3383 VSS.n3384 0.147342
R12523 VSS.n3384 VSS.n3385 0.147342
R12524 VSS.n3387 VSS.n3386 2.37296
R12525 VSS.n3388 VSS.n3387 0.127318
R12526 VSS.n3389 VSS.n3388 0.127318
R12527 VSS.t5 VSS.n3389 2.73618
R12528 VSS.n3362 VSS.n3367 4.5005
R12529 VSS.n3364 VSS.n3368 4.5005
R12530 VSS.n3365 VSS.n3369 4.5005
R12531 VSS.n3366 VSS.n3370 4.57324
R12532 VSS.n3362 VSS.n3360 0.147342
R12533 VSS.n3363 VSS.n3364 0.0732424
R12534 VSS.n3364 VSS.n3365 0.147342
R12535 VSS.n3367 VSS.n3371 0.0721009
R12536 VSS.n3372 VSS.n3368 4.5005
R12537 VSS.n3373 VSS.n3369 4.5005
R12538 VSS.n3374 VSS.n3370 4.5005
R12539 VSS.n3360 VSS.n3371 4.57442
R12540 VSS.n3367 VSS.n3368 0.147342
R12541 VSS.n3368 VSS.n3369 0.147342
R12542 VSS.n3369 VSS.n3370 0.147342
R12543 VSS.n3371 VSS.n3372 2.39784
R12544 VSS.n3372 VSS.n3373 0.147342
R12545 VSS.n3373 VSS.n3374 0.147342
R12546 VSS.n3374 VSS.t361 3.13212
R12547 VSS.n3347 VSS.n3352 4.5005
R12548 VSS.n3349 VSS.n3353 4.5005
R12549 VSS.n3350 VSS.n3354 4.5005
R12550 VSS.n3351 VSS.n3355 4.57324
R12551 VSS.n3347 VSS.n3345 0.147342
R12552 VSS.n3348 VSS.n3349 0.0732424
R12553 VSS.n3349 VSS.n3350 0.147342
R12554 VSS.n3352 VSS.n3356 0.0721009
R12555 VSS.n3357 VSS.n3353 4.5005
R12556 VSS.n3358 VSS.n3354 4.5005
R12557 VSS.n3359 VSS.n3355 4.5005
R12558 VSS.n3345 VSS.n3356 4.57442
R12559 VSS.n3352 VSS.n3353 0.147342
R12560 VSS.n3353 VSS.n3354 0.147342
R12561 VSS.n3354 VSS.n3355 0.147342
R12562 VSS.n3356 VSS.n3357 2.39784
R12563 VSS.n3357 VSS.n3358 0.147342
R12564 VSS.n3358 VSS.n3359 0.147342
R12565 VSS.n3359 VSS.t37 3.13212
R12566 VSS.n3332 VSS.n3337 4.5005
R12567 VSS.n3334 VSS.n3338 4.5005
R12568 VSS.n3335 VSS.n3339 4.5005
R12569 VSS.n3336 VSS.n3340 4.57324
R12570 VSS.n3332 VSS.n3330 0.147342
R12571 VSS.n3333 VSS.n3334 0.0732424
R12572 VSS.n3334 VSS.n3335 0.147342
R12573 VSS.n3337 VSS.n3341 0.0721009
R12574 VSS.n3342 VSS.n3338 4.5005
R12575 VSS.n3343 VSS.n3339 4.5005
R12576 VSS.n3344 VSS.n3340 4.5005
R12577 VSS.n3330 VSS.n3341 4.57442
R12578 VSS.n3337 VSS.n3338 0.147342
R12579 VSS.n3338 VSS.n3339 0.147342
R12580 VSS.n3339 VSS.n3340 0.147342
R12581 VSS.n3341 VSS.n3342 2.39784
R12582 VSS.n3342 VSS.n3343 0.147342
R12583 VSS.n3343 VSS.n3344 0.147342
R12584 VSS.n3344 VSS.t15 3.13212
R12585 VSS.n3322 VSS.n3317 4.5005
R12586 VSS.n3323 VSS.n3319 4.5005
R12587 VSS.n3324 VSS.n3320 4.5005
R12588 VSS.n3325 VSS.n3321 4.57324
R12589 VSS.n3315 VSS.n3317 0.147342
R12590 VSS.n3318 VSS.n3319 0.0732424
R12591 VSS.n3319 VSS.n3320 0.147342
R12592 VSS.n3326 VSS.n3322 0.0722544
R12593 VSS.n3327 VSS.n3323 4.5005
R12594 VSS.n3328 VSS.n3324 4.5005
R12595 VSS.n3329 VSS.n3325 4.5005
R12596 VSS.n3326 VSS.n3315 4.57426
R12597 VSS.n3322 VSS.n3323 0.147342
R12598 VSS.n3323 VSS.n3324 0.147342
R12599 VSS.n3324 VSS.n3325 0.147342
R12600 VSS.n3327 VSS.n3326 2.37296
R12601 VSS.n3328 VSS.n3327 0.127318
R12602 VSS.n3329 VSS.n3328 0.127318
R12603 VSS.t5 VSS.n3329 2.73618
R12604 VSS.n3302 VSS.n3307 4.5005
R12605 VSS.n3304 VSS.n3308 4.5005
R12606 VSS.n3305 VSS.n3309 4.5005
R12607 VSS.n3306 VSS.n3310 4.57324
R12608 VSS.n3302 VSS.n3300 0.147342
R12609 VSS.n3303 VSS.n3304 0.0732424
R12610 VSS.n3304 VSS.n3305 0.147342
R12611 VSS.n3307 VSS.n3311 0.0721009
R12612 VSS.n3312 VSS.n3308 4.5005
R12613 VSS.n3313 VSS.n3309 4.5005
R12614 VSS.n3314 VSS.n3310 4.5005
R12615 VSS.n3300 VSS.n3311 4.57442
R12616 VSS.n3307 VSS.n3308 0.147342
R12617 VSS.n3308 VSS.n3309 0.147342
R12618 VSS.n3309 VSS.n3310 0.147342
R12619 VSS.n3311 VSS.n3312 2.39784
R12620 VSS.n3312 VSS.n3313 0.147342
R12621 VSS.n3313 VSS.n3314 0.147342
R12622 VSS.n3314 VSS.t231 3.13212
R12623 VSS.n3287 VSS.n3292 4.5005
R12624 VSS.n3289 VSS.n3293 4.5005
R12625 VSS.n3290 VSS.n3294 4.5005
R12626 VSS.n3291 VSS.n3295 4.57324
R12627 VSS.n3287 VSS.n3285 0.147342
R12628 VSS.n3288 VSS.n3289 0.0732424
R12629 VSS.n3289 VSS.n3290 0.147342
R12630 VSS.n3292 VSS.n3296 0.0721009
R12631 VSS.n3297 VSS.n3293 4.5005
R12632 VSS.n3298 VSS.n3294 4.5005
R12633 VSS.n3299 VSS.n3295 4.5005
R12634 VSS.n3285 VSS.n3296 4.57442
R12635 VSS.n3292 VSS.n3293 0.147342
R12636 VSS.n3293 VSS.n3294 0.147342
R12637 VSS.n3294 VSS.n3295 0.147342
R12638 VSS.n3296 VSS.n3297 2.39784
R12639 VSS.n3297 VSS.n3298 0.147342
R12640 VSS.n3298 VSS.n3299 0.147342
R12641 VSS.n3299 VSS.t465 3.13212
R12642 VSS.n3272 VSS.n3277 4.5005
R12643 VSS.n3274 VSS.n3278 4.5005
R12644 VSS.n3275 VSS.n3279 4.5005
R12645 VSS.n3276 VSS.n3280 4.57324
R12646 VSS.n3272 VSS.n3270 0.147342
R12647 VSS.n3273 VSS.n3274 0.0732424
R12648 VSS.n3274 VSS.n3275 0.147342
R12649 VSS.n3277 VSS.n3281 0.0721009
R12650 VSS.n3282 VSS.n3278 4.5005
R12651 VSS.n3283 VSS.n3279 4.5005
R12652 VSS.n3284 VSS.n3280 4.5005
R12653 VSS.n3270 VSS.n3281 4.57442
R12654 VSS.n3277 VSS.n3278 0.147342
R12655 VSS.n3278 VSS.n3279 0.147342
R12656 VSS.n3279 VSS.n3280 0.147342
R12657 VSS.n3281 VSS.n3282 2.39784
R12658 VSS.n3282 VSS.n3283 0.147342
R12659 VSS.n3283 VSS.n3284 0.147342
R12660 VSS.n3284 VSS.t248 3.13212
R12661 VSS.n3257 VSS.n3262 4.5005
R12662 VSS.n3259 VSS.n3263 4.5005
R12663 VSS.n3260 VSS.n3264 4.5005
R12664 VSS.n3261 VSS.n3265 4.57324
R12665 VSS.n3257 VSS.n3255 0.147342
R12666 VSS.n3258 VSS.n3259 0.0732424
R12667 VSS.n3259 VSS.n3260 0.147342
R12668 VSS.n3262 VSS.n3266 0.0721009
R12669 VSS.n3267 VSS.n3263 4.5005
R12670 VSS.n3268 VSS.n3264 4.5005
R12671 VSS.n3269 VSS.n3265 4.5005
R12672 VSS.n3255 VSS.n3266 4.57442
R12673 VSS.n3262 VSS.n3263 0.147342
R12674 VSS.n3263 VSS.n3264 0.147342
R12675 VSS.n3264 VSS.n3265 0.147342
R12676 VSS.n3266 VSS.n3267 2.39784
R12677 VSS.n3267 VSS.n3268 0.147342
R12678 VSS.n3268 VSS.n3269 0.147342
R12679 VSS.n3269 VSS.t252 3.13212
R12680 VSS.n3247 VSS.n3242 4.5005
R12681 VSS.n3248 VSS.n3244 4.5005
R12682 VSS.n3249 VSS.n3245 4.5005
R12683 VSS.n3250 VSS.n3246 4.57324
R12684 VSS.n3240 VSS.n3242 0.147342
R12685 VSS.n3243 VSS.n3244 0.0732424
R12686 VSS.n3244 VSS.n3245 0.147342
R12687 VSS.n3251 VSS.n3247 0.0722544
R12688 VSS.n3252 VSS.n3248 4.5005
R12689 VSS.n3253 VSS.n3249 4.5005
R12690 VSS.n3254 VSS.n3250 4.5005
R12691 VSS.n3251 VSS.n3240 4.57426
R12692 VSS.n3247 VSS.n3248 0.147342
R12693 VSS.n3248 VSS.n3249 0.147342
R12694 VSS.n3249 VSS.n3250 0.147342
R12695 VSS.n3252 VSS.n3251 2.37296
R12696 VSS.n3253 VSS.n3252 0.127318
R12697 VSS.n3254 VSS.n3253 0.127318
R12698 VSS.t5 VSS.n3254 2.73618
R12699 VSS.n3227 VSS.n3232 4.5005
R12700 VSS.n3229 VSS.n3233 4.5005
R12701 VSS.n3230 VSS.n3234 4.5005
R12702 VSS.n3231 VSS.n3235 4.57324
R12703 VSS.n3227 VSS.n3225 0.147342
R12704 VSS.n3228 VSS.n3229 0.0732424
R12705 VSS.n3229 VSS.n3230 0.147342
R12706 VSS.n3232 VSS.n3236 0.0721009
R12707 VSS.n3237 VSS.n3233 4.5005
R12708 VSS.n3238 VSS.n3234 4.5005
R12709 VSS.n3239 VSS.n3235 4.5005
R12710 VSS.n3225 VSS.n3236 4.57442
R12711 VSS.n3232 VSS.n3233 0.147342
R12712 VSS.n3233 VSS.n3234 0.147342
R12713 VSS.n3234 VSS.n3235 0.147342
R12714 VSS.n3236 VSS.n3237 2.39784
R12715 VSS.n3237 VSS.n3238 0.147342
R12716 VSS.n3238 VSS.n3239 0.147342
R12717 VSS.n3239 VSS.t276 3.13212
R12718 VSS.n3212 VSS.n3217 4.5005
R12719 VSS.n3214 VSS.n3218 4.5005
R12720 VSS.n3215 VSS.n3219 4.5005
R12721 VSS.n3216 VSS.n3220 4.57324
R12722 VSS.n3212 VSS.n3210 0.147342
R12723 VSS.n3213 VSS.n3214 0.0732424
R12724 VSS.n3214 VSS.n3215 0.147342
R12725 VSS.n3217 VSS.n3221 0.0721009
R12726 VSS.n3222 VSS.n3218 4.5005
R12727 VSS.n3223 VSS.n3219 4.5005
R12728 VSS.n3224 VSS.n3220 4.5005
R12729 VSS.n3210 VSS.n3221 4.57442
R12730 VSS.n3217 VSS.n3218 0.147342
R12731 VSS.n3218 VSS.n3219 0.147342
R12732 VSS.n3219 VSS.n3220 0.147342
R12733 VSS.n3221 VSS.n3222 2.39784
R12734 VSS.n3222 VSS.n3223 0.147342
R12735 VSS.n3223 VSS.n3224 0.147342
R12736 VSS.n3224 VSS.t91 3.13212
R12737 VSS.n3197 VSS.n3202 4.5005
R12738 VSS.n3199 VSS.n3203 4.5005
R12739 VSS.n3200 VSS.n3204 4.5005
R12740 VSS.n3201 VSS.n3205 4.57324
R12741 VSS.n3197 VSS.n3195 0.147342
R12742 VSS.n3198 VSS.n3199 0.0732424
R12743 VSS.n3199 VSS.n3200 0.147342
R12744 VSS.n3202 VSS.n3206 0.0721009
R12745 VSS.n3207 VSS.n3203 4.5005
R12746 VSS.n3208 VSS.n3204 4.5005
R12747 VSS.n3209 VSS.n3205 4.5005
R12748 VSS.n3195 VSS.n3206 4.57442
R12749 VSS.n3202 VSS.n3203 0.147342
R12750 VSS.n3203 VSS.n3204 0.147342
R12751 VSS.n3204 VSS.n3205 0.147342
R12752 VSS.n3206 VSS.n3207 2.39784
R12753 VSS.n3207 VSS.n3208 0.147342
R12754 VSS.n3208 VSS.n3209 0.147342
R12755 VSS.n3209 VSS.t121 3.13212
R12756 VSS.n3187 VSS.n3182 4.5005
R12757 VSS.n3188 VSS.n3184 4.5005
R12758 VSS.n3189 VSS.n3185 4.5005
R12759 VSS.n3190 VSS.n3186 4.57324
R12760 VSS.n3180 VSS.n3182 0.147342
R12761 VSS.n3183 VSS.n3184 0.0732424
R12762 VSS.n3184 VSS.n3185 0.147342
R12763 VSS.n3191 VSS.n3187 0.0722544
R12764 VSS.n3192 VSS.n3188 4.5005
R12765 VSS.n3193 VSS.n3189 4.5005
R12766 VSS.n3194 VSS.n3190 4.5005
R12767 VSS.n3191 VSS.n3180 4.57426
R12768 VSS.n3187 VSS.n3188 0.147342
R12769 VSS.n3188 VSS.n3189 0.147342
R12770 VSS.n3189 VSS.n3190 0.147342
R12771 VSS.n3192 VSS.n3191 2.37296
R12772 VSS.n3193 VSS.n3192 0.127318
R12773 VSS.n3194 VSS.n3193 0.127318
R12774 VSS.t5 VSS.n3194 2.73618
R12775 VSS.n3167 VSS.n3172 4.5005
R12776 VSS.n3169 VSS.n3173 4.5005
R12777 VSS.n3170 VSS.n3174 4.5005
R12778 VSS.n3171 VSS.n3175 4.57324
R12779 VSS.n3167 VSS.n3165 0.147342
R12780 VSS.n3168 VSS.n3169 0.0732424
R12781 VSS.n3169 VSS.n3170 0.147342
R12782 VSS.n3172 VSS.n3176 0.0721009
R12783 VSS.n3177 VSS.n3173 4.5005
R12784 VSS.n3178 VSS.n3174 4.5005
R12785 VSS.n3179 VSS.n3175 4.5005
R12786 VSS.n3165 VSS.n3176 4.57442
R12787 VSS.n3172 VSS.n3173 0.147342
R12788 VSS.n3173 VSS.n3174 0.147342
R12789 VSS.n3174 VSS.n3175 0.147342
R12790 VSS.n3176 VSS.n3177 2.39784
R12791 VSS.n3177 VSS.n3178 0.147342
R12792 VSS.n3178 VSS.n3179 0.147342
R12793 VSS.n3179 VSS.t72 3.13212
R12794 VSS.n3152 VSS.n3157 4.5005
R12795 VSS.n3154 VSS.n3158 4.5005
R12796 VSS.n3155 VSS.n3159 4.5005
R12797 VSS.n3156 VSS.n3160 4.57324
R12798 VSS.n3152 VSS.n3150 0.147342
R12799 VSS.n3153 VSS.n3154 0.0732424
R12800 VSS.n3154 VSS.n3155 0.147342
R12801 VSS.n3157 VSS.n3161 0.0721009
R12802 VSS.n3162 VSS.n3158 4.5005
R12803 VSS.n3163 VSS.n3159 4.5005
R12804 VSS.n3164 VSS.n3160 4.5005
R12805 VSS.n3150 VSS.n3161 4.57442
R12806 VSS.n3157 VSS.n3158 0.147342
R12807 VSS.n3158 VSS.n3159 0.147342
R12808 VSS.n3159 VSS.n3160 0.147342
R12809 VSS.n3161 VSS.n3162 2.39784
R12810 VSS.n3162 VSS.n3163 0.147342
R12811 VSS.n3163 VSS.n3164 0.147342
R12812 VSS.n3164 VSS.t478 3.13212
R12813 VSS.n3137 VSS.n3142 4.5005
R12814 VSS.n3139 VSS.n3143 4.5005
R12815 VSS.n3140 VSS.n3144 4.5005
R12816 VSS.n3141 VSS.n3145 4.57324
R12817 VSS.n3137 VSS.n3135 0.147342
R12818 VSS.n3138 VSS.n3139 0.0732424
R12819 VSS.n3139 VSS.n3140 0.147342
R12820 VSS.n3142 VSS.n3146 0.0721009
R12821 VSS.n3147 VSS.n3143 4.5005
R12822 VSS.n3148 VSS.n3144 4.5005
R12823 VSS.n3149 VSS.n3145 4.5005
R12824 VSS.n3135 VSS.n3146 4.57442
R12825 VSS.n3142 VSS.n3143 0.147342
R12826 VSS.n3143 VSS.n3144 0.147342
R12827 VSS.n3144 VSS.n3145 0.147342
R12828 VSS.n3146 VSS.n3147 2.39784
R12829 VSS.n3147 VSS.n3148 0.147342
R12830 VSS.n3148 VSS.n3149 0.147342
R12831 VSS.n3149 VSS.t144 3.13212
R12832 VSS.n3122 VSS.n3127 4.5005
R12833 VSS.n3124 VSS.n3128 4.5005
R12834 VSS.n3125 VSS.n3129 4.5005
R12835 VSS.n3126 VSS.n3130 4.57324
R12836 VSS.n3122 VSS.n3120 0.147342
R12837 VSS.n3123 VSS.n3124 0.0732424
R12838 VSS.n3124 VSS.n3125 0.147342
R12839 VSS.n3127 VSS.n3131 0.0721009
R12840 VSS.n3132 VSS.n3128 4.5005
R12841 VSS.n3133 VSS.n3129 4.5005
R12842 VSS.n3134 VSS.n3130 4.5005
R12843 VSS.n3120 VSS.n3131 4.57442
R12844 VSS.n3127 VSS.n3128 0.147342
R12845 VSS.n3128 VSS.n3129 0.147342
R12846 VSS.n3129 VSS.n3130 0.147342
R12847 VSS.n3131 VSS.n3132 2.39784
R12848 VSS.n3132 VSS.n3133 0.147342
R12849 VSS.n3133 VSS.n3134 0.147342
R12850 VSS.n3134 VSS.t11 3.13212
R12851 VSS.n3107 VSS.n3112 4.5005
R12852 VSS.n3109 VSS.n3113 4.5005
R12853 VSS.n3110 VSS.n3114 4.5005
R12854 VSS.n3111 VSS.n3115 4.57324
R12855 VSS.n3107 VSS.n3105 0.147342
R12856 VSS.n3108 VSS.n3109 0.0732424
R12857 VSS.n3109 VSS.n3110 0.147342
R12858 VSS.n3112 VSS.n3116 0.0721009
R12859 VSS.n3117 VSS.n3113 4.5005
R12860 VSS.n3118 VSS.n3114 4.5005
R12861 VSS.n3119 VSS.n3115 4.5005
R12862 VSS.n3105 VSS.n3116 4.57442
R12863 VSS.n3112 VSS.n3113 0.147342
R12864 VSS.n3113 VSS.n3114 0.147342
R12865 VSS.n3114 VSS.n3115 0.147342
R12866 VSS.n3116 VSS.n3117 2.39784
R12867 VSS.n3117 VSS.n3118 0.147342
R12868 VSS.n3118 VSS.n3119 0.147342
R12869 VSS.n3119 VSS.t193 3.13212
R12870 VSS.n3092 VSS.n3097 4.5005
R12871 VSS.n3094 VSS.n3098 4.5005
R12872 VSS.n3095 VSS.n3099 4.5005
R12873 VSS.n3096 VSS.n3100 4.57324
R12874 VSS.n3092 VSS.n3090 0.147342
R12875 VSS.n3093 VSS.n3094 0.0732424
R12876 VSS.n3094 VSS.n3095 0.147342
R12877 VSS.n3097 VSS.n3101 0.0721009
R12878 VSS.n3102 VSS.n3098 4.5005
R12879 VSS.n3103 VSS.n3099 4.5005
R12880 VSS.n3104 VSS.n3100 4.5005
R12881 VSS.n3090 VSS.n3101 4.57442
R12882 VSS.n3097 VSS.n3098 0.147342
R12883 VSS.n3098 VSS.n3099 0.147342
R12884 VSS.n3099 VSS.n3100 0.147342
R12885 VSS.n3101 VSS.n3102 2.39784
R12886 VSS.n3102 VSS.n3103 0.147342
R12887 VSS.n3103 VSS.n3104 0.147342
R12888 VSS.n3104 VSS.t497 3.13212
R12889 VSS.n3082 VSS.n3077 4.5005
R12890 VSS.n3083 VSS.n3079 4.5005
R12891 VSS.n3084 VSS.n3080 4.5005
R12892 VSS.n3085 VSS.n3081 4.57324
R12893 VSS.n3075 VSS.n3077 0.147342
R12894 VSS.n3078 VSS.n3079 0.0732424
R12895 VSS.n3079 VSS.n3080 0.147342
R12896 VSS.n3086 VSS.n3082 0.0722544
R12897 VSS.n3087 VSS.n3083 4.5005
R12898 VSS.n3088 VSS.n3084 4.5005
R12899 VSS.n3089 VSS.n3085 4.5005
R12900 VSS.n3086 VSS.n3075 4.57426
R12901 VSS.n3082 VSS.n3083 0.147342
R12902 VSS.n3083 VSS.n3084 0.147342
R12903 VSS.n3084 VSS.n3085 0.147342
R12904 VSS.n3087 VSS.n3086 2.37296
R12905 VSS.n3088 VSS.n3087 0.127318
R12906 VSS.n3089 VSS.n3088 0.127318
R12907 VSS.t5 VSS.n3089 2.73618
R12908 VSS.n3062 VSS.n3067 4.5005
R12909 VSS.n3064 VSS.n3068 4.5005
R12910 VSS.n3065 VSS.n3069 4.5005
R12911 VSS.n3066 VSS.n3070 4.57324
R12912 VSS.n3062 VSS.n3060 0.147342
R12913 VSS.n3063 VSS.n3064 0.0732424
R12914 VSS.n3064 VSS.n3065 0.147342
R12915 VSS.n3067 VSS.n3071 0.0721009
R12916 VSS.n3072 VSS.n3068 4.5005
R12917 VSS.n3073 VSS.n3069 4.5005
R12918 VSS.n3074 VSS.n3070 4.5005
R12919 VSS.n3060 VSS.n3071 4.57442
R12920 VSS.n3067 VSS.n3068 0.147342
R12921 VSS.n3068 VSS.n3069 0.147342
R12922 VSS.n3069 VSS.n3070 0.147342
R12923 VSS.n3071 VSS.n3072 2.39784
R12924 VSS.n3072 VSS.n3073 0.147342
R12925 VSS.n3073 VSS.n3074 0.147342
R12926 VSS.n3074 VSS.t363 3.13212
R12927 VSS.n3047 VSS.n3052 4.5005
R12928 VSS.n3049 VSS.n3053 4.5005
R12929 VSS.n3050 VSS.n3054 4.5005
R12930 VSS.n3051 VSS.n3055 4.57324
R12931 VSS.n3047 VSS.n3045 0.147342
R12932 VSS.n3048 VSS.n3049 0.0732424
R12933 VSS.n3049 VSS.n3050 0.147342
R12934 VSS.n3052 VSS.n3056 0.0721009
R12935 VSS.n3057 VSS.n3053 4.5005
R12936 VSS.n3058 VSS.n3054 4.5005
R12937 VSS.n3059 VSS.n3055 4.5005
R12938 VSS.n3045 VSS.n3056 4.57442
R12939 VSS.n3052 VSS.n3053 0.147342
R12940 VSS.n3053 VSS.n3054 0.147342
R12941 VSS.n3054 VSS.n3055 0.147342
R12942 VSS.n3056 VSS.n3057 2.39784
R12943 VSS.n3057 VSS.n3058 0.147342
R12944 VSS.n3058 VSS.n3059 0.147342
R12945 VSS.n3059 VSS.t125 3.13212
R12946 VSS.n3032 VSS.n3037 4.5005
R12947 VSS.n3034 VSS.n3038 4.5005
R12948 VSS.n3035 VSS.n3039 4.5005
R12949 VSS.n3036 VSS.n3040 4.57324
R12950 VSS.n3032 VSS.n3030 0.147342
R12951 VSS.n3033 VSS.n3034 0.0732424
R12952 VSS.n3034 VSS.n3035 0.147342
R12953 VSS.n3037 VSS.n3041 0.0721009
R12954 VSS.n3042 VSS.n3038 4.5005
R12955 VSS.n3043 VSS.n3039 4.5005
R12956 VSS.n3044 VSS.n3040 4.5005
R12957 VSS.n3030 VSS.n3041 4.57442
R12958 VSS.n3037 VSS.n3038 0.147342
R12959 VSS.n3038 VSS.n3039 0.147342
R12960 VSS.n3039 VSS.n3040 0.147342
R12961 VSS.n3041 VSS.n3042 2.39784
R12962 VSS.n3042 VSS.n3043 0.147342
R12963 VSS.n3043 VSS.n3044 0.147342
R12964 VSS.n3044 VSS.t17 3.13212
R12965 VSS.n3022 VSS.n3017 4.5005
R12966 VSS.n3023 VSS.n3019 4.5005
R12967 VSS.n3024 VSS.n3020 4.5005
R12968 VSS.n3025 VSS.n3021 4.57324
R12969 VSS.n3015 VSS.n3017 0.147342
R12970 VSS.n3018 VSS.n3019 0.0732424
R12971 VSS.n3019 VSS.n3020 0.147342
R12972 VSS.n3026 VSS.n3022 0.0722544
R12973 VSS.n3027 VSS.n3023 4.5005
R12974 VSS.n3028 VSS.n3024 4.5005
R12975 VSS.n3029 VSS.n3025 4.5005
R12976 VSS.n3026 VSS.n3015 4.57426
R12977 VSS.n3022 VSS.n3023 0.147342
R12978 VSS.n3023 VSS.n3024 0.147342
R12979 VSS.n3024 VSS.n3025 0.147342
R12980 VSS.n3027 VSS.n3026 2.37296
R12981 VSS.n3028 VSS.n3027 0.127318
R12982 VSS.n3029 VSS.n3028 0.127318
R12983 VSS.t5 VSS.n3029 2.73618
R12984 VSS.n3002 VSS.n3007 4.5005
R12985 VSS.n3004 VSS.n3008 4.5005
R12986 VSS.n3005 VSS.n3009 4.5005
R12987 VSS.n3006 VSS.n3010 4.57324
R12988 VSS.n3002 VSS.n3000 0.147342
R12989 VSS.n3003 VSS.n3004 0.0732424
R12990 VSS.n3004 VSS.n3005 0.147342
R12991 VSS.n3007 VSS.n3011 0.0721009
R12992 VSS.n3012 VSS.n3008 4.5005
R12993 VSS.n3013 VSS.n3009 4.5005
R12994 VSS.n3014 VSS.n3010 4.5005
R12995 VSS.n3000 VSS.n3011 4.57442
R12996 VSS.n3007 VSS.n3008 0.147342
R12997 VSS.n3008 VSS.n3009 0.147342
R12998 VSS.n3009 VSS.n3010 0.147342
R12999 VSS.n3011 VSS.n3012 2.39784
R13000 VSS.n3012 VSS.n3013 0.147342
R13001 VSS.n3013 VSS.n3014 0.147342
R13002 VSS.n3014 VSS.t234 3.13212
R13003 VSS.n2987 VSS.n2992 4.5005
R13004 VSS.n2989 VSS.n2993 4.5005
R13005 VSS.n2990 VSS.n2994 4.5005
R13006 VSS.n2991 VSS.n2995 4.57324
R13007 VSS.n2987 VSS.n2985 0.147342
R13008 VSS.n2988 VSS.n2989 0.0732424
R13009 VSS.n2989 VSS.n2990 0.147342
R13010 VSS.n2992 VSS.n2996 0.0721009
R13011 VSS.n2997 VSS.n2993 4.5005
R13012 VSS.n2998 VSS.n2994 4.5005
R13013 VSS.n2999 VSS.n2995 4.5005
R13014 VSS.n2985 VSS.n2996 4.57442
R13015 VSS.n2992 VSS.n2993 0.147342
R13016 VSS.n2993 VSS.n2994 0.147342
R13017 VSS.n2994 VSS.n2995 0.147342
R13018 VSS.n2996 VSS.n2997 2.39784
R13019 VSS.n2997 VSS.n2998 0.147342
R13020 VSS.n2998 VSS.n2999 0.147342
R13021 VSS.n2999 VSS.t258 3.13212
R13022 VSS.n2972 VSS.n2977 4.5005
R13023 VSS.n2974 VSS.n2978 4.5005
R13024 VSS.n2975 VSS.n2979 4.5005
R13025 VSS.n2976 VSS.n2980 4.57324
R13026 VSS.n2972 VSS.n2970 0.147342
R13027 VSS.n2973 VSS.n2974 0.0732424
R13028 VSS.n2974 VSS.n2975 0.147342
R13029 VSS.n2977 VSS.n2981 0.0721009
R13030 VSS.n2982 VSS.n2978 4.5005
R13031 VSS.n2983 VSS.n2979 4.5005
R13032 VSS.n2984 VSS.n2980 4.5005
R13033 VSS.n2970 VSS.n2981 4.57442
R13034 VSS.n2977 VSS.n2978 0.147342
R13035 VSS.n2978 VSS.n2979 0.147342
R13036 VSS.n2979 VSS.n2980 0.147342
R13037 VSS.n2981 VSS.n2982 2.39784
R13038 VSS.n2982 VSS.n2983 0.147342
R13039 VSS.n2983 VSS.n2984 0.147342
R13040 VSS.n2984 VSS.t77 3.13212
R13041 VSS.n2957 VSS.n2962 4.5005
R13042 VSS.n2959 VSS.n2963 4.5005
R13043 VSS.n2960 VSS.n2964 4.5005
R13044 VSS.n2961 VSS.n2965 4.57324
R13045 VSS.n2957 VSS.n2955 0.147342
R13046 VSS.n2958 VSS.n2959 0.0732424
R13047 VSS.n2959 VSS.n2960 0.147342
R13048 VSS.n2962 VSS.n2966 0.0721009
R13049 VSS.n2967 VSS.n2963 4.5005
R13050 VSS.n2968 VSS.n2964 4.5005
R13051 VSS.n2969 VSS.n2965 4.5005
R13052 VSS.n2955 VSS.n2966 4.57442
R13053 VSS.n2962 VSS.n2963 0.147342
R13054 VSS.n2963 VSS.n2964 0.147342
R13055 VSS.n2964 VSS.n2965 0.147342
R13056 VSS.n2966 VSS.n2967 2.39784
R13057 VSS.n2967 VSS.n2968 0.147342
R13058 VSS.n2968 VSS.n2969 0.147342
R13059 VSS.n2969 VSS.t253 3.13212
R13060 VSS.n2947 VSS.n2942 4.5005
R13061 VSS.n2948 VSS.n2944 4.5005
R13062 VSS.n2949 VSS.n2945 4.5005
R13063 VSS.n2950 VSS.n2946 4.57324
R13064 VSS.n2940 VSS.n2942 0.147342
R13065 VSS.n2943 VSS.n2944 0.0732424
R13066 VSS.n2944 VSS.n2945 0.147342
R13067 VSS.n2951 VSS.n2947 0.0722544
R13068 VSS.n2952 VSS.n2948 4.5005
R13069 VSS.n2953 VSS.n2949 4.5005
R13070 VSS.n2954 VSS.n2950 4.5005
R13071 VSS.n2951 VSS.n2940 4.57426
R13072 VSS.n2947 VSS.n2948 0.147342
R13073 VSS.n2948 VSS.n2949 0.147342
R13074 VSS.n2949 VSS.n2950 0.147342
R13075 VSS.n2952 VSS.n2951 2.37296
R13076 VSS.n2953 VSS.n2952 0.127318
R13077 VSS.n2954 VSS.n2953 0.127318
R13078 VSS.t5 VSS.n2954 2.73618
R13079 VSS.n2927 VSS.n2932 4.5005
R13080 VSS.n2929 VSS.n2933 4.5005
R13081 VSS.n2930 VSS.n2934 4.5005
R13082 VSS.n2931 VSS.n2935 4.57324
R13083 VSS.n2927 VSS.n2925 0.147342
R13084 VSS.n2928 VSS.n2929 0.0732424
R13085 VSS.n2929 VSS.n2930 0.147342
R13086 VSS.n2932 VSS.n2936 0.0721009
R13087 VSS.n2937 VSS.n2933 4.5005
R13088 VSS.n2938 VSS.n2934 4.5005
R13089 VSS.n2939 VSS.n2935 4.5005
R13090 VSS.n2925 VSS.n2936 4.57442
R13091 VSS.n2932 VSS.n2933 0.147342
R13092 VSS.n2933 VSS.n2934 0.147342
R13093 VSS.n2934 VSS.n2935 0.147342
R13094 VSS.n2936 VSS.n2937 2.39784
R13095 VSS.n2937 VSS.n2938 0.147342
R13096 VSS.n2938 VSS.n2939 0.147342
R13097 VSS.n2939 VSS.t419 3.13212
R13098 VSS.n2912 VSS.n2917 4.5005
R13099 VSS.n2914 VSS.n2918 4.5005
R13100 VSS.n2915 VSS.n2919 4.5005
R13101 VSS.n2916 VSS.n2920 4.57324
R13102 VSS.n2912 VSS.n2910 0.147342
R13103 VSS.n2913 VSS.n2914 0.0732424
R13104 VSS.n2914 VSS.n2915 0.147342
R13105 VSS.n2917 VSS.n2921 0.0721009
R13106 VSS.n2922 VSS.n2918 4.5005
R13107 VSS.n2923 VSS.n2919 4.5005
R13108 VSS.n2924 VSS.n2920 4.5005
R13109 VSS.n2910 VSS.n2921 4.57442
R13110 VSS.n2917 VSS.n2918 0.147342
R13111 VSS.n2918 VSS.n2919 0.147342
R13112 VSS.n2919 VSS.n2920 0.147342
R13113 VSS.n2921 VSS.n2922 2.39784
R13114 VSS.n2922 VSS.n2923 0.147342
R13115 VSS.n2923 VSS.n2924 0.147342
R13116 VSS.n2924 VSS.t87 3.13212
R13117 VSS.n2897 VSS.n2902 4.5005
R13118 VSS.n2899 VSS.n2903 4.5005
R13119 VSS.n2900 VSS.n2904 4.5005
R13120 VSS.n2901 VSS.n2905 4.57324
R13121 VSS.n2897 VSS.n2895 0.147342
R13122 VSS.n2898 VSS.n2899 0.0732424
R13123 VSS.n2899 VSS.n2900 0.147342
R13124 VSS.n2902 VSS.n2906 0.0721009
R13125 VSS.n2907 VSS.n2903 4.5005
R13126 VSS.n2908 VSS.n2904 4.5005
R13127 VSS.n2909 VSS.n2905 4.5005
R13128 VSS.n2895 VSS.n2906 4.57442
R13129 VSS.n2902 VSS.n2903 0.147342
R13130 VSS.n2903 VSS.n2904 0.147342
R13131 VSS.n2904 VSS.n2905 0.147342
R13132 VSS.n2906 VSS.n2907 2.39784
R13133 VSS.n2907 VSS.n2908 0.147342
R13134 VSS.n2908 VSS.n2909 0.147342
R13135 VSS.n2909 VSS.t118 3.13212
R13136 VSS.n2887 VSS.n2882 4.5005
R13137 VSS.n2888 VSS.n2884 4.5005
R13138 VSS.n2889 VSS.n2885 4.5005
R13139 VSS.n2890 VSS.n2886 4.57324
R13140 VSS.n2880 VSS.n2882 0.147342
R13141 VSS.n2883 VSS.n2884 0.0732424
R13142 VSS.n2884 VSS.n2885 0.147342
R13143 VSS.n2891 VSS.n2887 0.0722544
R13144 VSS.n2892 VSS.n2888 4.5005
R13145 VSS.n2893 VSS.n2889 4.5005
R13146 VSS.n2894 VSS.n2890 4.5005
R13147 VSS.n2891 VSS.n2880 4.57426
R13148 VSS.n2887 VSS.n2888 0.147342
R13149 VSS.n2888 VSS.n2889 0.147342
R13150 VSS.n2889 VSS.n2890 0.147342
R13151 VSS.n2892 VSS.n2891 2.37296
R13152 VSS.n2893 VSS.n2892 0.127318
R13153 VSS.n2894 VSS.n2893 0.127318
R13154 VSS.t5 VSS.n2894 2.73618
R13155 VSS.n2867 VSS.n2872 4.5005
R13156 VSS.n2869 VSS.n2873 4.5005
R13157 VSS.n2870 VSS.n2874 4.5005
R13158 VSS.n2871 VSS.n2875 4.57324
R13159 VSS.n2867 VSS.n2865 0.147342
R13160 VSS.n2868 VSS.n2869 0.0732424
R13161 VSS.n2869 VSS.n2870 0.147342
R13162 VSS.n2872 VSS.n2876 0.0721009
R13163 VSS.n2877 VSS.n2873 4.5005
R13164 VSS.n2878 VSS.n2874 4.5005
R13165 VSS.n2879 VSS.n2875 4.5005
R13166 VSS.n2865 VSS.n2876 4.57442
R13167 VSS.n2872 VSS.n2873 0.147342
R13168 VSS.n2873 VSS.n2874 0.147342
R13169 VSS.n2874 VSS.n2875 0.147342
R13170 VSS.n2876 VSS.n2877 2.39784
R13171 VSS.n2877 VSS.n2878 0.147342
R13172 VSS.n2878 VSS.n2879 0.147342
R13173 VSS.n2879 VSS.t74 3.13212
R13174 VSS.n2852 VSS.n2857 4.5005
R13175 VSS.n2854 VSS.n2858 4.5005
R13176 VSS.n2855 VSS.n2859 4.5005
R13177 VSS.n2856 VSS.n2860 4.57324
R13178 VSS.n2852 VSS.n2850 0.147342
R13179 VSS.n2853 VSS.n2854 0.0732424
R13180 VSS.n2854 VSS.n2855 0.147342
R13181 VSS.n2857 VSS.n2861 0.0721009
R13182 VSS.n2862 VSS.n2858 4.5005
R13183 VSS.n2863 VSS.n2859 4.5005
R13184 VSS.n2864 VSS.n2860 4.5005
R13185 VSS.n2850 VSS.n2861 4.57442
R13186 VSS.n2857 VSS.n2858 0.147342
R13187 VSS.n2858 VSS.n2859 0.147342
R13188 VSS.n2859 VSS.n2860 0.147342
R13189 VSS.n2861 VSS.n2862 2.39784
R13190 VSS.n2862 VSS.n2863 0.147342
R13191 VSS.n2863 VSS.n2864 0.147342
R13192 VSS.n2864 VSS.t183 3.13212
R13193 VSS.n2837 VSS.n2842 4.5005
R13194 VSS.n2839 VSS.n2843 4.5005
R13195 VSS.n2840 VSS.n2844 4.5005
R13196 VSS.n2841 VSS.n2845 4.57324
R13197 VSS.n2837 VSS.n2835 0.147342
R13198 VSS.n2838 VSS.n2839 0.0732424
R13199 VSS.n2839 VSS.n2840 0.147342
R13200 VSS.n2842 VSS.n2846 0.0721009
R13201 VSS.n2847 VSS.n2843 4.5005
R13202 VSS.n2848 VSS.n2844 4.5005
R13203 VSS.n2849 VSS.n2845 4.5005
R13204 VSS.n2835 VSS.n2846 4.57442
R13205 VSS.n2842 VSS.n2843 0.147342
R13206 VSS.n2843 VSS.n2844 0.147342
R13207 VSS.n2844 VSS.n2845 0.147342
R13208 VSS.n2846 VSS.n2847 2.39784
R13209 VSS.n2847 VSS.n2848 0.147342
R13210 VSS.n2848 VSS.n2849 0.147342
R13211 VSS.n2849 VSS.t327 3.13212
R13212 VSS.n2822 VSS.n2827 4.5005
R13213 VSS.n2824 VSS.n2828 4.5005
R13214 VSS.n2825 VSS.n2829 4.5005
R13215 VSS.n2826 VSS.n2830 4.57324
R13216 VSS.n2822 VSS.n2820 0.147342
R13217 VSS.n2823 VSS.n2824 0.0732424
R13218 VSS.n2824 VSS.n2825 0.147342
R13219 VSS.n2827 VSS.n2831 0.0721009
R13220 VSS.n2832 VSS.n2828 4.5005
R13221 VSS.n2833 VSS.n2829 4.5005
R13222 VSS.n2834 VSS.n2830 4.5005
R13223 VSS.n2820 VSS.n2831 4.57442
R13224 VSS.n2827 VSS.n2828 0.147342
R13225 VSS.n2828 VSS.n2829 0.147342
R13226 VSS.n2829 VSS.n2830 0.147342
R13227 VSS.n2831 VSS.n2832 2.39784
R13228 VSS.n2832 VSS.n2833 0.147342
R13229 VSS.n2833 VSS.n2834 0.147342
R13230 VSS.n2834 VSS.t9 3.13212
R13231 VSS.n2807 VSS.n2812 4.5005
R13232 VSS.n2809 VSS.n2813 4.5005
R13233 VSS.n2810 VSS.n2814 4.5005
R13234 VSS.n2811 VSS.n2815 4.57324
R13235 VSS.n2807 VSS.n2805 0.147342
R13236 VSS.n2808 VSS.n2809 0.0732424
R13237 VSS.n2809 VSS.n2810 0.147342
R13238 VSS.n2812 VSS.n2816 0.0721009
R13239 VSS.n2817 VSS.n2813 4.5005
R13240 VSS.n2818 VSS.n2814 4.5005
R13241 VSS.n2819 VSS.n2815 4.5005
R13242 VSS.n2805 VSS.n2816 4.57442
R13243 VSS.n2812 VSS.n2813 0.147342
R13244 VSS.n2813 VSS.n2814 0.147342
R13245 VSS.n2814 VSS.n2815 0.147342
R13246 VSS.n2816 VSS.n2817 2.39784
R13247 VSS.n2817 VSS.n2818 0.147342
R13248 VSS.n2818 VSS.n2819 0.147342
R13249 VSS.n2819 VSS.t195 3.13212
R13250 VSS.n2792 VSS.n2797 4.5005
R13251 VSS.n2794 VSS.n2798 4.5005
R13252 VSS.n2795 VSS.n2799 4.5005
R13253 VSS.n2796 VSS.n2800 4.57324
R13254 VSS.n2792 VSS.n2790 0.147342
R13255 VSS.n2793 VSS.n2794 0.0732424
R13256 VSS.n2794 VSS.n2795 0.147342
R13257 VSS.n2797 VSS.n2801 0.0721009
R13258 VSS.n2802 VSS.n2798 4.5005
R13259 VSS.n2803 VSS.n2799 4.5005
R13260 VSS.n2804 VSS.n2800 4.5005
R13261 VSS.n2790 VSS.n2801 4.57442
R13262 VSS.n2797 VSS.n2798 0.147342
R13263 VSS.n2798 VSS.n2799 0.147342
R13264 VSS.n2799 VSS.n2800 0.147342
R13265 VSS.n2801 VSS.n2802 2.39784
R13266 VSS.n2802 VSS.n2803 0.147342
R13267 VSS.n2803 VSS.n2804 0.147342
R13268 VSS.n2804 VSS.t167 3.13212
R13269 VSS.n2782 VSS.n2777 4.5005
R13270 VSS.n2783 VSS.n2779 4.5005
R13271 VSS.n2784 VSS.n2780 4.5005
R13272 VSS.n2785 VSS.n2781 4.57324
R13273 VSS.n2775 VSS.n2777 0.147342
R13274 VSS.n2778 VSS.n2779 0.0732424
R13275 VSS.n2779 VSS.n2780 0.147342
R13276 VSS.n2786 VSS.n2782 0.0722544
R13277 VSS.n2787 VSS.n2783 4.5005
R13278 VSS.n2788 VSS.n2784 4.5005
R13279 VSS.n2789 VSS.n2785 4.5005
R13280 VSS.n2786 VSS.n2775 4.57426
R13281 VSS.n2782 VSS.n2783 0.147342
R13282 VSS.n2783 VSS.n2784 0.147342
R13283 VSS.n2784 VSS.n2785 0.147342
R13284 VSS.n2787 VSS.n2786 2.37296
R13285 VSS.n2788 VSS.n2787 0.127318
R13286 VSS.n2789 VSS.n2788 0.127318
R13287 VSS.t5 VSS.n2789 2.73618
R13288 VSS.n2762 VSS.n2767 4.5005
R13289 VSS.n2764 VSS.n2768 4.5005
R13290 VSS.n2765 VSS.n2769 4.5005
R13291 VSS.n2766 VSS.n2770 4.57324
R13292 VSS.n2762 VSS.n2760 0.147342
R13293 VSS.n2763 VSS.n2764 0.0732424
R13294 VSS.n2764 VSS.n2765 0.147342
R13295 VSS.n2767 VSS.n2771 0.0721009
R13296 VSS.n2772 VSS.n2768 4.5005
R13297 VSS.n2773 VSS.n2769 4.5005
R13298 VSS.n2774 VSS.n2770 4.5005
R13299 VSS.n2760 VSS.n2771 4.57442
R13300 VSS.n2767 VSS.n2768 0.147342
R13301 VSS.n2768 VSS.n2769 0.147342
R13302 VSS.n2769 VSS.n2770 0.147342
R13303 VSS.n2771 VSS.n2772 2.39784
R13304 VSS.n2772 VSS.n2773 0.147342
R13305 VSS.n2773 VSS.n2774 0.147342
R13306 VSS.n2774 VSS.t165 3.13212
R13307 VSS.n2747 VSS.n2752 4.5005
R13308 VSS.n2749 VSS.n2753 4.5005
R13309 VSS.n2750 VSS.n2754 4.5005
R13310 VSS.n2751 VSS.n2755 4.57324
R13311 VSS.n2747 VSS.n2745 0.147342
R13312 VSS.n2748 VSS.n2749 0.0732424
R13313 VSS.n2749 VSS.n2750 0.147342
R13314 VSS.n2752 VSS.n2756 0.0721009
R13315 VSS.n2757 VSS.n2753 4.5005
R13316 VSS.n2758 VSS.n2754 4.5005
R13317 VSS.n2759 VSS.n2755 4.5005
R13318 VSS.n2745 VSS.n2756 4.57442
R13319 VSS.n2752 VSS.n2753 0.147342
R13320 VSS.n2753 VSS.n2754 0.147342
R13321 VSS.n2754 VSS.n2755 0.147342
R13322 VSS.n2756 VSS.n2757 2.39784
R13323 VSS.n2757 VSS.n2758 0.147342
R13324 VSS.n2758 VSS.n2759 0.147342
R13325 VSS.n2759 VSS.t128 3.13212
R13326 VSS.n2732 VSS.n2737 4.5005
R13327 VSS.n2734 VSS.n2738 4.5005
R13328 VSS.n2735 VSS.n2739 4.5005
R13329 VSS.n2736 VSS.n2740 4.57324
R13330 VSS.n2732 VSS.n2730 0.147342
R13331 VSS.n2733 VSS.n2734 0.0732424
R13332 VSS.n2734 VSS.n2735 0.147342
R13333 VSS.n2737 VSS.n2741 0.0721009
R13334 VSS.n2742 VSS.n2738 4.5005
R13335 VSS.n2743 VSS.n2739 4.5005
R13336 VSS.n2744 VSS.n2740 4.5005
R13337 VSS.n2730 VSS.n2741 4.57442
R13338 VSS.n2737 VSS.n2738 0.147342
R13339 VSS.n2738 VSS.n2739 0.147342
R13340 VSS.n2739 VSS.n2740 0.147342
R13341 VSS.n2741 VSS.n2742 2.39784
R13342 VSS.n2742 VSS.n2743 0.147342
R13343 VSS.n2743 VSS.n2744 0.147342
R13344 VSS.n2744 VSS.t19 3.13212
R13345 VSS.n2722 VSS.n2717 4.5005
R13346 VSS.n2723 VSS.n2719 4.5005
R13347 VSS.n2724 VSS.n2720 4.5005
R13348 VSS.n2725 VSS.n2721 4.57324
R13349 VSS.n2715 VSS.n2717 0.147342
R13350 VSS.n2718 VSS.n2719 0.0732424
R13351 VSS.n2719 VSS.n2720 0.147342
R13352 VSS.n2726 VSS.n2722 0.0722544
R13353 VSS.n2727 VSS.n2723 4.5005
R13354 VSS.n2728 VSS.n2724 4.5005
R13355 VSS.n2729 VSS.n2725 4.5005
R13356 VSS.n2726 VSS.n2715 4.57426
R13357 VSS.n2722 VSS.n2723 0.147342
R13358 VSS.n2723 VSS.n2724 0.147342
R13359 VSS.n2724 VSS.n2725 0.147342
R13360 VSS.n2727 VSS.n2726 2.37296
R13361 VSS.n2728 VSS.n2727 0.127318
R13362 VSS.n2729 VSS.n2728 0.127318
R13363 VSS.t5 VSS.n2729 2.73618
R13364 VSS.n2702 VSS.n2707 4.5005
R13365 VSS.n2704 VSS.n2708 4.5005
R13366 VSS.n2705 VSS.n2709 4.5005
R13367 VSS.n2706 VSS.n2710 4.57324
R13368 VSS.n2702 VSS.n2700 0.147342
R13369 VSS.n2703 VSS.n2704 0.0732424
R13370 VSS.n2704 VSS.n2705 0.147342
R13371 VSS.n2707 VSS.n2711 0.0721009
R13372 VSS.n2712 VSS.n2708 4.5005
R13373 VSS.n2713 VSS.n2709 4.5005
R13374 VSS.n2714 VSS.n2710 4.5005
R13375 VSS.n2700 VSS.n2711 4.57442
R13376 VSS.n2707 VSS.n2708 0.147342
R13377 VSS.n2708 VSS.n2709 0.147342
R13378 VSS.n2709 VSS.n2710 0.147342
R13379 VSS.n2711 VSS.n2712 2.39784
R13380 VSS.n2712 VSS.n2713 0.147342
R13381 VSS.n2713 VSS.n2714 0.147342
R13382 VSS.n2714 VSS.t232 3.13212
R13383 VSS.n2687 VSS.n2692 4.5005
R13384 VSS.n2689 VSS.n2693 4.5005
R13385 VSS.n2690 VSS.n2694 4.5005
R13386 VSS.n2691 VSS.n2695 4.57324
R13387 VSS.n2687 VSS.n2685 0.147342
R13388 VSS.n2688 VSS.n2689 0.0732424
R13389 VSS.n2689 VSS.n2690 0.147342
R13390 VSS.n2692 VSS.n2696 0.0721009
R13391 VSS.n2697 VSS.n2693 4.5005
R13392 VSS.n2698 VSS.n2694 4.5005
R13393 VSS.n2699 VSS.n2695 4.5005
R13394 VSS.n2685 VSS.n2696 4.57442
R13395 VSS.n2692 VSS.n2693 0.147342
R13396 VSS.n2693 VSS.n2694 0.147342
R13397 VSS.n2694 VSS.n2695 0.147342
R13398 VSS.n2696 VSS.n2697 2.39784
R13399 VSS.n2697 VSS.n2698 0.147342
R13400 VSS.n2698 VSS.n2699 0.147342
R13401 VSS.n2699 VSS.t466 3.13212
R13402 VSS.n2672 VSS.n2677 4.5005
R13403 VSS.n2674 VSS.n2678 4.5005
R13404 VSS.n2675 VSS.n2679 4.5005
R13405 VSS.n2676 VSS.n2680 4.57324
R13406 VSS.n2672 VSS.n2670 0.147342
R13407 VSS.n2673 VSS.n2674 0.0732424
R13408 VSS.n2674 VSS.n2675 0.147342
R13409 VSS.n2677 VSS.n2681 0.0721009
R13410 VSS.n2682 VSS.n2678 4.5005
R13411 VSS.n2683 VSS.n2679 4.5005
R13412 VSS.n2684 VSS.n2680 4.5005
R13413 VSS.n2670 VSS.n2681 4.57442
R13414 VSS.n2677 VSS.n2678 0.147342
R13415 VSS.n2678 VSS.n2679 0.147342
R13416 VSS.n2679 VSS.n2680 0.147342
R13417 VSS.n2681 VSS.n2682 2.39784
R13418 VSS.n2682 VSS.n2683 0.147342
R13419 VSS.n2683 VSS.n2684 0.147342
R13420 VSS.n2684 VSS.t243 3.13212
R13421 VSS.n2657 VSS.n2662 4.5005
R13422 VSS.n2659 VSS.n2663 4.5005
R13423 VSS.n2660 VSS.n2664 4.5005
R13424 VSS.n2661 VSS.n2665 4.57324
R13425 VSS.n2657 VSS.n2655 0.147342
R13426 VSS.n2658 VSS.n2659 0.0732424
R13427 VSS.n2659 VSS.n2660 0.147342
R13428 VSS.n2662 VSS.n2666 0.0721009
R13429 VSS.n2667 VSS.n2663 4.5005
R13430 VSS.n2668 VSS.n2664 4.5005
R13431 VSS.n2669 VSS.n2665 4.5005
R13432 VSS.n2655 VSS.n2666 4.57442
R13433 VSS.n2662 VSS.n2663 0.147342
R13434 VSS.n2663 VSS.n2664 0.147342
R13435 VSS.n2664 VSS.n2665 0.147342
R13436 VSS.n2666 VSS.n2667 2.39784
R13437 VSS.n2667 VSS.n2668 0.147342
R13438 VSS.n2668 VSS.n2669 0.147342
R13439 VSS.n2669 VSS.t345 3.13212
R13440 VSS.n2647 VSS.n2642 4.5005
R13441 VSS.n2648 VSS.n2644 4.5005
R13442 VSS.n2649 VSS.n2645 4.5005
R13443 VSS.n2650 VSS.n2646 4.57324
R13444 VSS.n2640 VSS.n2642 0.147342
R13445 VSS.n2643 VSS.n2644 0.0732424
R13446 VSS.n2644 VSS.n2645 0.147342
R13447 VSS.n2651 VSS.n2647 0.0722544
R13448 VSS.n2652 VSS.n2648 4.5005
R13449 VSS.n2653 VSS.n2649 4.5005
R13450 VSS.n2654 VSS.n2650 4.5005
R13451 VSS.n2651 VSS.n2640 4.57426
R13452 VSS.n2647 VSS.n2648 0.147342
R13453 VSS.n2648 VSS.n2649 0.147342
R13454 VSS.n2649 VSS.n2650 0.147342
R13455 VSS.n2652 VSS.n2651 2.37296
R13456 VSS.n2653 VSS.n2652 0.127318
R13457 VSS.n2654 VSS.n2653 0.127318
R13458 VSS.t5 VSS.n2654 2.73618
R13459 VSS.n2627 VSS.n2632 4.5005
R13460 VSS.n2629 VSS.n2633 4.5005
R13461 VSS.n2630 VSS.n2634 4.5005
R13462 VSS.n2631 VSS.n2635 4.57324
R13463 VSS.n2627 VSS.n2625 0.147342
R13464 VSS.n2628 VSS.n2629 0.0732424
R13465 VSS.n2629 VSS.n2630 0.147342
R13466 VSS.n2632 VSS.n2636 0.0721009
R13467 VSS.n2637 VSS.n2633 4.5005
R13468 VSS.n2638 VSS.n2634 4.5005
R13469 VSS.n2639 VSS.n2635 4.5005
R13470 VSS.n2625 VSS.n2636 4.57442
R13471 VSS.n2632 VSS.n2633 0.147342
R13472 VSS.n2633 VSS.n2634 0.147342
R13473 VSS.n2634 VSS.n2635 0.147342
R13474 VSS.n2636 VSS.n2637 2.39784
R13475 VSS.n2637 VSS.n2638 0.147342
R13476 VSS.n2638 VSS.n2639 0.147342
R13477 VSS.n2639 VSS.t436 3.13212
R13478 VSS.n2612 VSS.n2617 4.5005
R13479 VSS.n2614 VSS.n2618 4.5005
R13480 VSS.n2615 VSS.n2619 4.5005
R13481 VSS.n2616 VSS.n2620 4.57324
R13482 VSS.n2612 VSS.n2610 0.147342
R13483 VSS.n2613 VSS.n2614 0.0732424
R13484 VSS.n2614 VSS.n2615 0.147342
R13485 VSS.n2617 VSS.n2621 0.0721009
R13486 VSS.n2622 VSS.n2618 4.5005
R13487 VSS.n2623 VSS.n2619 4.5005
R13488 VSS.n2624 VSS.n2620 4.5005
R13489 VSS.n2610 VSS.n2621 4.57442
R13490 VSS.n2617 VSS.n2618 0.147342
R13491 VSS.n2618 VSS.n2619 0.147342
R13492 VSS.n2619 VSS.n2620 0.147342
R13493 VSS.n2621 VSS.n2622 2.39784
R13494 VSS.n2622 VSS.n2623 0.147342
R13495 VSS.n2623 VSS.n2624 0.147342
R13496 VSS.n2624 VSS.t89 3.13212
R13497 VSS.n2597 VSS.n2602 4.5005
R13498 VSS.n2599 VSS.n2603 4.5005
R13499 VSS.n2600 VSS.n2604 4.5005
R13500 VSS.n2601 VSS.n2605 4.57324
R13501 VSS.n2597 VSS.n2595 0.147342
R13502 VSS.n2598 VSS.n2599 0.0732424
R13503 VSS.n2599 VSS.n2600 0.147342
R13504 VSS.n2602 VSS.n2606 0.0721009
R13505 VSS.n2607 VSS.n2603 4.5005
R13506 VSS.n2608 VSS.n2604 4.5005
R13507 VSS.n2609 VSS.n2605 4.5005
R13508 VSS.n2595 VSS.n2606 4.57442
R13509 VSS.n2602 VSS.n2603 0.147342
R13510 VSS.n2603 VSS.n2604 0.147342
R13511 VSS.n2604 VSS.n2605 0.147342
R13512 VSS.n2606 VSS.n2607 2.39784
R13513 VSS.n2607 VSS.n2608 0.147342
R13514 VSS.n2608 VSS.n2609 0.147342
R13515 VSS.n2609 VSS.t518 3.13212
R13516 VSS.n2587 VSS.n2582 4.5005
R13517 VSS.n2588 VSS.n2584 4.5005
R13518 VSS.n2589 VSS.n2585 4.5005
R13519 VSS.n2590 VSS.n2586 4.57324
R13520 VSS.n2580 VSS.n2582 0.147342
R13521 VSS.n2583 VSS.n2584 0.0732424
R13522 VSS.n2584 VSS.n2585 0.147342
R13523 VSS.n2591 VSS.n2587 0.0722544
R13524 VSS.n2592 VSS.n2588 4.5005
R13525 VSS.n2593 VSS.n2589 4.5005
R13526 VSS.n2594 VSS.n2590 4.5005
R13527 VSS.n2591 VSS.n2580 4.57426
R13528 VSS.n2587 VSS.n2588 0.147342
R13529 VSS.n2588 VSS.n2589 0.147342
R13530 VSS.n2589 VSS.n2590 0.147342
R13531 VSS.n2592 VSS.n2591 2.37296
R13532 VSS.n2593 VSS.n2592 0.127318
R13533 VSS.n2594 VSS.n2593 0.127318
R13534 VSS.t5 VSS.n2594 2.73618
R13535 VSS.n2567 VSS.n2572 4.5005
R13536 VSS.n2569 VSS.n2573 4.5005
R13537 VSS.n2570 VSS.n2574 4.5005
R13538 VSS.n2571 VSS.n2575 4.57324
R13539 VSS.n2567 VSS.n2565 0.147342
R13540 VSS.n2568 VSS.n2569 0.0732424
R13541 VSS.n2569 VSS.n2570 0.147342
R13542 VSS.n2572 VSS.n2576 0.0721009
R13543 VSS.n2577 VSS.n2573 4.5005
R13544 VSS.n2578 VSS.n2574 4.5005
R13545 VSS.n2579 VSS.n2575 4.5005
R13546 VSS.n2565 VSS.n2576 4.57442
R13547 VSS.n2572 VSS.n2573 0.147342
R13548 VSS.n2573 VSS.n2574 0.147342
R13549 VSS.n2574 VSS.n2575 0.147342
R13550 VSS.n2576 VSS.n2577 2.39784
R13551 VSS.n2577 VSS.n2578 0.147342
R13552 VSS.n2578 VSS.n2579 0.147342
R13553 VSS.n2579 VSS.t620 3.13212
R13554 VSS.n2552 VSS.n2557 4.5005
R13555 VSS.n2554 VSS.n2558 4.5005
R13556 VSS.n2555 VSS.n2559 4.5005
R13557 VSS.n2556 VSS.n2560 4.57324
R13558 VSS.n2552 VSS.n2550 0.147342
R13559 VSS.n2553 VSS.n2554 0.0732424
R13560 VSS.n2554 VSS.n2555 0.147342
R13561 VSS.n2557 VSS.n2561 0.0721009
R13562 VSS.n2562 VSS.n2558 4.5005
R13563 VSS.n2563 VSS.n2559 4.5005
R13564 VSS.n2564 VSS.n2560 4.5005
R13565 VSS.n2550 VSS.n2561 4.57442
R13566 VSS.n2557 VSS.n2558 0.147342
R13567 VSS.n2558 VSS.n2559 0.147342
R13568 VSS.n2559 VSS.n2560 0.147342
R13569 VSS.n2561 VSS.n2562 2.39784
R13570 VSS.n2562 VSS.n2563 0.147342
R13571 VSS.n2563 VSS.n2564 0.147342
R13572 VSS.n2564 VSS.t185 3.13212
R13573 VSS.n2537 VSS.n2542 4.5005
R13574 VSS.n2539 VSS.n2543 4.5005
R13575 VSS.n2540 VSS.n2544 4.5005
R13576 VSS.n2541 VSS.n2545 4.57324
R13577 VSS.n2537 VSS.n2535 0.147342
R13578 VSS.n2538 VSS.n2539 0.0732424
R13579 VSS.n2539 VSS.n2540 0.147342
R13580 VSS.n2542 VSS.n2546 0.0721009
R13581 VSS.n2547 VSS.n2543 4.5005
R13582 VSS.n2548 VSS.n2544 4.5005
R13583 VSS.n2549 VSS.n2545 4.5005
R13584 VSS.n2535 VSS.n2546 4.57442
R13585 VSS.n2542 VSS.n2543 0.147342
R13586 VSS.n2543 VSS.n2544 0.147342
R13587 VSS.n2544 VSS.n2545 0.147342
R13588 VSS.n2546 VSS.n2547 2.39784
R13589 VSS.n2547 VSS.n2548 0.147342
R13590 VSS.n2548 VSS.n2549 0.147342
R13591 VSS.n2549 VSS.t145 3.13212
R13592 VSS.n2522 VSS.n2527 4.5005
R13593 VSS.n2524 VSS.n2528 4.5005
R13594 VSS.n2525 VSS.n2529 4.5005
R13595 VSS.n2526 VSS.n2530 4.57324
R13596 VSS.n2522 VSS.n2520 0.147342
R13597 VSS.n2523 VSS.n2524 0.0732424
R13598 VSS.n2524 VSS.n2525 0.147342
R13599 VSS.n2527 VSS.n2531 0.0721009
R13600 VSS.n2532 VSS.n2528 4.5005
R13601 VSS.n2533 VSS.n2529 4.5005
R13602 VSS.n2534 VSS.n2530 4.5005
R13603 VSS.n2520 VSS.n2531 4.57442
R13604 VSS.n2527 VSS.n2528 0.147342
R13605 VSS.n2528 VSS.n2529 0.147342
R13606 VSS.n2529 VSS.n2530 0.147342
R13607 VSS.n2531 VSS.n2532 2.39784
R13608 VSS.n2532 VSS.n2533 0.147342
R13609 VSS.n2533 VSS.n2534 0.147342
R13610 VSS.n2534 VSS.t6 3.13212
R13611 VSS.n2507 VSS.n2512 4.5005
R13612 VSS.n2509 VSS.n2513 4.5005
R13613 VSS.n2510 VSS.n2514 4.5005
R13614 VSS.n2511 VSS.n2515 4.57324
R13615 VSS.n2507 VSS.n2505 0.147342
R13616 VSS.n2508 VSS.n2509 0.0732424
R13617 VSS.n2509 VSS.n2510 0.147342
R13618 VSS.n2512 VSS.n2516 0.0721009
R13619 VSS.n2517 VSS.n2513 4.5005
R13620 VSS.n2518 VSS.n2514 4.5005
R13621 VSS.n2519 VSS.n2515 4.5005
R13622 VSS.n2505 VSS.n2516 4.57442
R13623 VSS.n2512 VSS.n2513 0.147342
R13624 VSS.n2513 VSS.n2514 0.147342
R13625 VSS.n2514 VSS.n2515 0.147342
R13626 VSS.n2516 VSS.n2517 2.39784
R13627 VSS.n2517 VSS.n2518 0.147342
R13628 VSS.n2518 VSS.n2519 0.147342
R13629 VSS.n2519 VSS.t197 3.13212
R13630 VSS.n2492 VSS.n2497 4.5005
R13631 VSS.n2494 VSS.n2498 4.5005
R13632 VSS.n2495 VSS.n2499 4.5005
R13633 VSS.n2496 VSS.n2500 4.57324
R13634 VSS.n2492 VSS.n2490 0.147342
R13635 VSS.n2493 VSS.n2494 0.0732424
R13636 VSS.n2494 VSS.n2495 0.147342
R13637 VSS.n2497 VSS.n2501 0.0721009
R13638 VSS.n2502 VSS.n2498 4.5005
R13639 VSS.n2503 VSS.n2499 4.5005
R13640 VSS.n2504 VSS.n2500 4.5005
R13641 VSS.n2490 VSS.n2501 4.57442
R13642 VSS.n2497 VSS.n2498 0.147342
R13643 VSS.n2498 VSS.n2499 0.147342
R13644 VSS.n2499 VSS.n2500 0.147342
R13645 VSS.n2501 VSS.n2502 2.39784
R13646 VSS.n2502 VSS.n2503 0.147342
R13647 VSS.n2503 VSS.n2504 0.147342
R13648 VSS.n2504 VSS.t169 3.13212
R13649 VSS.n2482 VSS.n2477 4.5005
R13650 VSS.n2483 VSS.n2479 4.5005
R13651 VSS.n2484 VSS.n2480 4.5005
R13652 VSS.n2485 VSS.n2481 4.57324
R13653 VSS.n2475 VSS.n2477 0.147342
R13654 VSS.n2478 VSS.n2479 0.0732424
R13655 VSS.n2479 VSS.n2480 0.147342
R13656 VSS.n2486 VSS.n2482 0.0722544
R13657 VSS.n2487 VSS.n2483 4.5005
R13658 VSS.n2488 VSS.n2484 4.5005
R13659 VSS.n2489 VSS.n2485 4.5005
R13660 VSS.n2486 VSS.n2475 4.57426
R13661 VSS.n2482 VSS.n2483 0.147342
R13662 VSS.n2483 VSS.n2484 0.147342
R13663 VSS.n2484 VSS.n2485 0.147342
R13664 VSS.n2487 VSS.n2486 2.37296
R13665 VSS.n2488 VSS.n2487 0.127318
R13666 VSS.n2489 VSS.n2488 0.127318
R13667 VSS.t5 VSS.n2489 2.73618
R13668 VSS.n2462 VSS.n2467 4.5005
R13669 VSS.n2464 VSS.n2468 4.5005
R13670 VSS.n2465 VSS.n2469 4.5005
R13671 VSS.n2466 VSS.n2470 4.57324
R13672 VSS.n2462 VSS.n2460 0.147342
R13673 VSS.n2463 VSS.n2464 0.0732424
R13674 VSS.n2464 VSS.n2465 0.147342
R13675 VSS.n2467 VSS.n2471 0.0721009
R13676 VSS.n2472 VSS.n2468 4.5005
R13677 VSS.n2473 VSS.n2469 4.5005
R13678 VSS.n2474 VSS.n2470 4.5005
R13679 VSS.n2460 VSS.n2471 4.57442
R13680 VSS.n2467 VSS.n2468 0.147342
R13681 VSS.n2468 VSS.n2469 0.147342
R13682 VSS.n2469 VSS.n2470 0.147342
R13683 VSS.n2471 VSS.n2472 2.39784
R13684 VSS.n2472 VSS.n2473 0.147342
R13685 VSS.n2473 VSS.n2474 0.147342
R13686 VSS.n2474 VSS.t365 3.13212
R13687 VSS.n2447 VSS.n2452 4.5005
R13688 VSS.n2449 VSS.n2453 4.5005
R13689 VSS.n2450 VSS.n2454 4.5005
R13690 VSS.n2451 VSS.n2455 4.57324
R13691 VSS.n2447 VSS.n2445 0.147342
R13692 VSS.n2448 VSS.n2449 0.0732424
R13693 VSS.n2449 VSS.n2450 0.147342
R13694 VSS.n2452 VSS.n2456 0.0721009
R13695 VSS.n2457 VSS.n2453 4.5005
R13696 VSS.n2458 VSS.n2454 4.5005
R13697 VSS.n2459 VSS.n2455 4.5005
R13698 VSS.n2445 VSS.n2456 4.57442
R13699 VSS.n2452 VSS.n2453 0.147342
R13700 VSS.n2453 VSS.n2454 0.147342
R13701 VSS.n2454 VSS.n2455 0.147342
R13702 VSS.n2456 VSS.n2457 2.39784
R13703 VSS.n2457 VSS.n2458 0.147342
R13704 VSS.n2458 VSS.n2459 0.147342
R13705 VSS.n2459 VSS.t126 3.13212
R13706 VSS.n2432 VSS.n2437 4.5005
R13707 VSS.n2434 VSS.n2438 4.5005
R13708 VSS.n2435 VSS.n2439 4.5005
R13709 VSS.n2436 VSS.n2440 4.57324
R13710 VSS.n2432 VSS.n2430 0.147342
R13711 VSS.n2433 VSS.n2434 0.0732424
R13712 VSS.n2434 VSS.n2435 0.147342
R13713 VSS.n2437 VSS.n2441 0.0721009
R13714 VSS.n2442 VSS.n2438 4.5005
R13715 VSS.n2443 VSS.n2439 4.5005
R13716 VSS.n2444 VSS.n2440 4.5005
R13717 VSS.n2430 VSS.n2441 4.57442
R13718 VSS.n2437 VSS.n2438 0.147342
R13719 VSS.n2438 VSS.n2439 0.147342
R13720 VSS.n2439 VSS.n2440 0.147342
R13721 VSS.n2441 VSS.n2442 2.39784
R13722 VSS.n2442 VSS.n2443 0.147342
R13723 VSS.n2443 VSS.n2444 0.147342
R13724 VSS.n2444 VSS.t29 3.13212
R13725 VSS.n2422 VSS.n2417 4.5005
R13726 VSS.n2423 VSS.n2419 4.5005
R13727 VSS.n2424 VSS.n2420 4.5005
R13728 VSS.n2425 VSS.n2421 4.57324
R13729 VSS.n2415 VSS.n2417 0.147342
R13730 VSS.n2418 VSS.n2419 0.0732424
R13731 VSS.n2419 VSS.n2420 0.147342
R13732 VSS.n2426 VSS.n2422 0.0722544
R13733 VSS.n2427 VSS.n2423 4.5005
R13734 VSS.n2428 VSS.n2424 4.5005
R13735 VSS.n2429 VSS.n2425 4.5005
R13736 VSS.n2426 VSS.n2415 4.57426
R13737 VSS.n2422 VSS.n2423 0.147342
R13738 VSS.n2423 VSS.n2424 0.147342
R13739 VSS.n2424 VSS.n2425 0.147342
R13740 VSS.n2427 VSS.n2426 2.37296
R13741 VSS.n2428 VSS.n2427 0.127318
R13742 VSS.n2429 VSS.n2428 0.127318
R13743 VSS.t5 VSS.n2429 2.73618
R13744 VSS.n2402 VSS.n2407 4.5005
R13745 VSS.n2404 VSS.n2408 4.5005
R13746 VSS.n2405 VSS.n2409 4.5005
R13747 VSS.n2406 VSS.n2410 4.57324
R13748 VSS.n2402 VSS.n2400 0.147342
R13749 VSS.n2403 VSS.n2404 0.0732424
R13750 VSS.n2404 VSS.n2405 0.147342
R13751 VSS.n2407 VSS.n2411 0.0721009
R13752 VSS.n2412 VSS.n2408 4.5005
R13753 VSS.n2413 VSS.n2409 4.5005
R13754 VSS.n2414 VSS.n2410 4.5005
R13755 VSS.n2400 VSS.n2411 4.57442
R13756 VSS.n2407 VSS.n2408 0.147342
R13757 VSS.n2408 VSS.n2409 0.147342
R13758 VSS.n2409 VSS.n2410 0.147342
R13759 VSS.n2411 VSS.n2412 2.39784
R13760 VSS.n2412 VSS.n2413 0.147342
R13761 VSS.n2413 VSS.n2414 0.147342
R13762 VSS.n2414 VSS.t330 3.13212
R13763 VSS.n2387 VSS.n2392 4.5005
R13764 VSS.n2389 VSS.n2393 4.5005
R13765 VSS.n2390 VSS.n2394 4.5005
R13766 VSS.n2391 VSS.n2395 4.57324
R13767 VSS.n2387 VSS.n2385 0.147342
R13768 VSS.n2388 VSS.n2389 0.0732424
R13769 VSS.n2389 VSS.n2390 0.147342
R13770 VSS.n2392 VSS.n2396 0.0721009
R13771 VSS.n2397 VSS.n2393 4.5005
R13772 VSS.n2398 VSS.n2394 4.5005
R13773 VSS.n2399 VSS.n2395 4.5005
R13774 VSS.n2385 VSS.n2396 4.57442
R13775 VSS.n2392 VSS.n2393 0.147342
R13776 VSS.n2393 VSS.n2394 0.147342
R13777 VSS.n2394 VSS.n2395 0.147342
R13778 VSS.n2396 VSS.n2397 2.39784
R13779 VSS.n2397 VSS.n2398 0.147342
R13780 VSS.n2398 VSS.n2399 0.147342
R13781 VSS.n2399 VSS.t490 3.13212
R13782 VSS.n2361 VSS.n2362 0.0722544
R13783 VSS.n2363 VSS.n2364 4.5005
R13784 VSS.n2365 VSS.n2366 4.5005
R13785 VSS.n2367 VSS.n2368 4.5005
R13786 VSS.n2363 VSS.n2361 2.37296
R13787 VSS.n2365 VSS.n2363 0.127318
R13788 VSS.n2367 VSS.n2365 0.127318
R13789 VSS.t20 VSS.n2367 2.73618
R13790 VSS.n2362 VSS.n2027 4.5005
R13791 VSS.n2364 VSS.n2029 4.5005
R13792 VSS.n2366 VSS.n2030 4.5005
R13793 VSS.n2361 VSS.n2025 4.57426
R13794 VSS.n2362 VSS.n2364 0.147342
R13795 VSS.n2364 VSS.n2366 0.147342
R13796 VSS.n2366 VSS.n2368 0.147342
R13797 VSS.n2025 VSS.n2027 0.147342
R13798 VSS.n2028 VSS.n2029 0.0732424
R13799 VSS.n2029 VSS.n2030 0.147342
R13800 VSS.n2030 VSS.n2369 0.0732424
R13801 VSS.n2353 VSS.n2352 0.0722544
R13802 VSS.n2354 VSS.n2355 4.5005
R13803 VSS.n2356 VSS.n2357 4.5005
R13804 VSS.n2358 VSS.n2359 4.5005
R13805 VSS.n2352 VSS.n2354 2.37296
R13806 VSS.n2354 VSS.n2356 0.127318
R13807 VSS.n2356 VSS.n2358 0.127318
R13808 VSS.n2358 VSS.t20 2.73618
R13809 VSS.n1931 VSS.n2353 4.5005
R13810 VSS.n1933 VSS.n2355 4.5005
R13811 VSS.n1934 VSS.n2357 4.5005
R13812 VSS.n1929 VSS.n2352 4.57426
R13813 VSS.n2353 VSS.n2355 0.147342
R13814 VSS.n2355 VSS.n2357 0.147342
R13815 VSS.n2357 VSS.n2359 0.147342
R13816 VSS.n1931 VSS.n1929 0.147342
R13817 VSS.n1932 VSS.n1933 0.0732424
R13818 VSS.n1933 VSS.n1934 0.147342
R13819 VSS.n2360 VSS.n1934 0.0732424
R13820 VSS.n2344 VSS.n2343 0.0722544
R13821 VSS.n2345 VSS.n2346 4.5005
R13822 VSS.n2347 VSS.n2348 4.5005
R13823 VSS.n2349 VSS.n2350 4.5005
R13824 VSS.n2343 VSS.n2345 2.37296
R13825 VSS.n2345 VSS.n2347 0.127318
R13826 VSS.n2347 VSS.n2349 0.127318
R13827 VSS.n2349 VSS.t20 2.73618
R13828 VSS.n1880 VSS.n2344 4.5005
R13829 VSS.n1882 VSS.n2346 4.5005
R13830 VSS.n1883 VSS.n2348 4.5005
R13831 VSS.n1878 VSS.n2343 4.57426
R13832 VSS.n2344 VSS.n2346 0.147342
R13833 VSS.n2346 VSS.n2348 0.147342
R13834 VSS.n2348 VSS.n2350 0.147342
R13835 VSS.n1880 VSS.n1878 0.147342
R13836 VSS.n1881 VSS.n1882 0.0732424
R13837 VSS.n1882 VSS.n1883 0.147342
R13838 VSS.n2351 VSS.n1883 0.0732424
R13839 VSS.n2335 VSS.n2334 0.0722544
R13840 VSS.n2336 VSS.n2337 4.5005
R13841 VSS.n2338 VSS.n2339 4.5005
R13842 VSS.n2340 VSS.n2341 4.5005
R13843 VSS.n2334 VSS.n2336 2.37296
R13844 VSS.n2336 VSS.n2338 0.127318
R13845 VSS.n2338 VSS.n2340 0.127318
R13846 VSS.n2340 VSS.t20 2.73618
R13847 VSS.n1814 VSS.n2335 4.5005
R13848 VSS.n1816 VSS.n2337 4.5005
R13849 VSS.n1817 VSS.n2339 4.5005
R13850 VSS.n1812 VSS.n2334 4.57426
R13851 VSS.n2335 VSS.n2337 0.147342
R13852 VSS.n2337 VSS.n2339 0.147342
R13853 VSS.n2339 VSS.n2341 0.147342
R13854 VSS.n1814 VSS.n1812 0.147342
R13855 VSS.n1815 VSS.n1816 0.0732424
R13856 VSS.n1816 VSS.n1817 0.147342
R13857 VSS.n2342 VSS.n1817 0.0732424
R13858 VSS.n2326 VSS.n2325 0.0722544
R13859 VSS.n2327 VSS.n2328 4.5005
R13860 VSS.n2329 VSS.n2330 4.5005
R13861 VSS.n2331 VSS.n2332 4.5005
R13862 VSS.n2325 VSS.n2327 2.37296
R13863 VSS.n2327 VSS.n2329 0.127318
R13864 VSS.n2329 VSS.n2331 0.127318
R13865 VSS.n2331 VSS.t20 2.73618
R13866 VSS.n1763 VSS.n2326 4.5005
R13867 VSS.n1765 VSS.n2328 4.5005
R13868 VSS.n1766 VSS.n2330 4.5005
R13869 VSS.n1761 VSS.n2325 4.57426
R13870 VSS.n2326 VSS.n2328 0.147342
R13871 VSS.n2328 VSS.n2330 0.147342
R13872 VSS.n2330 VSS.n2332 0.147342
R13873 VSS.n1763 VSS.n1761 0.147342
R13874 VSS.n1764 VSS.n1765 0.0732424
R13875 VSS.n1765 VSS.n1766 0.147342
R13876 VSS.n2333 VSS.n1766 0.0732424
R13877 VSS.n2317 VSS.n2316 0.0722544
R13878 VSS.n2318 VSS.n2319 4.5005
R13879 VSS.n2320 VSS.n2321 4.5005
R13880 VSS.n2322 VSS.n2323 4.5005
R13881 VSS.n2316 VSS.n2318 2.37296
R13882 VSS.n2318 VSS.n2320 0.127318
R13883 VSS.n2320 VSS.n2322 0.127318
R13884 VSS.n2322 VSS.t20 2.73618
R13885 VSS.n1667 VSS.n2317 4.5005
R13886 VSS.n1669 VSS.n2319 4.5005
R13887 VSS.n1670 VSS.n2321 4.5005
R13888 VSS.n1665 VSS.n2316 4.57426
R13889 VSS.n2317 VSS.n2319 0.147342
R13890 VSS.n2319 VSS.n2321 0.147342
R13891 VSS.n2321 VSS.n2323 0.147342
R13892 VSS.n1667 VSS.n1665 0.147342
R13893 VSS.n1668 VSS.n1669 0.0732424
R13894 VSS.n1669 VSS.n1670 0.147342
R13895 VSS.n2324 VSS.n1670 0.0732424
R13896 VSS.n2308 VSS.n2307 0.0722544
R13897 VSS.n2309 VSS.n2310 4.5005
R13898 VSS.n2311 VSS.n2312 4.5005
R13899 VSS.n2313 VSS.n2314 4.5005
R13900 VSS.n2307 VSS.n2309 2.37296
R13901 VSS.n2309 VSS.n2311 0.127318
R13902 VSS.n2311 VSS.n2313 0.127318
R13903 VSS.n2313 VSS.t20 2.73618
R13904 VSS.n1616 VSS.n2308 4.5005
R13905 VSS.n1618 VSS.n2310 4.5005
R13906 VSS.n1619 VSS.n2312 4.5005
R13907 VSS.n1614 VSS.n2307 4.57426
R13908 VSS.n2308 VSS.n2310 0.147342
R13909 VSS.n2310 VSS.n2312 0.147342
R13910 VSS.n2312 VSS.n2314 0.147342
R13911 VSS.n1616 VSS.n1614 0.147342
R13912 VSS.n1617 VSS.n1618 0.0732424
R13913 VSS.n1618 VSS.n1619 0.147342
R13914 VSS.n2315 VSS.n1619 0.0732424
R13915 VSS.n2299 VSS.n2298 0.0722544
R13916 VSS.n2300 VSS.n2301 4.5005
R13917 VSS.n2302 VSS.n2303 4.5005
R13918 VSS.n2304 VSS.n2305 4.5005
R13919 VSS.n2298 VSS.n2300 2.37296
R13920 VSS.n2300 VSS.n2302 0.127318
R13921 VSS.n2302 VSS.n2304 0.127318
R13922 VSS.n2304 VSS.t20 2.73618
R13923 VSS.n1550 VSS.n2299 4.5005
R13924 VSS.n1552 VSS.n2301 4.5005
R13925 VSS.n1553 VSS.n2303 4.5005
R13926 VSS.n1548 VSS.n2298 4.57426
R13927 VSS.n2299 VSS.n2301 0.147342
R13928 VSS.n2301 VSS.n2303 0.147342
R13929 VSS.n2303 VSS.n2305 0.147342
R13930 VSS.n1550 VSS.n1548 0.147342
R13931 VSS.n1551 VSS.n1552 0.0732424
R13932 VSS.n1552 VSS.n1553 0.147342
R13933 VSS.n2306 VSS.n1553 0.0732424
R13934 VSS.n2290 VSS.n2289 0.0722544
R13935 VSS.n2291 VSS.n2292 4.5005
R13936 VSS.n2293 VSS.n2294 4.5005
R13937 VSS.n2295 VSS.n2296 4.5005
R13938 VSS.n2289 VSS.n2291 2.37296
R13939 VSS.n2291 VSS.n2293 0.127318
R13940 VSS.n2293 VSS.n2295 0.127318
R13941 VSS.n2295 VSS.t20 2.73618
R13942 VSS.n1499 VSS.n2290 4.5005
R13943 VSS.n1501 VSS.n2292 4.5005
R13944 VSS.n1502 VSS.n2294 4.5005
R13945 VSS.n1497 VSS.n2289 4.57426
R13946 VSS.n2290 VSS.n2292 0.147342
R13947 VSS.n2292 VSS.n2294 0.147342
R13948 VSS.n2294 VSS.n2296 0.147342
R13949 VSS.n1499 VSS.n1497 0.147342
R13950 VSS.n1500 VSS.n1501 0.0732424
R13951 VSS.n1501 VSS.n1502 0.147342
R13952 VSS.n2297 VSS.n1502 0.0732424
R13953 VSS.n2280 VSS.n2281 0.0722544
R13954 VSS.n2282 VSS.n2283 4.5005
R13955 VSS.n2284 VSS.n2285 4.5005
R13956 VSS.n2286 VSS.n2287 4.5005
R13957 VSS.n2282 VSS.n2280 2.37296
R13958 VSS.n2284 VSS.n2282 0.127318
R13959 VSS.n2286 VSS.n2284 0.127318
R13960 VSS.t20 VSS.n2286 2.73618
R13961 VSS.n2281 VSS.n1403 4.5005
R13962 VSS.n2283 VSS.n1405 4.5005
R13963 VSS.n2285 VSS.n1406 4.5005
R13964 VSS.n2280 VSS.n1401 4.57426
R13965 VSS.n2281 VSS.n2283 0.147342
R13966 VSS.n2283 VSS.n2285 0.147342
R13967 VSS.n2285 VSS.n2287 0.147342
R13968 VSS.n1401 VSS.n1403 0.147342
R13969 VSS.n1404 VSS.n1405 0.0732424
R13970 VSS.n1405 VSS.n1406 0.147342
R13971 VSS.n1406 VSS.n2288 0.0732424
R13972 VSS.n2271 VSS.n2272 0.0722544
R13973 VSS.n2273 VSS.n2274 4.5005
R13974 VSS.n2275 VSS.n2276 4.5005
R13975 VSS.n2277 VSS.n2278 4.5005
R13976 VSS.n2273 VSS.n2271 2.37296
R13977 VSS.n2275 VSS.n2273 0.127318
R13978 VSS.n2277 VSS.n2275 0.127318
R13979 VSS.t20 VSS.n2277 2.73618
R13980 VSS.n2272 VSS.n1352 4.5005
R13981 VSS.n2274 VSS.n1354 4.5005
R13982 VSS.n2276 VSS.n1355 4.5005
R13983 VSS.n2271 VSS.n1350 4.57426
R13984 VSS.n2272 VSS.n2274 0.147342
R13985 VSS.n2274 VSS.n2276 0.147342
R13986 VSS.n2276 VSS.n2278 0.147342
R13987 VSS.n1350 VSS.n1352 0.147342
R13988 VSS.n1353 VSS.n1354 0.0732424
R13989 VSS.n1354 VSS.n1355 0.147342
R13990 VSS.n1355 VSS.n2279 0.0732424
R13991 VSS.n2262 VSS.n2263 0.0722544
R13992 VSS.n2264 VSS.n2265 4.5005
R13993 VSS.n2266 VSS.n2267 4.5005
R13994 VSS.n2268 VSS.n2269 4.5005
R13995 VSS.n2264 VSS.n2262 2.37296
R13996 VSS.n2266 VSS.n2264 0.127318
R13997 VSS.n2268 VSS.n2266 0.127318
R13998 VSS.t20 VSS.n2268 2.73618
R13999 VSS.n2263 VSS.n1286 4.5005
R14000 VSS.n2265 VSS.n1288 4.5005
R14001 VSS.n2267 VSS.n1289 4.5005
R14002 VSS.n2262 VSS.n1284 4.57426
R14003 VSS.n2263 VSS.n2265 0.147342
R14004 VSS.n2265 VSS.n2267 0.147342
R14005 VSS.n2267 VSS.n2269 0.147342
R14006 VSS.n1284 VSS.n1286 0.147342
R14007 VSS.n1287 VSS.n1288 0.0732424
R14008 VSS.n1288 VSS.n1289 0.147342
R14009 VSS.n1289 VSS.n2270 0.0732424
R14010 VSS.n2253 VSS.n2254 0.0722544
R14011 VSS.n2255 VSS.n2256 4.5005
R14012 VSS.n2257 VSS.n2258 4.5005
R14013 VSS.n2259 VSS.n2260 4.5005
R14014 VSS.n2255 VSS.n2253 2.37296
R14015 VSS.n2257 VSS.n2255 0.127318
R14016 VSS.n2259 VSS.n2257 0.127318
R14017 VSS.t20 VSS.n2259 2.73618
R14018 VSS.n2254 VSS.n1235 4.5005
R14019 VSS.n2256 VSS.n1237 4.5005
R14020 VSS.n2258 VSS.n1238 4.5005
R14021 VSS.n2253 VSS.n1233 4.57426
R14022 VSS.n2254 VSS.n2256 0.147342
R14023 VSS.n2256 VSS.n2258 0.147342
R14024 VSS.n2258 VSS.n2260 0.147342
R14025 VSS.n1233 VSS.n1235 0.147342
R14026 VSS.n1236 VSS.n1237 0.0732424
R14027 VSS.n1237 VSS.n1238 0.147342
R14028 VSS.n1238 VSS.n2261 0.0732424
R14029 VSS.n2244 VSS.n2245 0.0722544
R14030 VSS.n2246 VSS.n2247 4.5005
R14031 VSS.n2248 VSS.n2249 4.5005
R14032 VSS.n2250 VSS.n2251 4.5005
R14033 VSS.n2246 VSS.n2244 2.37296
R14034 VSS.n2248 VSS.n2246 0.127318
R14035 VSS.n2250 VSS.n2248 0.127318
R14036 VSS.t20 VSS.n2250 2.73618
R14037 VSS.n2245 VSS.n1139 4.5005
R14038 VSS.n2247 VSS.n1141 4.5005
R14039 VSS.n2249 VSS.n1142 4.5005
R14040 VSS.n2244 VSS.n1137 4.57426
R14041 VSS.n2245 VSS.n2247 0.147342
R14042 VSS.n2247 VSS.n2249 0.147342
R14043 VSS.n2249 VSS.n2251 0.147342
R14044 VSS.n1137 VSS.n1139 0.147342
R14045 VSS.n1140 VSS.n1141 0.0732424
R14046 VSS.n1141 VSS.n1142 0.147342
R14047 VSS.n1142 VSS.n2252 0.0732424
R14048 VSS.n2235 VSS.n2236 0.0722544
R14049 VSS.n2237 VSS.n2238 4.5005
R14050 VSS.n2239 VSS.n2240 4.5005
R14051 VSS.n2241 VSS.n2242 4.5005
R14052 VSS.n2237 VSS.n2235 2.37296
R14053 VSS.n2239 VSS.n2237 0.127318
R14054 VSS.n2241 VSS.n2239 0.127318
R14055 VSS.t20 VSS.n2241 2.73618
R14056 VSS.n2236 VSS.n1088 4.5005
R14057 VSS.n2238 VSS.n1090 4.5005
R14058 VSS.n2240 VSS.n1091 4.5005
R14059 VSS.n2235 VSS.n1086 4.57426
R14060 VSS.n2236 VSS.n2238 0.147342
R14061 VSS.n2238 VSS.n2240 0.147342
R14062 VSS.n2240 VSS.n2242 0.147342
R14063 VSS.n1086 VSS.n1088 0.147342
R14064 VSS.n1089 VSS.n1090 0.0732424
R14065 VSS.n1090 VSS.n1091 0.147342
R14066 VSS.n1091 VSS.n2243 0.0732424
R14067 VSS.n2226 VSS.n2227 0.0722544
R14068 VSS.n2228 VSS.n2229 4.5005
R14069 VSS.n2230 VSS.n2231 4.5005
R14070 VSS.n2232 VSS.n2233 4.5005
R14071 VSS.n2228 VSS.n2226 2.37296
R14072 VSS.n2230 VSS.n2228 0.127318
R14073 VSS.n2232 VSS.n2230 0.127318
R14074 VSS.t20 VSS.n2232 2.73618
R14075 VSS.n2227 VSS.n1022 4.5005
R14076 VSS.n2229 VSS.n1024 4.5005
R14077 VSS.n2231 VSS.n1025 4.5005
R14078 VSS.n2226 VSS.n1020 4.57426
R14079 VSS.n2227 VSS.n2229 0.147342
R14080 VSS.n2229 VSS.n2231 0.147342
R14081 VSS.n2231 VSS.n2233 0.147342
R14082 VSS.n1020 VSS.n1022 0.147342
R14083 VSS.n1023 VSS.n1024 0.0732424
R14084 VSS.n1024 VSS.n1025 0.147342
R14085 VSS.n1025 VSS.n2234 0.0732424
R14086 VSS.n2217 VSS.n2218 0.0722544
R14087 VSS.n2219 VSS.n2220 4.5005
R14088 VSS.n2221 VSS.n2222 4.5005
R14089 VSS.n2223 VSS.n2224 4.5005
R14090 VSS.n2219 VSS.n2217 2.37296
R14091 VSS.n2221 VSS.n2219 0.127318
R14092 VSS.n2223 VSS.n2221 0.127318
R14093 VSS.t20 VSS.n2223 2.73618
R14094 VSS.n2218 VSS.n971 4.5005
R14095 VSS.n2220 VSS.n973 4.5005
R14096 VSS.n2222 VSS.n974 4.5005
R14097 VSS.n2217 VSS.n969 4.57426
R14098 VSS.n2218 VSS.n2220 0.147342
R14099 VSS.n2220 VSS.n2222 0.147342
R14100 VSS.n2222 VSS.n2224 0.147342
R14101 VSS.n969 VSS.n971 0.147342
R14102 VSS.n972 VSS.n973 0.0732424
R14103 VSS.n973 VSS.n974 0.147342
R14104 VSS.n974 VSS.n2225 0.0732424
R14105 VSS.n2208 VSS.n2209 0.0722544
R14106 VSS.n2210 VSS.n2211 4.5005
R14107 VSS.n2212 VSS.n2213 4.5005
R14108 VSS.n2214 VSS.n2215 4.5005
R14109 VSS.n2210 VSS.n2208 2.37296
R14110 VSS.n2212 VSS.n2210 0.127318
R14111 VSS.n2214 VSS.n2212 0.127318
R14112 VSS.t20 VSS.n2214 2.73618
R14113 VSS.n2209 VSS.n875 4.5005
R14114 VSS.n2211 VSS.n877 4.5005
R14115 VSS.n2213 VSS.n878 4.5005
R14116 VSS.n2208 VSS.n873 4.57426
R14117 VSS.n2209 VSS.n2211 0.147342
R14118 VSS.n2211 VSS.n2213 0.147342
R14119 VSS.n2213 VSS.n2215 0.147342
R14120 VSS.n873 VSS.n875 0.147342
R14121 VSS.n876 VSS.n877 0.0732424
R14122 VSS.n877 VSS.n878 0.147342
R14123 VSS.n878 VSS.n2216 0.0732424
R14124 VSS.n2199 VSS.n2200 0.0722544
R14125 VSS.n2201 VSS.n2202 4.5005
R14126 VSS.n2203 VSS.n2204 4.5005
R14127 VSS.n2205 VSS.n2206 4.5005
R14128 VSS.n2201 VSS.n2199 2.37296
R14129 VSS.n2203 VSS.n2201 0.127318
R14130 VSS.n2205 VSS.n2203 0.127318
R14131 VSS.t20 VSS.n2205 2.73618
R14132 VSS.n2200 VSS.n824 4.5005
R14133 VSS.n2202 VSS.n826 4.5005
R14134 VSS.n2204 VSS.n827 4.5005
R14135 VSS.n2199 VSS.n822 4.57426
R14136 VSS.n2200 VSS.n2202 0.147342
R14137 VSS.n2202 VSS.n2204 0.147342
R14138 VSS.n2204 VSS.n2206 0.147342
R14139 VSS.n822 VSS.n824 0.147342
R14140 VSS.n825 VSS.n826 0.0732424
R14141 VSS.n826 VSS.n827 0.147342
R14142 VSS.n827 VSS.n2207 0.0732424
R14143 VSS.n2190 VSS.n2191 0.0722544
R14144 VSS.n2192 VSS.n2193 4.5005
R14145 VSS.n2194 VSS.n2195 4.5005
R14146 VSS.n2196 VSS.n2197 4.5005
R14147 VSS.n2192 VSS.n2190 2.37296
R14148 VSS.n2194 VSS.n2192 0.127318
R14149 VSS.n2196 VSS.n2194 0.127318
R14150 VSS.t20 VSS.n2196 2.73618
R14151 VSS.n2191 VSS.n758 4.5005
R14152 VSS.n2193 VSS.n760 4.5005
R14153 VSS.n2195 VSS.n761 4.5005
R14154 VSS.n2190 VSS.n756 4.57426
R14155 VSS.n2191 VSS.n2193 0.147342
R14156 VSS.n2193 VSS.n2195 0.147342
R14157 VSS.n2195 VSS.n2197 0.147342
R14158 VSS.n756 VSS.n758 0.147342
R14159 VSS.n759 VSS.n760 0.0732424
R14160 VSS.n760 VSS.n761 0.147342
R14161 VSS.n761 VSS.n2198 0.0732424
R14162 VSS.n2181 VSS.n2182 0.0722544
R14163 VSS.n2183 VSS.n2184 4.5005
R14164 VSS.n2185 VSS.n2186 4.5005
R14165 VSS.n2187 VSS.n2188 4.5005
R14166 VSS.n2183 VSS.n2181 2.37296
R14167 VSS.n2185 VSS.n2183 0.127318
R14168 VSS.n2187 VSS.n2185 0.127318
R14169 VSS.t20 VSS.n2187 2.73618
R14170 VSS.n2182 VSS.n707 4.5005
R14171 VSS.n2184 VSS.n709 4.5005
R14172 VSS.n2186 VSS.n710 4.5005
R14173 VSS.n2181 VSS.n705 4.57426
R14174 VSS.n2182 VSS.n2184 0.147342
R14175 VSS.n2184 VSS.n2186 0.147342
R14176 VSS.n2186 VSS.n2188 0.147342
R14177 VSS.n705 VSS.n707 0.147342
R14178 VSS.n708 VSS.n709 0.0732424
R14179 VSS.n709 VSS.n710 0.147342
R14180 VSS.n710 VSS.n2189 0.0732424
R14181 VSS.n2172 VSS.n2173 0.0722544
R14182 VSS.n2174 VSS.n2175 4.5005
R14183 VSS.n2176 VSS.n2177 4.5005
R14184 VSS.n2178 VSS.n2179 4.5005
R14185 VSS.n2174 VSS.n2172 2.37296
R14186 VSS.n2176 VSS.n2174 0.127318
R14187 VSS.n2178 VSS.n2176 0.127318
R14188 VSS.t20 VSS.n2178 2.73618
R14189 VSS.n2173 VSS.n611 4.5005
R14190 VSS.n2175 VSS.n613 4.5005
R14191 VSS.n2177 VSS.n614 4.5005
R14192 VSS.n2172 VSS.n609 4.57426
R14193 VSS.n2173 VSS.n2175 0.147342
R14194 VSS.n2175 VSS.n2177 0.147342
R14195 VSS.n2177 VSS.n2179 0.147342
R14196 VSS.n609 VSS.n611 0.147342
R14197 VSS.n612 VSS.n613 0.0732424
R14198 VSS.n613 VSS.n614 0.147342
R14199 VSS.n614 VSS.n2180 0.0732424
R14200 VSS.n2163 VSS.n2164 0.0722544
R14201 VSS.n2165 VSS.n2166 4.5005
R14202 VSS.n2167 VSS.n2168 4.5005
R14203 VSS.n2169 VSS.n2170 4.5005
R14204 VSS.n2165 VSS.n2163 2.37296
R14205 VSS.n2167 VSS.n2165 0.127318
R14206 VSS.n2169 VSS.n2167 0.127318
R14207 VSS.t20 VSS.n2169 2.73618
R14208 VSS.n2164 VSS.n560 4.5005
R14209 VSS.n2166 VSS.n562 4.5005
R14210 VSS.n2168 VSS.n563 4.5005
R14211 VSS.n2163 VSS.n558 4.57426
R14212 VSS.n2164 VSS.n2166 0.147342
R14213 VSS.n2166 VSS.n2168 0.147342
R14214 VSS.n2168 VSS.n2170 0.147342
R14215 VSS.n558 VSS.n560 0.147342
R14216 VSS.n561 VSS.n562 0.0732424
R14217 VSS.n562 VSS.n563 0.147342
R14218 VSS.n563 VSS.n2171 0.0732424
R14219 VSS.n2154 VSS.n2155 0.0722544
R14220 VSS.n2156 VSS.n2157 4.5005
R14221 VSS.n2158 VSS.n2159 4.5005
R14222 VSS.n2160 VSS.n2161 4.5005
R14223 VSS.n2156 VSS.n2154 2.37296
R14224 VSS.n2158 VSS.n2156 0.127318
R14225 VSS.n2160 VSS.n2158 0.127318
R14226 VSS.t20 VSS.n2160 2.73618
R14227 VSS.n2155 VSS.n494 4.5005
R14228 VSS.n2157 VSS.n496 4.5005
R14229 VSS.n2159 VSS.n497 4.5005
R14230 VSS.n2154 VSS.n492 4.57426
R14231 VSS.n2155 VSS.n2157 0.147342
R14232 VSS.n2157 VSS.n2159 0.147342
R14233 VSS.n2159 VSS.n2161 0.147342
R14234 VSS.n492 VSS.n494 0.147342
R14235 VSS.n495 VSS.n496 0.0732424
R14236 VSS.n496 VSS.n497 0.147342
R14237 VSS.n497 VSS.n2162 0.0732424
R14238 VSS.n2145 VSS.n2146 0.0722544
R14239 VSS.n2147 VSS.n2148 4.5005
R14240 VSS.n2149 VSS.n2150 4.5005
R14241 VSS.n2151 VSS.n2152 4.5005
R14242 VSS.n2147 VSS.n2145 2.37296
R14243 VSS.n2149 VSS.n2147 0.127318
R14244 VSS.n2151 VSS.n2149 0.127318
R14245 VSS.t20 VSS.n2151 2.73618
R14246 VSS.n2146 VSS.n443 4.5005
R14247 VSS.n2148 VSS.n445 4.5005
R14248 VSS.n2150 VSS.n446 4.5005
R14249 VSS.n2145 VSS.n441 4.57426
R14250 VSS.n2146 VSS.n2148 0.147342
R14251 VSS.n2148 VSS.n2150 0.147342
R14252 VSS.n2150 VSS.n2152 0.147342
R14253 VSS.n441 VSS.n443 0.147342
R14254 VSS.n444 VSS.n445 0.0732424
R14255 VSS.n445 VSS.n446 0.147342
R14256 VSS.n446 VSS.n2153 0.0732424
R14257 VSS.n2136 VSS.n2137 0.0722544
R14258 VSS.n2138 VSS.n2139 4.5005
R14259 VSS.n2140 VSS.n2141 4.5005
R14260 VSS.n2142 VSS.n2143 4.5005
R14261 VSS.n2138 VSS.n2136 2.37296
R14262 VSS.n2140 VSS.n2138 0.127318
R14263 VSS.n2142 VSS.n2140 0.127318
R14264 VSS.t20 VSS.n2142 2.73618
R14265 VSS.n2137 VSS.n347 4.5005
R14266 VSS.n2139 VSS.n349 4.5005
R14267 VSS.n2141 VSS.n350 4.5005
R14268 VSS.n2136 VSS.n345 4.57426
R14269 VSS.n2137 VSS.n2139 0.147342
R14270 VSS.n2139 VSS.n2141 0.147342
R14271 VSS.n2141 VSS.n2143 0.147342
R14272 VSS.n345 VSS.n347 0.147342
R14273 VSS.n348 VSS.n349 0.0732424
R14274 VSS.n349 VSS.n350 0.147342
R14275 VSS.n350 VSS.n2144 0.0732424
R14276 VSS.n2127 VSS.n2128 0.0722544
R14277 VSS.n2129 VSS.n2130 4.5005
R14278 VSS.n2131 VSS.n2132 4.5005
R14279 VSS.n2133 VSS.n2134 4.5005
R14280 VSS.n2129 VSS.n2127 2.37296
R14281 VSS.n2131 VSS.n2129 0.127318
R14282 VSS.n2133 VSS.n2131 0.127318
R14283 VSS.t20 VSS.n2133 2.73618
R14284 VSS.n2128 VSS.n296 4.5005
R14285 VSS.n2130 VSS.n298 4.5005
R14286 VSS.n2132 VSS.n299 4.5005
R14287 VSS.n2127 VSS.n294 4.57426
R14288 VSS.n2128 VSS.n2130 0.147342
R14289 VSS.n2130 VSS.n2132 0.147342
R14290 VSS.n2132 VSS.n2134 0.147342
R14291 VSS.n294 VSS.n296 0.147342
R14292 VSS.n297 VSS.n298 0.0732424
R14293 VSS.n298 VSS.n299 0.147342
R14294 VSS.n299 VSS.n2135 0.0732424
R14295 VSS.n2118 VSS.n2119 0.0722544
R14296 VSS.n2120 VSS.n2121 4.5005
R14297 VSS.n2122 VSS.n2123 4.5005
R14298 VSS.n2124 VSS.n2125 4.5005
R14299 VSS.n2120 VSS.n2118 2.37296
R14300 VSS.n2122 VSS.n2120 0.127318
R14301 VSS.n2124 VSS.n2122 0.127318
R14302 VSS.t20 VSS.n2124 2.73618
R14303 VSS.n2119 VSS.n230 4.5005
R14304 VSS.n2121 VSS.n232 4.5005
R14305 VSS.n2123 VSS.n233 4.5005
R14306 VSS.n2118 VSS.n228 4.57426
R14307 VSS.n2119 VSS.n2121 0.147342
R14308 VSS.n2121 VSS.n2123 0.147342
R14309 VSS.n2123 VSS.n2125 0.147342
R14310 VSS.n228 VSS.n230 0.147342
R14311 VSS.n231 VSS.n232 0.0732424
R14312 VSS.n232 VSS.n233 0.147342
R14313 VSS.n233 VSS.n2126 0.0732424
R14314 VSS.n2109 VSS.n2110 0.0722544
R14315 VSS.n2111 VSS.n2112 4.5005
R14316 VSS.n2113 VSS.n2114 4.5005
R14317 VSS.n2115 VSS.n2116 4.5005
R14318 VSS.n2111 VSS.n2109 2.37296
R14319 VSS.n2113 VSS.n2111 0.127318
R14320 VSS.n2115 VSS.n2113 0.127318
R14321 VSS.t20 VSS.n2115 2.73618
R14322 VSS.n2110 VSS.n179 4.5005
R14323 VSS.n2112 VSS.n181 4.5005
R14324 VSS.n2114 VSS.n182 4.5005
R14325 VSS.n2109 VSS.n177 4.57426
R14326 VSS.n2110 VSS.n2112 0.147342
R14327 VSS.n2112 VSS.n2114 0.147342
R14328 VSS.n2114 VSS.n2116 0.147342
R14329 VSS.n177 VSS.n179 0.147342
R14330 VSS.n180 VSS.n181 0.0732424
R14331 VSS.n181 VSS.n182 0.147342
R14332 VSS.n182 VSS.n2117 0.0732424
R14333 VSS.n2099 VSS.n2100 0.0722544
R14334 VSS.n2101 VSS.n2102 4.5005
R14335 VSS.n2103 VSS.n2104 4.5005
R14336 VSS.n2105 VSS.n2106 4.5005
R14337 VSS.n2101 VSS.n2099 2.37296
R14338 VSS.n2103 VSS.n2101 0.127318
R14339 VSS.n2105 VSS.n2103 0.127318
R14340 VSS.t20 VSS.n2105 2.73618
R14341 VSS.n2100 VSS.n83 4.5005
R14342 VSS.n2102 VSS.n85 4.5005
R14343 VSS.n2104 VSS.n86 4.5005
R14344 VSS.n2099 VSS.n81 4.57426
R14345 VSS.n2100 VSS.n2102 0.147342
R14346 VSS.n2102 VSS.n2104 0.147342
R14347 VSS.n2104 VSS.n2106 0.147342
R14348 VSS.n81 VSS.n83 0.147342
R14349 VSS.n84 VSS.n85 0.0732424
R14350 VSS.n85 VSS.n86 0.147342
R14351 VSS.n86 VSS.n2107 0.0732424
R14352 VSS.n2090 VSS.n2091 0.0722544
R14353 VSS.n2092 VSS.n2093 4.5005
R14354 VSS.n2094 VSS.n2095 4.5005
R14355 VSS.n2096 VSS.n2097 4.5005
R14356 VSS.n2092 VSS.n2090 2.37296
R14357 VSS.n2094 VSS.n2092 0.127318
R14358 VSS.n2096 VSS.n2094 0.127318
R14359 VSS.t20 VSS.n2096 2.73618
R14360 VSS.n2091 VSS.n32 4.5005
R14361 VSS.n2093 VSS.n34 4.5005
R14362 VSS.n2095 VSS.n35 4.5005
R14363 VSS.n2090 VSS.n30 4.57426
R14364 VSS.n2091 VSS.n2093 0.147342
R14365 VSS.n2093 VSS.n2095 0.147342
R14366 VSS.n2095 VSS.n2097 0.147342
R14367 VSS.n30 VSS.n32 0.147342
R14368 VSS.n33 VSS.n34 0.0732424
R14369 VSS.n34 VSS.n35 0.147342
R14370 VSS.n35 VSS.n2098 0.0732424
R14371 VSS.n2063 VSS.n2068 4.5005
R14372 VSS.n2065 VSS.n2069 4.5005
R14373 VSS.n2066 VSS.n2070 4.5005
R14374 VSS.n2067 VSS.n2071 4.57324
R14375 VSS.n2063 VSS.n2061 0.147342
R14376 VSS.n2064 VSS.n2065 0.0732424
R14377 VSS.n2065 VSS.n2066 0.147342
R14378 VSS.n2068 VSS.n2072 0.0721009
R14379 VSS.n2073 VSS.n2069 4.5005
R14380 VSS.n2074 VSS.n2070 4.5005
R14381 VSS.n2075 VSS.n2071 4.5005
R14382 VSS.n2061 VSS.n2072 4.57442
R14383 VSS.n2068 VSS.n2069 0.147342
R14384 VSS.n2069 VSS.n2070 0.147342
R14385 VSS.n2070 VSS.n2071 0.147342
R14386 VSS.n2072 VSS.n2073 2.39784
R14387 VSS.n2073 VSS.n2074 0.147342
R14388 VSS.n2074 VSS.n2075 0.147342
R14389 VSS.n2075 VSS.t561 3.13212
R14390 VSS.n2048 VSS.n2053 4.5005
R14391 VSS.n2050 VSS.n2054 4.5005
R14392 VSS.n2051 VSS.n2055 4.5005
R14393 VSS.n2052 VSS.n2056 4.57324
R14394 VSS.n2048 VSS.n2046 0.147342
R14395 VSS.n2049 VSS.n2050 0.0732424
R14396 VSS.n2050 VSS.n2051 0.147342
R14397 VSS.n2053 VSS.n2057 0.0721009
R14398 VSS.n2058 VSS.n2054 4.5005
R14399 VSS.n2059 VSS.n2055 4.5005
R14400 VSS.n2060 VSS.n2056 4.5005
R14401 VSS.n2046 VSS.n2057 4.57442
R14402 VSS.n2053 VSS.n2054 0.147342
R14403 VSS.n2054 VSS.n2055 0.147342
R14404 VSS.n2055 VSS.n2056 0.147342
R14405 VSS.n2057 VSS.n2058 2.39784
R14406 VSS.n2058 VSS.n2059 0.147342
R14407 VSS.n2059 VSS.n2060 0.147342
R14408 VSS.n2060 VSS.t377 3.13212
R14409 VSS.n2033 VSS.n2038 4.5005
R14410 VSS.n2035 VSS.n2039 4.5005
R14411 VSS.n2036 VSS.n2040 4.5005
R14412 VSS.n2037 VSS.n2041 4.57324
R14413 VSS.n2033 VSS.n2031 0.147342
R14414 VSS.n2034 VSS.n2035 0.0732424
R14415 VSS.n2035 VSS.n2036 0.147342
R14416 VSS.n2038 VSS.n2042 0.0721009
R14417 VSS.n2043 VSS.n2039 4.5005
R14418 VSS.n2044 VSS.n2040 4.5005
R14419 VSS.n2045 VSS.n2041 4.5005
R14420 VSS.n2031 VSS.n2042 4.57442
R14421 VSS.n2038 VSS.n2039 0.147342
R14422 VSS.n2039 VSS.n2040 0.147342
R14423 VSS.n2040 VSS.n2041 0.147342
R14424 VSS.n2042 VSS.n2043 2.39784
R14425 VSS.n2043 VSS.n2044 0.147342
R14426 VSS.n2044 VSS.n2045 0.147342
R14427 VSS.n2045 VSS.t596 3.13212
R14428 VSS.n2012 VSS.n2017 4.5005
R14429 VSS.n2014 VSS.n2018 4.5005
R14430 VSS.n2015 VSS.n2019 4.5005
R14431 VSS.n2016 VSS.n2020 4.57324
R14432 VSS.n2012 VSS.n2010 0.147342
R14433 VSS.n2013 VSS.n2014 0.0732424
R14434 VSS.n2014 VSS.n2015 0.147342
R14435 VSS.n2017 VSS.n2021 0.0721009
R14436 VSS.n2022 VSS.n2018 4.5005
R14437 VSS.n2023 VSS.n2019 4.5005
R14438 VSS.n2024 VSS.n2020 4.5005
R14439 VSS.n2010 VSS.n2021 4.57442
R14440 VSS.n2017 VSS.n2018 0.147342
R14441 VSS.n2018 VSS.n2019 0.147342
R14442 VSS.n2019 VSS.n2020 0.147342
R14443 VSS.n2021 VSS.n2022 2.39784
R14444 VSS.n2022 VSS.n2023 0.147342
R14445 VSS.n2023 VSS.n2024 0.147342
R14446 VSS.n2024 VSS.t368 3.13212
R14447 VSS.n1997 VSS.n2002 4.5005
R14448 VSS.n1999 VSS.n2003 4.5005
R14449 VSS.n2000 VSS.n2004 4.5005
R14450 VSS.n2001 VSS.n2005 4.57324
R14451 VSS.n1997 VSS.n1995 0.147342
R14452 VSS.n1998 VSS.n1999 0.0732424
R14453 VSS.n1999 VSS.n2000 0.147342
R14454 VSS.n2002 VSS.n2006 0.0721009
R14455 VSS.n2007 VSS.n2003 4.5005
R14456 VSS.n2008 VSS.n2004 4.5005
R14457 VSS.n2009 VSS.n2005 4.5005
R14458 VSS.n1995 VSS.n2006 4.57442
R14459 VSS.n2002 VSS.n2003 0.147342
R14460 VSS.n2003 VSS.n2004 0.147342
R14461 VSS.n2004 VSS.n2005 0.147342
R14462 VSS.n2006 VSS.n2007 2.39784
R14463 VSS.n2007 VSS.n2008 0.147342
R14464 VSS.n2008 VSS.n2009 0.147342
R14465 VSS.n2009 VSS.t344 3.13212
R14466 VSS.n1982 VSS.n1987 4.5005
R14467 VSS.n1984 VSS.n1988 4.5005
R14468 VSS.n1985 VSS.n1989 4.5005
R14469 VSS.n1986 VSS.n1990 4.57324
R14470 VSS.n1982 VSS.n1980 0.147342
R14471 VSS.n1983 VSS.n1984 0.0732424
R14472 VSS.n1984 VSS.n1985 0.147342
R14473 VSS.n1987 VSS.n1991 0.0721009
R14474 VSS.n1992 VSS.n1988 4.5005
R14475 VSS.n1993 VSS.n1989 4.5005
R14476 VSS.n1994 VSS.n1990 4.5005
R14477 VSS.n1980 VSS.n1991 4.57442
R14478 VSS.n1987 VSS.n1988 0.147342
R14479 VSS.n1988 VSS.n1989 0.147342
R14480 VSS.n1989 VSS.n1990 0.147342
R14481 VSS.n1991 VSS.n1992 2.39784
R14482 VSS.n1992 VSS.n1993 0.147342
R14483 VSS.n1993 VSS.n1994 0.147342
R14484 VSS.n1994 VSS.t426 3.13212
R14485 VSS.n1967 VSS.n1972 4.5005
R14486 VSS.n1969 VSS.n1973 4.5005
R14487 VSS.n1970 VSS.n1974 4.5005
R14488 VSS.n1971 VSS.n1975 4.57324
R14489 VSS.n1967 VSS.n1965 0.147342
R14490 VSS.n1968 VSS.n1969 0.0732424
R14491 VSS.n1969 VSS.n1970 0.147342
R14492 VSS.n1972 VSS.n1976 0.0721009
R14493 VSS.n1977 VSS.n1973 4.5005
R14494 VSS.n1978 VSS.n1974 4.5005
R14495 VSS.n1979 VSS.n1975 4.5005
R14496 VSS.n1965 VSS.n1976 4.57442
R14497 VSS.n1972 VSS.n1973 0.147342
R14498 VSS.n1973 VSS.n1974 0.147342
R14499 VSS.n1974 VSS.n1975 0.147342
R14500 VSS.n1976 VSS.n1977 2.39784
R14501 VSS.n1977 VSS.n1978 0.147342
R14502 VSS.n1978 VSS.n1979 0.147342
R14503 VSS.n1979 VSS.t81 3.13212
R14504 VSS.n1952 VSS.n1957 4.5005
R14505 VSS.n1954 VSS.n1958 4.5005
R14506 VSS.n1955 VSS.n1959 4.5005
R14507 VSS.n1956 VSS.n1960 4.57324
R14508 VSS.n1952 VSS.n1950 0.147342
R14509 VSS.n1953 VSS.n1954 0.0732424
R14510 VSS.n1954 VSS.n1955 0.147342
R14511 VSS.n1957 VSS.n1961 0.0721009
R14512 VSS.n1962 VSS.n1958 4.5005
R14513 VSS.n1963 VSS.n1959 4.5005
R14514 VSS.n1964 VSS.n1960 4.5005
R14515 VSS.n1950 VSS.n1961 4.57442
R14516 VSS.n1957 VSS.n1958 0.147342
R14517 VSS.n1958 VSS.n1959 0.147342
R14518 VSS.n1959 VSS.n1960 0.147342
R14519 VSS.n1961 VSS.n1962 2.39784
R14520 VSS.n1962 VSS.n1963 0.147342
R14521 VSS.n1963 VSS.n1964 0.147342
R14522 VSS.n1964 VSS.t24 3.13212
R14523 VSS.n1937 VSS.n1942 4.5005
R14524 VSS.n1939 VSS.n1943 4.5005
R14525 VSS.n1940 VSS.n1944 4.5005
R14526 VSS.n1941 VSS.n1945 4.57324
R14527 VSS.n1937 VSS.n1935 0.147342
R14528 VSS.n1938 VSS.n1939 0.0732424
R14529 VSS.n1939 VSS.n1940 0.147342
R14530 VSS.n1942 VSS.n1946 0.0721009
R14531 VSS.n1947 VSS.n1943 4.5005
R14532 VSS.n1948 VSS.n1944 4.5005
R14533 VSS.n1949 VSS.n1945 4.5005
R14534 VSS.n1935 VSS.n1946 4.57442
R14535 VSS.n1942 VSS.n1943 0.147342
R14536 VSS.n1943 VSS.n1944 0.147342
R14537 VSS.n1944 VSS.n1945 0.147342
R14538 VSS.n1946 VSS.n1947 2.39784
R14539 VSS.n1947 VSS.n1948 0.147342
R14540 VSS.n1948 VSS.n1949 0.147342
R14541 VSS.n1949 VSS.t396 3.13212
R14542 VSS.n1916 VSS.n1921 4.5005
R14543 VSS.n1918 VSS.n1922 4.5005
R14544 VSS.n1919 VSS.n1923 4.5005
R14545 VSS.n1920 VSS.n1924 4.57324
R14546 VSS.n1916 VSS.n1914 0.147342
R14547 VSS.n1917 VSS.n1918 0.0732424
R14548 VSS.n1918 VSS.n1919 0.147342
R14549 VSS.n1921 VSS.n1925 0.0721009
R14550 VSS.n1926 VSS.n1922 4.5005
R14551 VSS.n1927 VSS.n1923 4.5005
R14552 VSS.n1928 VSS.n1924 4.5005
R14553 VSS.n1914 VSS.n1925 4.57442
R14554 VSS.n1921 VSS.n1922 0.147342
R14555 VSS.n1922 VSS.n1923 0.147342
R14556 VSS.n1923 VSS.n1924 0.147342
R14557 VSS.n1925 VSS.n1926 2.39784
R14558 VSS.n1926 VSS.n1927 0.147342
R14559 VSS.n1927 VSS.n1928 0.147342
R14560 VSS.n1928 VSS.t316 3.13212
R14561 VSS.n1901 VSS.n1906 4.5005
R14562 VSS.n1903 VSS.n1907 4.5005
R14563 VSS.n1904 VSS.n1908 4.5005
R14564 VSS.n1905 VSS.n1909 4.57324
R14565 VSS.n1901 VSS.n1899 0.147342
R14566 VSS.n1902 VSS.n1903 0.0732424
R14567 VSS.n1903 VSS.n1904 0.147342
R14568 VSS.n1906 VSS.n1910 0.0721009
R14569 VSS.n1911 VSS.n1907 4.5005
R14570 VSS.n1912 VSS.n1908 4.5005
R14571 VSS.n1913 VSS.n1909 4.5005
R14572 VSS.n1899 VSS.n1910 4.57442
R14573 VSS.n1906 VSS.n1907 0.147342
R14574 VSS.n1907 VSS.n1908 0.147342
R14575 VSS.n1908 VSS.n1909 0.147342
R14576 VSS.n1910 VSS.n1911 2.39784
R14577 VSS.n1911 VSS.n1912 0.147342
R14578 VSS.n1912 VSS.n1913 0.147342
R14579 VSS.n1913 VSS.t335 3.13212
R14580 VSS.n1886 VSS.n1891 4.5005
R14581 VSS.n1888 VSS.n1892 4.5005
R14582 VSS.n1889 VSS.n1893 4.5005
R14583 VSS.n1890 VSS.n1894 4.57324
R14584 VSS.n1886 VSS.n1884 0.147342
R14585 VSS.n1887 VSS.n1888 0.0732424
R14586 VSS.n1888 VSS.n1889 0.147342
R14587 VSS.n1891 VSS.n1895 0.0721009
R14588 VSS.n1896 VSS.n1892 4.5005
R14589 VSS.n1897 VSS.n1893 4.5005
R14590 VSS.n1898 VSS.n1894 4.5005
R14591 VSS.n1884 VSS.n1895 4.57442
R14592 VSS.n1891 VSS.n1892 0.147342
R14593 VSS.n1892 VSS.n1893 0.147342
R14594 VSS.n1893 VSS.n1894 0.147342
R14595 VSS.n1895 VSS.n1896 2.39784
R14596 VSS.n1896 VSS.n1897 0.147342
R14597 VSS.n1897 VSS.n1898 0.147342
R14598 VSS.n1898 VSS.t393 3.13212
R14599 VSS.n1865 VSS.n1870 4.5005
R14600 VSS.n1867 VSS.n1871 4.5005
R14601 VSS.n1868 VSS.n1872 4.5005
R14602 VSS.n1869 VSS.n1873 4.57324
R14603 VSS.n1865 VSS.n1863 0.147342
R14604 VSS.n1866 VSS.n1867 0.0732424
R14605 VSS.n1867 VSS.n1868 0.147342
R14606 VSS.n1870 VSS.n1874 0.0721009
R14607 VSS.n1875 VSS.n1871 4.5005
R14608 VSS.n1876 VSS.n1872 4.5005
R14609 VSS.n1877 VSS.n1873 4.5005
R14610 VSS.n1863 VSS.n1874 4.57442
R14611 VSS.n1870 VSS.n1871 0.147342
R14612 VSS.n1871 VSS.n1872 0.147342
R14613 VSS.n1872 VSS.n1873 0.147342
R14614 VSS.n1874 VSS.n1875 2.39784
R14615 VSS.n1875 VSS.n1876 0.147342
R14616 VSS.n1876 VSS.n1877 0.147342
R14617 VSS.n1877 VSS.t381 3.13212
R14618 VSS.n1850 VSS.n1855 4.5005
R14619 VSS.n1852 VSS.n1856 4.5005
R14620 VSS.n1853 VSS.n1857 4.5005
R14621 VSS.n1854 VSS.n1858 4.57324
R14622 VSS.n1850 VSS.n1848 0.147342
R14623 VSS.n1851 VSS.n1852 0.0732424
R14624 VSS.n1852 VSS.n1853 0.147342
R14625 VSS.n1855 VSS.n1859 0.0721009
R14626 VSS.n1860 VSS.n1856 4.5005
R14627 VSS.n1861 VSS.n1857 4.5005
R14628 VSS.n1862 VSS.n1858 4.5005
R14629 VSS.n1848 VSS.n1859 4.57442
R14630 VSS.n1855 VSS.n1856 0.147342
R14631 VSS.n1856 VSS.n1857 0.147342
R14632 VSS.n1857 VSS.n1858 0.147342
R14633 VSS.n1859 VSS.n1860 2.39784
R14634 VSS.n1860 VSS.n1861 0.147342
R14635 VSS.n1861 VSS.n1862 0.147342
R14636 VSS.n1862 VSS.t174 3.13212
R14637 VSS.n1835 VSS.n1840 4.5005
R14638 VSS.n1837 VSS.n1841 4.5005
R14639 VSS.n1838 VSS.n1842 4.5005
R14640 VSS.n1839 VSS.n1843 4.57324
R14641 VSS.n1835 VSS.n1833 0.147342
R14642 VSS.n1836 VSS.n1837 0.0732424
R14643 VSS.n1837 VSS.n1838 0.147342
R14644 VSS.n1840 VSS.n1844 0.0721009
R14645 VSS.n1845 VSS.n1841 4.5005
R14646 VSS.n1846 VSS.n1842 4.5005
R14647 VSS.n1847 VSS.n1843 4.5005
R14648 VSS.n1833 VSS.n1844 4.57442
R14649 VSS.n1840 VSS.n1841 0.147342
R14650 VSS.n1841 VSS.n1842 0.147342
R14651 VSS.n1842 VSS.n1843 0.147342
R14652 VSS.n1844 VSS.n1845 2.39784
R14653 VSS.n1845 VSS.n1846 0.147342
R14654 VSS.n1846 VSS.n1847 0.147342
R14655 VSS.n1847 VSS.t225 3.13212
R14656 VSS.n1820 VSS.n1825 4.5005
R14657 VSS.n1822 VSS.n1826 4.5005
R14658 VSS.n1823 VSS.n1827 4.5005
R14659 VSS.n1824 VSS.n1828 4.57324
R14660 VSS.n1820 VSS.n1818 0.147342
R14661 VSS.n1821 VSS.n1822 0.0732424
R14662 VSS.n1822 VSS.n1823 0.147342
R14663 VSS.n1825 VSS.n1829 0.0721009
R14664 VSS.n1830 VSS.n1826 4.5005
R14665 VSS.n1831 VSS.n1827 4.5005
R14666 VSS.n1832 VSS.n1828 4.5005
R14667 VSS.n1818 VSS.n1829 4.57442
R14668 VSS.n1825 VSS.n1826 0.147342
R14669 VSS.n1826 VSS.n1827 0.147342
R14670 VSS.n1827 VSS.n1828 0.147342
R14671 VSS.n1829 VSS.n1830 2.39784
R14672 VSS.n1830 VSS.n1831 0.147342
R14673 VSS.n1831 VSS.n1832 0.147342
R14674 VSS.n1832 VSS.t304 3.13212
R14675 VSS.n1799 VSS.n1804 4.5005
R14676 VSS.n1801 VSS.n1805 4.5005
R14677 VSS.n1802 VSS.n1806 4.5005
R14678 VSS.n1803 VSS.n1807 4.57324
R14679 VSS.n1799 VSS.n1797 0.147342
R14680 VSS.n1800 VSS.n1801 0.0732424
R14681 VSS.n1801 VSS.n1802 0.147342
R14682 VSS.n1804 VSS.n1808 0.0721009
R14683 VSS.n1809 VSS.n1805 4.5005
R14684 VSS.n1810 VSS.n1806 4.5005
R14685 VSS.n1811 VSS.n1807 4.5005
R14686 VSS.n1797 VSS.n1808 4.57442
R14687 VSS.n1804 VSS.n1805 0.147342
R14688 VSS.n1805 VSS.n1806 0.147342
R14689 VSS.n1806 VSS.n1807 0.147342
R14690 VSS.n1808 VSS.n1809 2.39784
R14691 VSS.n1809 VSS.n1810 0.147342
R14692 VSS.n1810 VSS.n1811 0.147342
R14693 VSS.n1811 VSS.t434 3.13212
R14694 VSS.n1784 VSS.n1789 4.5005
R14695 VSS.n1786 VSS.n1790 4.5005
R14696 VSS.n1787 VSS.n1791 4.5005
R14697 VSS.n1788 VSS.n1792 4.57324
R14698 VSS.n1784 VSS.n1782 0.147342
R14699 VSS.n1785 VSS.n1786 0.0732424
R14700 VSS.n1786 VSS.n1787 0.147342
R14701 VSS.n1789 VSS.n1793 0.0721009
R14702 VSS.n1794 VSS.n1790 4.5005
R14703 VSS.n1795 VSS.n1791 4.5005
R14704 VSS.n1796 VSS.n1792 4.5005
R14705 VSS.n1782 VSS.n1793 4.57442
R14706 VSS.n1789 VSS.n1790 0.147342
R14707 VSS.n1790 VSS.n1791 0.147342
R14708 VSS.n1791 VSS.n1792 0.147342
R14709 VSS.n1793 VSS.n1794 2.39784
R14710 VSS.n1794 VSS.n1795 0.147342
R14711 VSS.n1795 VSS.n1796 0.147342
R14712 VSS.n1796 VSS.t373 3.13212
R14713 VSS.n1769 VSS.n1774 4.5005
R14714 VSS.n1771 VSS.n1775 4.5005
R14715 VSS.n1772 VSS.n1776 4.5005
R14716 VSS.n1773 VSS.n1777 4.57324
R14717 VSS.n1769 VSS.n1767 0.147342
R14718 VSS.n1770 VSS.n1771 0.0732424
R14719 VSS.n1771 VSS.n1772 0.147342
R14720 VSS.n1774 VSS.n1778 0.0721009
R14721 VSS.n1779 VSS.n1775 4.5005
R14722 VSS.n1780 VSS.n1776 4.5005
R14723 VSS.n1781 VSS.n1777 4.5005
R14724 VSS.n1767 VSS.n1778 4.57442
R14725 VSS.n1774 VSS.n1775 0.147342
R14726 VSS.n1775 VSS.n1776 0.147342
R14727 VSS.n1776 VSS.n1777 0.147342
R14728 VSS.n1778 VSS.n1779 2.39784
R14729 VSS.n1779 VSS.n1780 0.147342
R14730 VSS.n1780 VSS.n1781 0.147342
R14731 VSS.n1781 VSS.t594 3.13212
R14732 VSS.n1748 VSS.n1753 4.5005
R14733 VSS.n1750 VSS.n1754 4.5005
R14734 VSS.n1751 VSS.n1755 4.5005
R14735 VSS.n1752 VSS.n1756 4.57324
R14736 VSS.n1748 VSS.n1746 0.147342
R14737 VSS.n1749 VSS.n1750 0.0732424
R14738 VSS.n1750 VSS.n1751 0.147342
R14739 VSS.n1753 VSS.n1757 0.0721009
R14740 VSS.n1758 VSS.n1754 4.5005
R14741 VSS.n1759 VSS.n1755 4.5005
R14742 VSS.n1760 VSS.n1756 4.5005
R14743 VSS.n1746 VSS.n1757 4.57442
R14744 VSS.n1753 VSS.n1754 0.147342
R14745 VSS.n1754 VSS.n1755 0.147342
R14746 VSS.n1755 VSS.n1756 0.147342
R14747 VSS.n1757 VSS.n1758 2.39784
R14748 VSS.n1758 VSS.n1759 0.147342
R14749 VSS.n1759 VSS.n1760 0.147342
R14750 VSS.n1760 VSS.t371 3.13212
R14751 VSS.n1733 VSS.n1738 4.5005
R14752 VSS.n1735 VSS.n1739 4.5005
R14753 VSS.n1736 VSS.n1740 4.5005
R14754 VSS.n1737 VSS.n1741 4.57324
R14755 VSS.n1733 VSS.n1731 0.147342
R14756 VSS.n1734 VSS.n1735 0.0732424
R14757 VSS.n1735 VSS.n1736 0.147342
R14758 VSS.n1738 VSS.n1742 0.0721009
R14759 VSS.n1743 VSS.n1739 4.5005
R14760 VSS.n1744 VSS.n1740 4.5005
R14761 VSS.n1745 VSS.n1741 4.5005
R14762 VSS.n1731 VSS.n1742 4.57442
R14763 VSS.n1738 VSS.n1739 0.147342
R14764 VSS.n1739 VSS.n1740 0.147342
R14765 VSS.n1740 VSS.n1741 0.147342
R14766 VSS.n1742 VSS.n1743 2.39784
R14767 VSS.n1743 VSS.n1744 0.147342
R14768 VSS.n1744 VSS.n1745 0.147342
R14769 VSS.n1745 VSS.t581 3.13212
R14770 VSS.n1718 VSS.n1723 4.5005
R14771 VSS.n1720 VSS.n1724 4.5005
R14772 VSS.n1721 VSS.n1725 4.5005
R14773 VSS.n1722 VSS.n1726 4.57324
R14774 VSS.n1718 VSS.n1716 0.147342
R14775 VSS.n1719 VSS.n1720 0.0732424
R14776 VSS.n1720 VSS.n1721 0.147342
R14777 VSS.n1723 VSS.n1727 0.0721009
R14778 VSS.n1728 VSS.n1724 4.5005
R14779 VSS.n1729 VSS.n1725 4.5005
R14780 VSS.n1730 VSS.n1726 4.5005
R14781 VSS.n1716 VSS.n1727 4.57442
R14782 VSS.n1723 VSS.n1724 0.147342
R14783 VSS.n1724 VSS.n1725 0.147342
R14784 VSS.n1725 VSS.n1726 0.147342
R14785 VSS.n1727 VSS.n1728 2.39784
R14786 VSS.n1728 VSS.n1729 0.147342
R14787 VSS.n1729 VSS.n1730 0.147342
R14788 VSS.n1730 VSS.t272 3.13212
R14789 VSS.n1703 VSS.n1708 4.5005
R14790 VSS.n1705 VSS.n1709 4.5005
R14791 VSS.n1706 VSS.n1710 4.5005
R14792 VSS.n1707 VSS.n1711 4.57324
R14793 VSS.n1703 VSS.n1701 0.147342
R14794 VSS.n1704 VSS.n1705 0.0732424
R14795 VSS.n1705 VSS.n1706 0.147342
R14796 VSS.n1708 VSS.n1712 0.0721009
R14797 VSS.n1713 VSS.n1709 4.5005
R14798 VSS.n1714 VSS.n1710 4.5005
R14799 VSS.n1715 VSS.n1711 4.5005
R14800 VSS.n1701 VSS.n1712 4.57442
R14801 VSS.n1708 VSS.n1709 0.147342
R14802 VSS.n1709 VSS.n1710 0.147342
R14803 VSS.n1710 VSS.n1711 0.147342
R14804 VSS.n1712 VSS.n1713 2.39784
R14805 VSS.n1713 VSS.n1714 0.147342
R14806 VSS.n1714 VSS.n1715 0.147342
R14807 VSS.n1715 VSS.t503 3.13212
R14808 VSS.n1688 VSS.n1693 4.5005
R14809 VSS.n1690 VSS.n1694 4.5005
R14810 VSS.n1691 VSS.n1695 4.5005
R14811 VSS.n1692 VSS.n1696 4.57324
R14812 VSS.n1688 VSS.n1686 0.147342
R14813 VSS.n1689 VSS.n1690 0.0732424
R14814 VSS.n1690 VSS.n1691 0.147342
R14815 VSS.n1693 VSS.n1697 0.0721009
R14816 VSS.n1698 VSS.n1694 4.5005
R14817 VSS.n1699 VSS.n1695 4.5005
R14818 VSS.n1700 VSS.n1696 4.5005
R14819 VSS.n1686 VSS.n1697 4.57442
R14820 VSS.n1693 VSS.n1694 0.147342
R14821 VSS.n1694 VSS.n1695 0.147342
R14822 VSS.n1695 VSS.n1696 0.147342
R14823 VSS.n1697 VSS.n1698 2.39784
R14824 VSS.n1698 VSS.n1699 0.147342
R14825 VSS.n1699 VSS.n1700 0.147342
R14826 VSS.n1700 VSS.t26 3.13212
R14827 VSS.n1673 VSS.n1678 4.5005
R14828 VSS.n1675 VSS.n1679 4.5005
R14829 VSS.n1676 VSS.n1680 4.5005
R14830 VSS.n1677 VSS.n1681 4.57324
R14831 VSS.n1673 VSS.n1671 0.147342
R14832 VSS.n1674 VSS.n1675 0.0732424
R14833 VSS.n1675 VSS.n1676 0.147342
R14834 VSS.n1678 VSS.n1682 0.0721009
R14835 VSS.n1683 VSS.n1679 4.5005
R14836 VSS.n1684 VSS.n1680 4.5005
R14837 VSS.n1685 VSS.n1681 4.5005
R14838 VSS.n1671 VSS.n1682 4.57442
R14839 VSS.n1678 VSS.n1679 0.147342
R14840 VSS.n1679 VSS.n1680 0.147342
R14841 VSS.n1680 VSS.n1681 0.147342
R14842 VSS.n1682 VSS.n1683 2.39784
R14843 VSS.n1683 VSS.n1684 0.147342
R14844 VSS.n1684 VSS.n1685 0.147342
R14845 VSS.n1685 VSS.t355 3.13212
R14846 VSS.n1652 VSS.n1657 4.5005
R14847 VSS.n1654 VSS.n1658 4.5005
R14848 VSS.n1655 VSS.n1659 4.5005
R14849 VSS.n1656 VSS.n1660 4.57324
R14850 VSS.n1652 VSS.n1650 0.147342
R14851 VSS.n1653 VSS.n1654 0.0732424
R14852 VSS.n1654 VSS.n1655 0.147342
R14853 VSS.n1657 VSS.n1661 0.0721009
R14854 VSS.n1662 VSS.n1658 4.5005
R14855 VSS.n1663 VSS.n1659 4.5005
R14856 VSS.n1664 VSS.n1660 4.5005
R14857 VSS.n1650 VSS.n1661 4.57442
R14858 VSS.n1657 VSS.n1658 0.147342
R14859 VSS.n1658 VSS.n1659 0.147342
R14860 VSS.n1659 VSS.n1660 0.147342
R14861 VSS.n1661 VSS.n1662 2.39784
R14862 VSS.n1662 VSS.n1663 0.147342
R14863 VSS.n1663 VSS.n1664 0.147342
R14864 VSS.n1664 VSS.t358 3.13212
R14865 VSS.n1637 VSS.n1642 4.5005
R14866 VSS.n1639 VSS.n1643 4.5005
R14867 VSS.n1640 VSS.n1644 4.5005
R14868 VSS.n1641 VSS.n1645 4.57324
R14869 VSS.n1637 VSS.n1635 0.147342
R14870 VSS.n1638 VSS.n1639 0.0732424
R14871 VSS.n1639 VSS.n1640 0.147342
R14872 VSS.n1642 VSS.n1646 0.0721009
R14873 VSS.n1647 VSS.n1643 4.5005
R14874 VSS.n1648 VSS.n1644 4.5005
R14875 VSS.n1649 VSS.n1645 4.5005
R14876 VSS.n1635 VSS.n1646 4.57442
R14877 VSS.n1642 VSS.n1643 0.147342
R14878 VSS.n1643 VSS.n1644 0.147342
R14879 VSS.n1644 VSS.n1645 0.147342
R14880 VSS.n1646 VSS.n1647 2.39784
R14881 VSS.n1647 VSS.n1648 0.147342
R14882 VSS.n1648 VSS.n1649 0.147342
R14883 VSS.n1649 VSS.t338 3.13212
R14884 VSS.n1622 VSS.n1627 4.5005
R14885 VSS.n1624 VSS.n1628 4.5005
R14886 VSS.n1625 VSS.n1629 4.5005
R14887 VSS.n1626 VSS.n1630 4.57324
R14888 VSS.n1622 VSS.n1620 0.147342
R14889 VSS.n1623 VSS.n1624 0.0732424
R14890 VSS.n1624 VSS.n1625 0.147342
R14891 VSS.n1627 VSS.n1631 0.0721009
R14892 VSS.n1632 VSS.n1628 4.5005
R14893 VSS.n1633 VSS.n1629 4.5005
R14894 VSS.n1634 VSS.n1630 4.5005
R14895 VSS.n1620 VSS.n1631 4.57442
R14896 VSS.n1627 VSS.n1628 0.147342
R14897 VSS.n1628 VSS.n1629 0.147342
R14898 VSS.n1629 VSS.n1630 0.147342
R14899 VSS.n1631 VSS.n1632 2.39784
R14900 VSS.n1632 VSS.n1633 0.147342
R14901 VSS.n1633 VSS.n1634 0.147342
R14902 VSS.n1634 VSS.t321 3.13212
R14903 VSS.n1601 VSS.n1606 4.5005
R14904 VSS.n1603 VSS.n1607 4.5005
R14905 VSS.n1604 VSS.n1608 4.5005
R14906 VSS.n1605 VSS.n1609 4.57324
R14907 VSS.n1601 VSS.n1599 0.147342
R14908 VSS.n1602 VSS.n1603 0.0732424
R14909 VSS.n1603 VSS.n1604 0.147342
R14910 VSS.n1606 VSS.n1610 0.0721009
R14911 VSS.n1611 VSS.n1607 4.5005
R14912 VSS.n1612 VSS.n1608 4.5005
R14913 VSS.n1613 VSS.n1609 4.5005
R14914 VSS.n1599 VSS.n1610 4.57442
R14915 VSS.n1606 VSS.n1607 0.147342
R14916 VSS.n1607 VSS.n1608 0.147342
R14917 VSS.n1608 VSS.n1609 0.147342
R14918 VSS.n1610 VSS.n1611 2.39784
R14919 VSS.n1611 VSS.n1612 0.147342
R14920 VSS.n1612 VSS.n1613 0.147342
R14921 VSS.n1613 VSS.t387 3.13212
R14922 VSS.n1586 VSS.n1591 4.5005
R14923 VSS.n1588 VSS.n1592 4.5005
R14924 VSS.n1589 VSS.n1593 4.5005
R14925 VSS.n1590 VSS.n1594 4.57324
R14926 VSS.n1586 VSS.n1584 0.147342
R14927 VSS.n1587 VSS.n1588 0.0732424
R14928 VSS.n1588 VSS.n1589 0.147342
R14929 VSS.n1591 VSS.n1595 0.0721009
R14930 VSS.n1596 VSS.n1592 4.5005
R14931 VSS.n1597 VSS.n1593 4.5005
R14932 VSS.n1598 VSS.n1594 4.5005
R14933 VSS.n1584 VSS.n1595 4.57442
R14934 VSS.n1591 VSS.n1592 0.147342
R14935 VSS.n1592 VSS.n1593 0.147342
R14936 VSS.n1593 VSS.n1594 0.147342
R14937 VSS.n1595 VSS.n1596 2.39784
R14938 VSS.n1596 VSS.n1597 0.147342
R14939 VSS.n1597 VSS.n1598 0.147342
R14940 VSS.n1598 VSS.t177 3.13212
R14941 VSS.n1571 VSS.n1576 4.5005
R14942 VSS.n1573 VSS.n1577 4.5005
R14943 VSS.n1574 VSS.n1578 4.5005
R14944 VSS.n1575 VSS.n1579 4.57324
R14945 VSS.n1571 VSS.n1569 0.147342
R14946 VSS.n1572 VSS.n1573 0.0732424
R14947 VSS.n1573 VSS.n1574 0.147342
R14948 VSS.n1576 VSS.n1580 0.0721009
R14949 VSS.n1581 VSS.n1577 4.5005
R14950 VSS.n1582 VSS.n1578 4.5005
R14951 VSS.n1583 VSS.n1579 4.5005
R14952 VSS.n1569 VSS.n1580 4.57442
R14953 VSS.n1576 VSS.n1577 0.147342
R14954 VSS.n1577 VSS.n1578 0.147342
R14955 VSS.n1578 VSS.n1579 0.147342
R14956 VSS.n1580 VSS.n1581 2.39784
R14957 VSS.n1581 VSS.n1582 0.147342
R14958 VSS.n1582 VSS.n1583 0.147342
R14959 VSS.n1583 VSS.t222 3.13212
R14960 VSS.n1556 VSS.n1561 4.5005
R14961 VSS.n1558 VSS.n1562 4.5005
R14962 VSS.n1559 VSS.n1563 4.5005
R14963 VSS.n1560 VSS.n1564 4.57324
R14964 VSS.n1556 VSS.n1554 0.147342
R14965 VSS.n1557 VSS.n1558 0.0732424
R14966 VSS.n1558 VSS.n1559 0.147342
R14967 VSS.n1561 VSS.n1565 0.0721009
R14968 VSS.n1566 VSS.n1562 4.5005
R14969 VSS.n1567 VSS.n1563 4.5005
R14970 VSS.n1568 VSS.n1564 4.5005
R14971 VSS.n1554 VSS.n1565 4.57442
R14972 VSS.n1561 VSS.n1562 0.147342
R14973 VSS.n1562 VSS.n1563 0.147342
R14974 VSS.n1563 VSS.n1564 0.147342
R14975 VSS.n1565 VSS.n1566 2.39784
R14976 VSS.n1566 VSS.n1567 0.147342
R14977 VSS.n1567 VSS.n1568 0.147342
R14978 VSS.n1568 VSS.t306 3.13212
R14979 VSS.n1535 VSS.n1540 4.5005
R14980 VSS.n1537 VSS.n1541 4.5005
R14981 VSS.n1538 VSS.n1542 4.5005
R14982 VSS.n1539 VSS.n1543 4.57324
R14983 VSS.n1535 VSS.n1533 0.147342
R14984 VSS.n1536 VSS.n1537 0.0732424
R14985 VSS.n1537 VSS.n1538 0.147342
R14986 VSS.n1540 VSS.n1544 0.0721009
R14987 VSS.n1545 VSS.n1541 4.5005
R14988 VSS.n1546 VSS.n1542 4.5005
R14989 VSS.n1547 VSS.n1543 4.5005
R14990 VSS.n1533 VSS.n1544 4.57442
R14991 VSS.n1540 VSS.n1541 0.147342
R14992 VSS.n1541 VSS.n1542 0.147342
R14993 VSS.n1542 VSS.n1543 0.147342
R14994 VSS.n1544 VSS.n1545 2.39784
R14995 VSS.n1545 VSS.n1546 0.147342
R14996 VSS.n1546 VSS.n1547 0.147342
R14997 VSS.n1547 VSS.t559 3.13212
R14998 VSS.n1520 VSS.n1525 4.5005
R14999 VSS.n1522 VSS.n1526 4.5005
R15000 VSS.n1523 VSS.n1527 4.5005
R15001 VSS.n1524 VSS.n1528 4.57324
R15002 VSS.n1520 VSS.n1518 0.147342
R15003 VSS.n1521 VSS.n1522 0.0732424
R15004 VSS.n1522 VSS.n1523 0.147342
R15005 VSS.n1525 VSS.n1529 0.0721009
R15006 VSS.n1530 VSS.n1526 4.5005
R15007 VSS.n1531 VSS.n1527 4.5005
R15008 VSS.n1532 VSS.n1528 4.5005
R15009 VSS.n1518 VSS.n1529 4.57442
R15010 VSS.n1525 VSS.n1526 0.147342
R15011 VSS.n1526 VSS.n1527 0.147342
R15012 VSS.n1527 VSS.n1528 0.147342
R15013 VSS.n1529 VSS.n1530 2.39784
R15014 VSS.n1530 VSS.n1531 0.147342
R15015 VSS.n1531 VSS.n1532 0.147342
R15016 VSS.n1532 VSS.t376 3.13212
R15017 VSS.n1505 VSS.n1510 4.5005
R15018 VSS.n1507 VSS.n1511 4.5005
R15019 VSS.n1508 VSS.n1512 4.5005
R15020 VSS.n1509 VSS.n1513 4.57324
R15021 VSS.n1505 VSS.n1503 0.147342
R15022 VSS.n1506 VSS.n1507 0.0732424
R15023 VSS.n1507 VSS.n1508 0.147342
R15024 VSS.n1510 VSS.n1514 0.0721009
R15025 VSS.n1515 VSS.n1511 4.5005
R15026 VSS.n1516 VSS.n1512 4.5005
R15027 VSS.n1517 VSS.n1513 4.5005
R15028 VSS.n1503 VSS.n1514 4.57442
R15029 VSS.n1510 VSS.n1511 0.147342
R15030 VSS.n1511 VSS.n1512 0.147342
R15031 VSS.n1512 VSS.n1513 0.147342
R15032 VSS.n1514 VSS.n1515 2.39784
R15033 VSS.n1515 VSS.n1516 0.147342
R15034 VSS.n1516 VSS.n1517 0.147342
R15035 VSS.n1517 VSS.t597 3.13212
R15036 VSS.n1484 VSS.n1489 4.5005
R15037 VSS.n1486 VSS.n1490 4.5005
R15038 VSS.n1487 VSS.n1491 4.5005
R15039 VSS.n1488 VSS.n1492 4.57324
R15040 VSS.n1484 VSS.n1482 0.147342
R15041 VSS.n1485 VSS.n1486 0.0732424
R15042 VSS.n1486 VSS.n1487 0.147342
R15043 VSS.n1489 VSS.n1493 0.0721009
R15044 VSS.n1494 VSS.n1490 4.5005
R15045 VSS.n1495 VSS.n1491 4.5005
R15046 VSS.n1496 VSS.n1492 4.5005
R15047 VSS.n1482 VSS.n1493 4.57442
R15048 VSS.n1489 VSS.n1490 0.147342
R15049 VSS.n1490 VSS.n1491 0.147342
R15050 VSS.n1491 VSS.n1492 0.147342
R15051 VSS.n1493 VSS.n1494 2.39784
R15052 VSS.n1494 VSS.n1495 0.147342
R15053 VSS.n1495 VSS.n1496 0.147342
R15054 VSS.n1496 VSS.t369 3.13212
R15055 VSS.n1469 VSS.n1474 4.5005
R15056 VSS.n1471 VSS.n1475 4.5005
R15057 VSS.n1472 VSS.n1476 4.5005
R15058 VSS.n1473 VSS.n1477 4.57324
R15059 VSS.n1469 VSS.n1467 0.147342
R15060 VSS.n1470 VSS.n1471 0.0732424
R15061 VSS.n1471 VSS.n1472 0.147342
R15062 VSS.n1474 VSS.n1478 0.0721009
R15063 VSS.n1479 VSS.n1475 4.5005
R15064 VSS.n1480 VSS.n1476 4.5005
R15065 VSS.n1481 VSS.n1477 4.5005
R15066 VSS.n1467 VSS.n1478 4.57442
R15067 VSS.n1474 VSS.n1475 0.147342
R15068 VSS.n1475 VSS.n1476 0.147342
R15069 VSS.n1476 VSS.n1477 0.147342
R15070 VSS.n1478 VSS.n1479 2.39784
R15071 VSS.n1479 VSS.n1480 0.147342
R15072 VSS.n1480 VSS.n1481 0.147342
R15073 VSS.n1481 VSS.t343 3.13212
R15074 VSS.n1454 VSS.n1459 4.5005
R15075 VSS.n1456 VSS.n1460 4.5005
R15076 VSS.n1457 VSS.n1461 4.5005
R15077 VSS.n1458 VSS.n1462 4.57324
R15078 VSS.n1454 VSS.n1452 0.147342
R15079 VSS.n1455 VSS.n1456 0.0732424
R15080 VSS.n1456 VSS.n1457 0.147342
R15081 VSS.n1459 VSS.n1463 0.0721009
R15082 VSS.n1464 VSS.n1460 4.5005
R15083 VSS.n1465 VSS.n1461 4.5005
R15084 VSS.n1466 VSS.n1462 4.5005
R15085 VSS.n1452 VSS.n1463 4.57442
R15086 VSS.n1459 VSS.n1460 0.147342
R15087 VSS.n1460 VSS.n1461 0.147342
R15088 VSS.n1461 VSS.n1462 0.147342
R15089 VSS.n1463 VSS.n1464 2.39784
R15090 VSS.n1464 VSS.n1465 0.147342
R15091 VSS.n1465 VSS.n1466 0.147342
R15092 VSS.n1466 VSS.t429 3.13212
R15093 VSS.n1439 VSS.n1444 4.5005
R15094 VSS.n1441 VSS.n1445 4.5005
R15095 VSS.n1442 VSS.n1446 4.5005
R15096 VSS.n1443 VSS.n1447 4.57324
R15097 VSS.n1439 VSS.n1437 0.147342
R15098 VSS.n1440 VSS.n1441 0.0732424
R15099 VSS.n1441 VSS.n1442 0.147342
R15100 VSS.n1444 VSS.n1448 0.0721009
R15101 VSS.n1449 VSS.n1445 4.5005
R15102 VSS.n1450 VSS.n1446 4.5005
R15103 VSS.n1451 VSS.n1447 4.5005
R15104 VSS.n1437 VSS.n1448 4.57442
R15105 VSS.n1444 VSS.n1445 0.147342
R15106 VSS.n1445 VSS.n1446 0.147342
R15107 VSS.n1446 VSS.n1447 0.147342
R15108 VSS.n1448 VSS.n1449 2.39784
R15109 VSS.n1449 VSS.n1450 0.147342
R15110 VSS.n1450 VSS.n1451 0.147342
R15111 VSS.n1451 VSS.t80 3.13212
R15112 VSS.n1424 VSS.n1429 4.5005
R15113 VSS.n1426 VSS.n1430 4.5005
R15114 VSS.n1427 VSS.n1431 4.5005
R15115 VSS.n1428 VSS.n1432 4.57324
R15116 VSS.n1424 VSS.n1422 0.147342
R15117 VSS.n1425 VSS.n1426 0.0732424
R15118 VSS.n1426 VSS.n1427 0.147342
R15119 VSS.n1429 VSS.n1433 0.0721009
R15120 VSS.n1434 VSS.n1430 4.5005
R15121 VSS.n1435 VSS.n1431 4.5005
R15122 VSS.n1436 VSS.n1432 4.5005
R15123 VSS.n1422 VSS.n1433 4.57442
R15124 VSS.n1429 VSS.n1430 0.147342
R15125 VSS.n1430 VSS.n1431 0.147342
R15126 VSS.n1431 VSS.n1432 0.147342
R15127 VSS.n1433 VSS.n1434 2.39784
R15128 VSS.n1434 VSS.n1435 0.147342
R15129 VSS.n1435 VSS.n1436 0.147342
R15130 VSS.n1436 VSS.t28 3.13212
R15131 VSS.n1409 VSS.n1414 4.5005
R15132 VSS.n1411 VSS.n1415 4.5005
R15133 VSS.n1412 VSS.n1416 4.5005
R15134 VSS.n1413 VSS.n1417 4.57324
R15135 VSS.n1409 VSS.n1407 0.147342
R15136 VSS.n1410 VSS.n1411 0.0732424
R15137 VSS.n1411 VSS.n1412 0.147342
R15138 VSS.n1414 VSS.n1418 0.0721009
R15139 VSS.n1419 VSS.n1415 4.5005
R15140 VSS.n1420 VSS.n1416 4.5005
R15141 VSS.n1421 VSS.n1417 4.5005
R15142 VSS.n1407 VSS.n1418 4.57442
R15143 VSS.n1414 VSS.n1415 0.147342
R15144 VSS.n1415 VSS.n1416 0.147342
R15145 VSS.n1416 VSS.n1417 0.147342
R15146 VSS.n1418 VSS.n1419 2.39784
R15147 VSS.n1419 VSS.n1420 0.147342
R15148 VSS.n1420 VSS.n1421 0.147342
R15149 VSS.n1421 VSS.t353 3.13212
R15150 VSS.n1388 VSS.n1393 4.5005
R15151 VSS.n1390 VSS.n1394 4.5005
R15152 VSS.n1391 VSS.n1395 4.5005
R15153 VSS.n1392 VSS.n1396 4.57324
R15154 VSS.n1388 VSS.n1386 0.147342
R15155 VSS.n1389 VSS.n1390 0.0732424
R15156 VSS.n1390 VSS.n1391 0.147342
R15157 VSS.n1393 VSS.n1397 0.0721009
R15158 VSS.n1398 VSS.n1394 4.5005
R15159 VSS.n1399 VSS.n1395 4.5005
R15160 VSS.n1400 VSS.n1396 4.5005
R15161 VSS.n1386 VSS.n1397 4.57442
R15162 VSS.n1393 VSS.n1394 0.147342
R15163 VSS.n1394 VSS.n1395 0.147342
R15164 VSS.n1395 VSS.n1396 0.147342
R15165 VSS.n1397 VSS.n1398 2.39784
R15166 VSS.n1398 VSS.n1399 0.147342
R15167 VSS.n1399 VSS.n1400 0.147342
R15168 VSS.n1400 VSS.t313 3.13212
R15169 VSS.n1373 VSS.n1378 4.5005
R15170 VSS.n1375 VSS.n1379 4.5005
R15171 VSS.n1376 VSS.n1380 4.5005
R15172 VSS.n1377 VSS.n1381 4.57324
R15173 VSS.n1373 VSS.n1371 0.147342
R15174 VSS.n1374 VSS.n1375 0.0732424
R15175 VSS.n1375 VSS.n1376 0.147342
R15176 VSS.n1378 VSS.n1382 0.0721009
R15177 VSS.n1383 VSS.n1379 4.5005
R15178 VSS.n1384 VSS.n1380 4.5005
R15179 VSS.n1385 VSS.n1381 4.5005
R15180 VSS.n1371 VSS.n1382 4.57442
R15181 VSS.n1378 VSS.n1379 0.147342
R15182 VSS.n1379 VSS.n1380 0.147342
R15183 VSS.n1380 VSS.n1381 0.147342
R15184 VSS.n1382 VSS.n1383 2.39784
R15185 VSS.n1383 VSS.n1384 0.147342
R15186 VSS.n1384 VSS.n1385 0.147342
R15187 VSS.n1385 VSS.t340 3.13212
R15188 VSS.n1358 VSS.n1363 4.5005
R15189 VSS.n1360 VSS.n1364 4.5005
R15190 VSS.n1361 VSS.n1365 4.5005
R15191 VSS.n1362 VSS.n1366 4.57324
R15192 VSS.n1358 VSS.n1356 0.147342
R15193 VSS.n1359 VSS.n1360 0.0732424
R15194 VSS.n1360 VSS.n1361 0.147342
R15195 VSS.n1363 VSS.n1367 0.0721009
R15196 VSS.n1368 VSS.n1364 4.5005
R15197 VSS.n1369 VSS.n1365 4.5005
R15198 VSS.n1370 VSS.n1366 4.5005
R15199 VSS.n1356 VSS.n1367 4.57442
R15200 VSS.n1363 VSS.n1364 0.147342
R15201 VSS.n1364 VSS.n1365 0.147342
R15202 VSS.n1365 VSS.n1366 0.147342
R15203 VSS.n1367 VSS.n1368 2.39784
R15204 VSS.n1368 VSS.n1369 0.147342
R15205 VSS.n1369 VSS.n1370 0.147342
R15206 VSS.n1370 VSS.t323 3.13212
R15207 VSS.n1337 VSS.n1342 4.5005
R15208 VSS.n1339 VSS.n1343 4.5005
R15209 VSS.n1340 VSS.n1344 4.5005
R15210 VSS.n1341 VSS.n1345 4.57324
R15211 VSS.n1337 VSS.n1335 0.147342
R15212 VSS.n1338 VSS.n1339 0.0732424
R15213 VSS.n1339 VSS.n1340 0.147342
R15214 VSS.n1342 VSS.n1346 0.0721009
R15215 VSS.n1347 VSS.n1343 4.5005
R15216 VSS.n1348 VSS.n1344 4.5005
R15217 VSS.n1349 VSS.n1345 4.5005
R15218 VSS.n1335 VSS.n1346 4.57442
R15219 VSS.n1342 VSS.n1343 0.147342
R15220 VSS.n1343 VSS.n1344 0.147342
R15221 VSS.n1344 VSS.n1345 0.147342
R15222 VSS.n1346 VSS.n1347 2.39784
R15223 VSS.n1347 VSS.n1348 0.147342
R15224 VSS.n1348 VSS.n1349 0.147342
R15225 VSS.n1349 VSS.t388 3.13212
R15226 VSS.n1322 VSS.n1327 4.5005
R15227 VSS.n1324 VSS.n1328 4.5005
R15228 VSS.n1325 VSS.n1329 4.5005
R15229 VSS.n1326 VSS.n1330 4.57324
R15230 VSS.n1322 VSS.n1320 0.147342
R15231 VSS.n1323 VSS.n1324 0.0732424
R15232 VSS.n1324 VSS.n1325 0.147342
R15233 VSS.n1327 VSS.n1331 0.0721009
R15234 VSS.n1332 VSS.n1328 4.5005
R15235 VSS.n1333 VSS.n1329 4.5005
R15236 VSS.n1334 VSS.n1330 4.5005
R15237 VSS.n1320 VSS.n1331 4.57442
R15238 VSS.n1327 VSS.n1328 0.147342
R15239 VSS.n1328 VSS.n1329 0.147342
R15240 VSS.n1329 VSS.n1330 0.147342
R15241 VSS.n1331 VSS.n1332 2.39784
R15242 VSS.n1332 VSS.n1333 0.147342
R15243 VSS.n1333 VSS.n1334 0.147342
R15244 VSS.n1334 VSS.t460 3.13212
R15245 VSS.n1307 VSS.n1312 4.5005
R15246 VSS.n1309 VSS.n1313 4.5005
R15247 VSS.n1310 VSS.n1314 4.5005
R15248 VSS.n1311 VSS.n1315 4.57324
R15249 VSS.n1307 VSS.n1305 0.147342
R15250 VSS.n1308 VSS.n1309 0.0732424
R15251 VSS.n1309 VSS.n1310 0.147342
R15252 VSS.n1312 VSS.n1316 0.0721009
R15253 VSS.n1317 VSS.n1313 4.5005
R15254 VSS.n1318 VSS.n1314 4.5005
R15255 VSS.n1319 VSS.n1315 4.5005
R15256 VSS.n1305 VSS.n1316 4.57442
R15257 VSS.n1312 VSS.n1313 0.147342
R15258 VSS.n1313 VSS.n1314 0.147342
R15259 VSS.n1314 VSS.n1315 0.147342
R15260 VSS.n1316 VSS.n1317 2.39784
R15261 VSS.n1317 VSS.n1318 0.147342
R15262 VSS.n1318 VSS.n1319 0.147342
R15263 VSS.n1319 VSS.t219 3.13212
R15264 VSS.n1292 VSS.n1297 4.5005
R15265 VSS.n1294 VSS.n1298 4.5005
R15266 VSS.n1295 VSS.n1299 4.5005
R15267 VSS.n1296 VSS.n1300 4.57324
R15268 VSS.n1292 VSS.n1290 0.147342
R15269 VSS.n1293 VSS.n1294 0.0732424
R15270 VSS.n1294 VSS.n1295 0.147342
R15271 VSS.n1297 VSS.n1301 0.0721009
R15272 VSS.n1302 VSS.n1298 4.5005
R15273 VSS.n1303 VSS.n1299 4.5005
R15274 VSS.n1304 VSS.n1300 4.5005
R15275 VSS.n1290 VSS.n1301 4.57442
R15276 VSS.n1297 VSS.n1298 0.147342
R15277 VSS.n1298 VSS.n1299 0.147342
R15278 VSS.n1299 VSS.n1300 0.147342
R15279 VSS.n1301 VSS.n1302 2.39784
R15280 VSS.n1302 VSS.n1303 0.147342
R15281 VSS.n1303 VSS.n1304 0.147342
R15282 VSS.n1304 VSS.t291 3.13212
R15283 VSS.n1271 VSS.n1276 4.5005
R15284 VSS.n1273 VSS.n1277 4.5005
R15285 VSS.n1274 VSS.n1278 4.5005
R15286 VSS.n1275 VSS.n1279 4.57324
R15287 VSS.n1271 VSS.n1269 0.147342
R15288 VSS.n1272 VSS.n1273 0.0732424
R15289 VSS.n1273 VSS.n1274 0.147342
R15290 VSS.n1276 VSS.n1280 0.0721009
R15291 VSS.n1281 VSS.n1277 4.5005
R15292 VSS.n1282 VSS.n1278 4.5005
R15293 VSS.n1283 VSS.n1279 4.5005
R15294 VSS.n1269 VSS.n1280 4.57442
R15295 VSS.n1276 VSS.n1277 0.147342
R15296 VSS.n1277 VSS.n1278 0.147342
R15297 VSS.n1278 VSS.n1279 0.147342
R15298 VSS.n1280 VSS.n1281 2.39784
R15299 VSS.n1281 VSS.n1282 0.147342
R15300 VSS.n1282 VSS.n1283 0.147342
R15301 VSS.n1283 VSS.t562 3.13212
R15302 VSS.n1256 VSS.n1261 4.5005
R15303 VSS.n1258 VSS.n1262 4.5005
R15304 VSS.n1259 VSS.n1263 4.5005
R15305 VSS.n1260 VSS.n1264 4.57324
R15306 VSS.n1256 VSS.n1254 0.147342
R15307 VSS.n1257 VSS.n1258 0.0732424
R15308 VSS.n1258 VSS.n1259 0.147342
R15309 VSS.n1261 VSS.n1265 0.0721009
R15310 VSS.n1266 VSS.n1262 4.5005
R15311 VSS.n1267 VSS.n1263 4.5005
R15312 VSS.n1268 VSS.n1264 4.5005
R15313 VSS.n1254 VSS.n1265 4.57442
R15314 VSS.n1261 VSS.n1262 0.147342
R15315 VSS.n1262 VSS.n1263 0.147342
R15316 VSS.n1263 VSS.n1264 0.147342
R15317 VSS.n1265 VSS.n1266 2.39784
R15318 VSS.n1266 VSS.n1267 0.147342
R15319 VSS.n1267 VSS.n1268 0.147342
R15320 VSS.n1268 VSS.t379 3.13212
R15321 VSS.n1241 VSS.n1246 4.5005
R15322 VSS.n1243 VSS.n1247 4.5005
R15323 VSS.n1244 VSS.n1248 4.5005
R15324 VSS.n1245 VSS.n1249 4.57324
R15325 VSS.n1241 VSS.n1239 0.147342
R15326 VSS.n1242 VSS.n1243 0.0732424
R15327 VSS.n1243 VSS.n1244 0.147342
R15328 VSS.n1246 VSS.n1250 0.0721009
R15329 VSS.n1251 VSS.n1247 4.5005
R15330 VSS.n1252 VSS.n1248 4.5005
R15331 VSS.n1253 VSS.n1249 4.5005
R15332 VSS.n1239 VSS.n1250 4.57442
R15333 VSS.n1246 VSS.n1247 0.147342
R15334 VSS.n1247 VSS.n1248 0.147342
R15335 VSS.n1248 VSS.n1249 0.147342
R15336 VSS.n1250 VSS.n1251 2.39784
R15337 VSS.n1251 VSS.n1252 0.147342
R15338 VSS.n1252 VSS.n1253 0.147342
R15339 VSS.n1253 VSS.t270 3.13212
R15340 VSS.n1220 VSS.n1225 4.5005
R15341 VSS.n1222 VSS.n1226 4.5005
R15342 VSS.n1223 VSS.n1227 4.5005
R15343 VSS.n1224 VSS.n1228 4.57324
R15344 VSS.n1220 VSS.n1218 0.147342
R15345 VSS.n1221 VSS.n1222 0.0732424
R15346 VSS.n1222 VSS.n1223 0.147342
R15347 VSS.n1225 VSS.n1229 0.0721009
R15348 VSS.n1230 VSS.n1226 4.5005
R15349 VSS.n1231 VSS.n1227 4.5005
R15350 VSS.n1232 VSS.n1228 4.5005
R15351 VSS.n1218 VSS.n1229 4.57442
R15352 VSS.n1225 VSS.n1226 0.147342
R15353 VSS.n1226 VSS.n1227 0.147342
R15354 VSS.n1227 VSS.n1228 0.147342
R15355 VSS.n1229 VSS.n1230 2.39784
R15356 VSS.n1230 VSS.n1231 0.147342
R15357 VSS.n1231 VSS.n1232 0.147342
R15358 VSS.n1232 VSS.t289 3.13212
R15359 VSS.n1205 VSS.n1210 4.5005
R15360 VSS.n1207 VSS.n1211 4.5005
R15361 VSS.n1208 VSS.n1212 4.5005
R15362 VSS.n1209 VSS.n1213 4.57324
R15363 VSS.n1205 VSS.n1203 0.147342
R15364 VSS.n1206 VSS.n1207 0.0732424
R15365 VSS.n1207 VSS.n1208 0.147342
R15366 VSS.n1210 VSS.n1214 0.0721009
R15367 VSS.n1215 VSS.n1211 4.5005
R15368 VSS.n1216 VSS.n1212 4.5005
R15369 VSS.n1217 VSS.n1213 4.5005
R15370 VSS.n1203 VSS.n1214 4.57442
R15371 VSS.n1210 VSS.n1211 0.147342
R15372 VSS.n1211 VSS.n1212 0.147342
R15373 VSS.n1212 VSS.n1213 0.147342
R15374 VSS.n1214 VSS.n1215 2.39784
R15375 VSS.n1215 VSS.n1216 0.147342
R15376 VSS.n1216 VSS.n1217 0.147342
R15377 VSS.n1217 VSS.t579 3.13212
R15378 VSS.n1190 VSS.n1195 4.5005
R15379 VSS.n1192 VSS.n1196 4.5005
R15380 VSS.n1193 VSS.n1197 4.5005
R15381 VSS.n1194 VSS.n1198 4.57324
R15382 VSS.n1190 VSS.n1188 0.147342
R15383 VSS.n1191 VSS.n1192 0.0732424
R15384 VSS.n1192 VSS.n1193 0.147342
R15385 VSS.n1195 VSS.n1199 0.0721009
R15386 VSS.n1200 VSS.n1196 4.5005
R15387 VSS.n1201 VSS.n1197 4.5005
R15388 VSS.n1202 VSS.n1198 4.5005
R15389 VSS.n1188 VSS.n1199 4.57442
R15390 VSS.n1195 VSS.n1196 0.147342
R15391 VSS.n1196 VSS.n1197 0.147342
R15392 VSS.n1197 VSS.n1198 0.147342
R15393 VSS.n1199 VSS.n1200 2.39784
R15394 VSS.n1200 VSS.n1201 0.147342
R15395 VSS.n1201 VSS.n1202 0.147342
R15396 VSS.n1202 VSS.t152 3.13212
R15397 VSS.n1175 VSS.n1180 4.5005
R15398 VSS.n1177 VSS.n1181 4.5005
R15399 VSS.n1178 VSS.n1182 4.5005
R15400 VSS.n1179 VSS.n1183 4.57324
R15401 VSS.n1175 VSS.n1173 0.147342
R15402 VSS.n1176 VSS.n1177 0.0732424
R15403 VSS.n1177 VSS.n1178 0.147342
R15404 VSS.n1180 VSS.n1184 0.0721009
R15405 VSS.n1185 VSS.n1181 4.5005
R15406 VSS.n1186 VSS.n1182 4.5005
R15407 VSS.n1187 VSS.n1183 4.5005
R15408 VSS.n1173 VSS.n1184 4.57442
R15409 VSS.n1180 VSS.n1181 0.147342
R15410 VSS.n1181 VSS.n1182 0.147342
R15411 VSS.n1182 VSS.n1183 0.147342
R15412 VSS.n1184 VSS.n1185 2.39784
R15413 VSS.n1185 VSS.n1186 0.147342
R15414 VSS.n1186 VSS.n1187 0.147342
R15415 VSS.n1187 VSS.t83 3.13212
R15416 VSS.n1160 VSS.n1165 4.5005
R15417 VSS.n1162 VSS.n1166 4.5005
R15418 VSS.n1163 VSS.n1167 4.5005
R15419 VSS.n1164 VSS.n1168 4.57324
R15420 VSS.n1160 VSS.n1158 0.147342
R15421 VSS.n1161 VSS.n1162 0.0732424
R15422 VSS.n1162 VSS.n1163 0.147342
R15423 VSS.n1165 VSS.n1169 0.0721009
R15424 VSS.n1170 VSS.n1166 4.5005
R15425 VSS.n1171 VSS.n1167 4.5005
R15426 VSS.n1172 VSS.n1168 4.5005
R15427 VSS.n1158 VSS.n1169 4.57442
R15428 VSS.n1165 VSS.n1166 0.147342
R15429 VSS.n1166 VSS.n1167 0.147342
R15430 VSS.n1167 VSS.n1168 0.147342
R15431 VSS.n1169 VSS.n1170 2.39784
R15432 VSS.n1170 VSS.n1171 0.147342
R15433 VSS.n1171 VSS.n1172 0.147342
R15434 VSS.n1172 VSS.t23 3.13212
R15435 VSS.n1145 VSS.n1150 4.5005
R15436 VSS.n1147 VSS.n1151 4.5005
R15437 VSS.n1148 VSS.n1152 4.5005
R15438 VSS.n1149 VSS.n1153 4.57324
R15439 VSS.n1145 VSS.n1143 0.147342
R15440 VSS.n1146 VSS.n1147 0.0732424
R15441 VSS.n1147 VSS.n1148 0.147342
R15442 VSS.n1150 VSS.n1154 0.0721009
R15443 VSS.n1155 VSS.n1151 4.5005
R15444 VSS.n1156 VSS.n1152 4.5005
R15445 VSS.n1157 VSS.n1153 4.5005
R15446 VSS.n1143 VSS.n1154 4.57442
R15447 VSS.n1150 VSS.n1151 0.147342
R15448 VSS.n1151 VSS.n1152 0.147342
R15449 VSS.n1152 VSS.n1153 0.147342
R15450 VSS.n1154 VSS.n1155 2.39784
R15451 VSS.n1155 VSS.n1156 0.147342
R15452 VSS.n1156 VSS.n1157 0.147342
R15453 VSS.n1157 VSS.t356 3.13212
R15454 VSS.n1124 VSS.n1129 4.5005
R15455 VSS.n1126 VSS.n1130 4.5005
R15456 VSS.n1127 VSS.n1131 4.5005
R15457 VSS.n1128 VSS.n1132 4.57324
R15458 VSS.n1124 VSS.n1122 0.147342
R15459 VSS.n1125 VSS.n1126 0.0732424
R15460 VSS.n1126 VSS.n1127 0.147342
R15461 VSS.n1129 VSS.n1133 0.0721009
R15462 VSS.n1134 VSS.n1130 4.5005
R15463 VSS.n1135 VSS.n1131 4.5005
R15464 VSS.n1136 VSS.n1132 4.5005
R15465 VSS.n1122 VSS.n1133 4.57442
R15466 VSS.n1129 VSS.n1130 0.147342
R15467 VSS.n1130 VSS.n1131 0.147342
R15468 VSS.n1131 VSS.n1132 0.147342
R15469 VSS.n1133 VSS.n1134 2.39784
R15470 VSS.n1134 VSS.n1135 0.147342
R15471 VSS.n1135 VSS.n1136 0.147342
R15472 VSS.n1136 VSS.t317 3.13212
R15473 VSS.n1109 VSS.n1114 4.5005
R15474 VSS.n1111 VSS.n1115 4.5005
R15475 VSS.n1112 VSS.n1116 4.5005
R15476 VSS.n1113 VSS.n1117 4.57324
R15477 VSS.n1109 VSS.n1107 0.147342
R15478 VSS.n1110 VSS.n1111 0.0732424
R15479 VSS.n1111 VSS.n1112 0.147342
R15480 VSS.n1114 VSS.n1118 0.0721009
R15481 VSS.n1119 VSS.n1115 4.5005
R15482 VSS.n1120 VSS.n1116 4.5005
R15483 VSS.n1121 VSS.n1117 4.5005
R15484 VSS.n1107 VSS.n1118 4.57442
R15485 VSS.n1114 VSS.n1115 0.147342
R15486 VSS.n1115 VSS.n1116 0.147342
R15487 VSS.n1116 VSS.n1117 0.147342
R15488 VSS.n1118 VSS.n1119 2.39784
R15489 VSS.n1119 VSS.n1120 0.147342
R15490 VSS.n1120 VSS.n1121 0.147342
R15491 VSS.n1121 VSS.t341 3.13212
R15492 VSS.n1094 VSS.n1099 4.5005
R15493 VSS.n1096 VSS.n1100 4.5005
R15494 VSS.n1097 VSS.n1101 4.5005
R15495 VSS.n1098 VSS.n1102 4.57324
R15496 VSS.n1094 VSS.n1092 0.147342
R15497 VSS.n1095 VSS.n1096 0.0732424
R15498 VSS.n1096 VSS.n1097 0.147342
R15499 VSS.n1099 VSS.n1103 0.0721009
R15500 VSS.n1104 VSS.n1100 4.5005
R15501 VSS.n1105 VSS.n1101 4.5005
R15502 VSS.n1106 VSS.n1102 4.5005
R15503 VSS.n1092 VSS.n1103 4.57442
R15504 VSS.n1099 VSS.n1100 0.147342
R15505 VSS.n1100 VSS.n1101 0.147342
R15506 VSS.n1101 VSS.n1102 0.147342
R15507 VSS.n1103 VSS.n1104 2.39784
R15508 VSS.n1104 VSS.n1105 0.147342
R15509 VSS.n1105 VSS.n1106 0.147342
R15510 VSS.n1106 VSS.t392 3.13212
R15511 VSS.n1073 VSS.n1078 4.5005
R15512 VSS.n1075 VSS.n1079 4.5005
R15513 VSS.n1076 VSS.n1080 4.5005
R15514 VSS.n1077 VSS.n1081 4.57324
R15515 VSS.n1073 VSS.n1071 0.147342
R15516 VSS.n1074 VSS.n1075 0.0732424
R15517 VSS.n1075 VSS.n1076 0.147342
R15518 VSS.n1078 VSS.n1082 0.0721009
R15519 VSS.n1083 VSS.n1079 4.5005
R15520 VSS.n1084 VSS.n1080 4.5005
R15521 VSS.n1085 VSS.n1081 4.5005
R15522 VSS.n1071 VSS.n1082 4.57442
R15523 VSS.n1078 VSS.n1079 0.147342
R15524 VSS.n1079 VSS.n1080 0.147342
R15525 VSS.n1080 VSS.n1081 0.147342
R15526 VSS.n1082 VSS.n1083 2.39784
R15527 VSS.n1083 VSS.n1084 0.147342
R15528 VSS.n1084 VSS.n1085 0.147342
R15529 VSS.n1085 VSS.t384 3.13212
R15530 VSS.n1058 VSS.n1063 4.5005
R15531 VSS.n1060 VSS.n1064 4.5005
R15532 VSS.n1061 VSS.n1065 4.5005
R15533 VSS.n1062 VSS.n1066 4.57324
R15534 VSS.n1058 VSS.n1056 0.147342
R15535 VSS.n1059 VSS.n1060 0.0732424
R15536 VSS.n1060 VSS.n1061 0.147342
R15537 VSS.n1063 VSS.n1067 0.0721009
R15538 VSS.n1068 VSS.n1064 4.5005
R15539 VSS.n1069 VSS.n1065 4.5005
R15540 VSS.n1070 VSS.n1066 4.5005
R15541 VSS.n1056 VSS.n1067 4.57442
R15542 VSS.n1063 VSS.n1064 0.147342
R15543 VSS.n1064 VSS.n1065 0.147342
R15544 VSS.n1065 VSS.n1066 0.147342
R15545 VSS.n1067 VSS.n1068 2.39784
R15546 VSS.n1068 VSS.n1069 0.147342
R15547 VSS.n1069 VSS.n1070 0.147342
R15548 VSS.n1070 VSS.t462 3.13212
R15549 VSS.n1043 VSS.n1048 4.5005
R15550 VSS.n1045 VSS.n1049 4.5005
R15551 VSS.n1046 VSS.n1050 4.5005
R15552 VSS.n1047 VSS.n1051 4.57324
R15553 VSS.n1043 VSS.n1041 0.147342
R15554 VSS.n1044 VSS.n1045 0.0732424
R15555 VSS.n1045 VSS.n1046 0.147342
R15556 VSS.n1048 VSS.n1052 0.0721009
R15557 VSS.n1053 VSS.n1049 4.5005
R15558 VSS.n1054 VSS.n1050 4.5005
R15559 VSS.n1055 VSS.n1051 4.5005
R15560 VSS.n1041 VSS.n1052 4.57442
R15561 VSS.n1048 VSS.n1049 0.147342
R15562 VSS.n1049 VSS.n1050 0.147342
R15563 VSS.n1050 VSS.n1051 0.147342
R15564 VSS.n1052 VSS.n1053 2.39784
R15565 VSS.n1053 VSS.n1054 0.147342
R15566 VSS.n1054 VSS.n1055 0.147342
R15567 VSS.n1055 VSS.t223 3.13212
R15568 VSS.n1028 VSS.n1033 4.5005
R15569 VSS.n1030 VSS.n1034 4.5005
R15570 VSS.n1031 VSS.n1035 4.5005
R15571 VSS.n1032 VSS.n1036 4.57324
R15572 VSS.n1028 VSS.n1026 0.147342
R15573 VSS.n1029 VSS.n1030 0.0732424
R15574 VSS.n1030 VSS.n1031 0.147342
R15575 VSS.n1033 VSS.n1037 0.0721009
R15576 VSS.n1038 VSS.n1034 4.5005
R15577 VSS.n1039 VSS.n1035 4.5005
R15578 VSS.n1040 VSS.n1036 4.5005
R15579 VSS.n1026 VSS.n1037 4.57442
R15580 VSS.n1033 VSS.n1034 0.147342
R15581 VSS.n1034 VSS.n1035 0.147342
R15582 VSS.n1035 VSS.n1036 0.147342
R15583 VSS.n1037 VSS.n1038 2.39784
R15584 VSS.n1038 VSS.n1039 0.147342
R15585 VSS.n1039 VSS.n1040 0.147342
R15586 VSS.n1040 VSS.t293 3.13212
R15587 VSS.n1007 VSS.n1012 4.5005
R15588 VSS.n1009 VSS.n1013 4.5005
R15589 VSS.n1010 VSS.n1014 4.5005
R15590 VSS.n1011 VSS.n1015 4.57324
R15591 VSS.n1007 VSS.n1005 0.147342
R15592 VSS.n1008 VSS.n1009 0.0732424
R15593 VSS.n1009 VSS.n1010 0.147342
R15594 VSS.n1012 VSS.n1016 0.0721009
R15595 VSS.n1017 VSS.n1013 4.5005
R15596 VSS.n1018 VSS.n1014 4.5005
R15597 VSS.n1019 VSS.n1015 4.5005
R15598 VSS.n1005 VSS.n1016 4.57442
R15599 VSS.n1012 VSS.n1013 0.147342
R15600 VSS.n1013 VSS.n1014 0.147342
R15601 VSS.n1014 VSS.n1015 0.147342
R15602 VSS.n1016 VSS.n1017 2.39784
R15603 VSS.n1017 VSS.n1018 0.147342
R15604 VSS.n1018 VSS.n1019 0.147342
R15605 VSS.n1019 VSS.t433 3.13212
R15606 VSS.n992 VSS.n997 4.5005
R15607 VSS.n994 VSS.n998 4.5005
R15608 VSS.n995 VSS.n999 4.5005
R15609 VSS.n996 VSS.n1000 4.57324
R15610 VSS.n992 VSS.n990 0.147342
R15611 VSS.n993 VSS.n994 0.0732424
R15612 VSS.n994 VSS.n995 0.147342
R15613 VSS.n997 VSS.n1001 0.0721009
R15614 VSS.n1002 VSS.n998 4.5005
R15615 VSS.n1003 VSS.n999 4.5005
R15616 VSS.n1004 VSS.n1000 4.5005
R15617 VSS.n990 VSS.n1001 4.57442
R15618 VSS.n997 VSS.n998 0.147342
R15619 VSS.n998 VSS.n999 0.147342
R15620 VSS.n999 VSS.n1000 0.147342
R15621 VSS.n1001 VSS.n1002 2.39784
R15622 VSS.n1002 VSS.n1003 0.147342
R15623 VSS.n1003 VSS.n1004 0.147342
R15624 VSS.n1004 VSS.t374 3.13212
R15625 VSS.n977 VSS.n982 4.5005
R15626 VSS.n979 VSS.n983 4.5005
R15627 VSS.n980 VSS.n984 4.5005
R15628 VSS.n981 VSS.n985 4.57324
R15629 VSS.n977 VSS.n975 0.147342
R15630 VSS.n978 VSS.n979 0.0732424
R15631 VSS.n979 VSS.n980 0.147342
R15632 VSS.n982 VSS.n986 0.0721009
R15633 VSS.n987 VSS.n983 4.5005
R15634 VSS.n988 VSS.n984 4.5005
R15635 VSS.n989 VSS.n985 4.5005
R15636 VSS.n975 VSS.n986 4.57442
R15637 VSS.n982 VSS.n983 0.147342
R15638 VSS.n983 VSS.n984 0.147342
R15639 VSS.n984 VSS.n985 0.147342
R15640 VSS.n986 VSS.n987 2.39784
R15641 VSS.n987 VSS.n988 0.147342
R15642 VSS.n988 VSS.n989 0.147342
R15643 VSS.n989 VSS.t271 3.13212
R15644 VSS.n956 VSS.n961 4.5005
R15645 VSS.n958 VSS.n962 4.5005
R15646 VSS.n959 VSS.n963 4.5005
R15647 VSS.n960 VSS.n964 4.57324
R15648 VSS.n956 VSS.n954 0.147342
R15649 VSS.n957 VSS.n958 0.0732424
R15650 VSS.n958 VSS.n959 0.147342
R15651 VSS.n961 VSS.n965 0.0721009
R15652 VSS.n966 VSS.n962 4.5005
R15653 VSS.n967 VSS.n963 4.5005
R15654 VSS.n968 VSS.n964 4.5005
R15655 VSS.n954 VSS.n965 4.57442
R15656 VSS.n961 VSS.n962 0.147342
R15657 VSS.n962 VSS.n963 0.147342
R15658 VSS.n963 VSS.n964 0.147342
R15659 VSS.n965 VSS.n966 2.39784
R15660 VSS.n966 VSS.n967 0.147342
R15661 VSS.n967 VSS.n968 0.147342
R15662 VSS.n968 VSS.t367 3.13212
R15663 VSS.n941 VSS.n946 4.5005
R15664 VSS.n943 VSS.n947 4.5005
R15665 VSS.n944 VSS.n948 4.5005
R15666 VSS.n945 VSS.n949 4.57324
R15667 VSS.n941 VSS.n939 0.147342
R15668 VSS.n942 VSS.n943 0.0732424
R15669 VSS.n943 VSS.n944 0.147342
R15670 VSS.n946 VSS.n950 0.0721009
R15671 VSS.n951 VSS.n947 4.5005
R15672 VSS.n952 VSS.n948 4.5005
R15673 VSS.n953 VSS.n949 4.5005
R15674 VSS.n939 VSS.n950 4.57442
R15675 VSS.n946 VSS.n947 0.147342
R15676 VSS.n947 VSS.n948 0.147342
R15677 VSS.n948 VSS.n949 0.147342
R15678 VSS.n950 VSS.n951 2.39784
R15679 VSS.n951 VSS.n952 0.147342
R15680 VSS.n952 VSS.n953 0.147342
R15681 VSS.n953 VSS.t580 3.13212
R15682 VSS.n926 VSS.n931 4.5005
R15683 VSS.n928 VSS.n932 4.5005
R15684 VSS.n929 VSS.n933 4.5005
R15685 VSS.n930 VSS.n934 4.57324
R15686 VSS.n926 VSS.n924 0.147342
R15687 VSS.n927 VSS.n928 0.0732424
R15688 VSS.n928 VSS.n929 0.147342
R15689 VSS.n931 VSS.n935 0.0721009
R15690 VSS.n936 VSS.n932 4.5005
R15691 VSS.n937 VSS.n933 4.5005
R15692 VSS.n938 VSS.n934 4.5005
R15693 VSS.n924 VSS.n935 4.57442
R15694 VSS.n931 VSS.n932 0.147342
R15695 VSS.n932 VSS.n933 0.147342
R15696 VSS.n933 VSS.n934 0.147342
R15697 VSS.n935 VSS.n936 2.39784
R15698 VSS.n936 VSS.n937 0.147342
R15699 VSS.n937 VSS.n938 0.147342
R15700 VSS.n938 VSS.t275 3.13212
R15701 VSS.n911 VSS.n916 4.5005
R15702 VSS.n913 VSS.n917 4.5005
R15703 VSS.n914 VSS.n918 4.5005
R15704 VSS.n915 VSS.n919 4.57324
R15705 VSS.n911 VSS.n909 0.147342
R15706 VSS.n912 VSS.n913 0.0732424
R15707 VSS.n913 VSS.n914 0.147342
R15708 VSS.n916 VSS.n920 0.0721009
R15709 VSS.n921 VSS.n917 4.5005
R15710 VSS.n922 VSS.n918 4.5005
R15711 VSS.n923 VSS.n919 4.5005
R15712 VSS.n909 VSS.n920 4.57442
R15713 VSS.n916 VSS.n917 0.147342
R15714 VSS.n917 VSS.n918 0.147342
R15715 VSS.n918 VSS.n919 0.147342
R15716 VSS.n920 VSS.n921 2.39784
R15717 VSS.n921 VSS.n922 0.147342
R15718 VSS.n922 VSS.n923 0.147342
R15719 VSS.n923 VSS.t84 3.13212
R15720 VSS.n896 VSS.n901 4.5005
R15721 VSS.n898 VSS.n902 4.5005
R15722 VSS.n899 VSS.n903 4.5005
R15723 VSS.n900 VSS.n904 4.57324
R15724 VSS.n896 VSS.n894 0.147342
R15725 VSS.n897 VSS.n898 0.0732424
R15726 VSS.n898 VSS.n899 0.147342
R15727 VSS.n901 VSS.n905 0.0721009
R15728 VSS.n906 VSS.n902 4.5005
R15729 VSS.n907 VSS.n903 4.5005
R15730 VSS.n908 VSS.n904 4.5005
R15731 VSS.n894 VSS.n905 4.57442
R15732 VSS.n901 VSS.n902 0.147342
R15733 VSS.n902 VSS.n903 0.147342
R15734 VSS.n903 VSS.n904 0.147342
R15735 VSS.n905 VSS.n906 2.39784
R15736 VSS.n906 VSS.n907 0.147342
R15737 VSS.n907 VSS.n908 0.147342
R15738 VSS.n908 VSS.t22 3.13212
R15739 VSS.n881 VSS.n886 4.5005
R15740 VSS.n883 VSS.n887 4.5005
R15741 VSS.n884 VSS.n888 4.5005
R15742 VSS.n885 VSS.n889 4.57324
R15743 VSS.n881 VSS.n879 0.147342
R15744 VSS.n882 VSS.n883 0.0732424
R15745 VSS.n883 VSS.n884 0.147342
R15746 VSS.n886 VSS.n890 0.0721009
R15747 VSS.n891 VSS.n887 4.5005
R15748 VSS.n892 VSS.n888 4.5005
R15749 VSS.n893 VSS.n889 4.5005
R15750 VSS.n879 VSS.n890 4.57442
R15751 VSS.n886 VSS.n887 0.147342
R15752 VSS.n887 VSS.n888 0.147342
R15753 VSS.n888 VSS.n889 0.147342
R15754 VSS.n890 VSS.n891 2.39784
R15755 VSS.n891 VSS.n892 0.147342
R15756 VSS.n892 VSS.n893 0.147342
R15757 VSS.n893 VSS.t505 3.13212
R15758 VSS.n860 VSS.n865 4.5005
R15759 VSS.n862 VSS.n866 4.5005
R15760 VSS.n863 VSS.n867 4.5005
R15761 VSS.n864 VSS.n868 4.57324
R15762 VSS.n860 VSS.n858 0.147342
R15763 VSS.n861 VSS.n862 0.0732424
R15764 VSS.n862 VSS.n863 0.147342
R15765 VSS.n865 VSS.n869 0.0721009
R15766 VSS.n870 VSS.n866 4.5005
R15767 VSS.n871 VSS.n867 4.5005
R15768 VSS.n872 VSS.n868 4.5005
R15769 VSS.n858 VSS.n869 4.57442
R15770 VSS.n865 VSS.n866 0.147342
R15771 VSS.n866 VSS.n867 0.147342
R15772 VSS.n867 VSS.n868 0.147342
R15773 VSS.n869 VSS.n870 2.39784
R15774 VSS.n870 VSS.n871 0.147342
R15775 VSS.n871 VSS.n872 0.147342
R15776 VSS.n872 VSS.t357 3.13212
R15777 VSS.n845 VSS.n850 4.5005
R15778 VSS.n847 VSS.n851 4.5005
R15779 VSS.n848 VSS.n852 4.5005
R15780 VSS.n849 VSS.n853 4.57324
R15781 VSS.n845 VSS.n843 0.147342
R15782 VSS.n846 VSS.n847 0.0732424
R15783 VSS.n847 VSS.n848 0.147342
R15784 VSS.n850 VSS.n854 0.0721009
R15785 VSS.n855 VSS.n851 4.5005
R15786 VSS.n856 VSS.n852 4.5005
R15787 VSS.n857 VSS.n853 4.5005
R15788 VSS.n843 VSS.n854 4.57442
R15789 VSS.n850 VSS.n851 0.147342
R15790 VSS.n851 VSS.n852 0.147342
R15791 VSS.n852 VSS.n853 0.147342
R15792 VSS.n854 VSS.n855 2.39784
R15793 VSS.n855 VSS.n856 0.147342
R15794 VSS.n856 VSS.n857 0.147342
R15795 VSS.n857 VSS.t342 3.13212
R15796 VSS.n830 VSS.n835 4.5005
R15797 VSS.n832 VSS.n836 4.5005
R15798 VSS.n833 VSS.n837 4.5005
R15799 VSS.n834 VSS.n838 4.57324
R15800 VSS.n830 VSS.n828 0.147342
R15801 VSS.n831 VSS.n832 0.0732424
R15802 VSS.n832 VSS.n833 0.147342
R15803 VSS.n835 VSS.n839 0.0721009
R15804 VSS.n840 VSS.n836 4.5005
R15805 VSS.n841 VSS.n837 4.5005
R15806 VSS.n842 VSS.n838 4.5005
R15807 VSS.n828 VSS.n839 4.57442
R15808 VSS.n835 VSS.n836 0.147342
R15809 VSS.n836 VSS.n837 0.147342
R15810 VSS.n837 VSS.n838 0.147342
R15811 VSS.n839 VSS.n840 2.39784
R15812 VSS.n840 VSS.n841 0.147342
R15813 VSS.n841 VSS.n842 0.147342
R15814 VSS.n842 VSS.t320 3.13212
R15815 VSS.n809 VSS.n814 4.5005
R15816 VSS.n811 VSS.n815 4.5005
R15817 VSS.n812 VSS.n816 4.5005
R15818 VSS.n813 VSS.n817 4.57324
R15819 VSS.n809 VSS.n807 0.147342
R15820 VSS.n810 VSS.n811 0.0732424
R15821 VSS.n811 VSS.n812 0.147342
R15822 VSS.n814 VSS.n818 0.0721009
R15823 VSS.n819 VSS.n815 4.5005
R15824 VSS.n820 VSS.n816 4.5005
R15825 VSS.n821 VSS.n817 4.5005
R15826 VSS.n807 VSS.n818 4.57442
R15827 VSS.n814 VSS.n815 0.147342
R15828 VSS.n815 VSS.n816 0.147342
R15829 VSS.n816 VSS.n817 0.147342
R15830 VSS.n818 VSS.n819 2.39784
R15831 VSS.n819 VSS.n820 0.147342
R15832 VSS.n820 VSS.n821 0.147342
R15833 VSS.n821 VSS.t382 3.13212
R15834 VSS.n794 VSS.n799 4.5005
R15835 VSS.n796 VSS.n800 4.5005
R15836 VSS.n797 VSS.n801 4.5005
R15837 VSS.n798 VSS.n802 4.57324
R15838 VSS.n794 VSS.n792 0.147342
R15839 VSS.n795 VSS.n796 0.0732424
R15840 VSS.n796 VSS.n797 0.147342
R15841 VSS.n799 VSS.n803 0.0721009
R15842 VSS.n804 VSS.n800 4.5005
R15843 VSS.n805 VSS.n801 4.5005
R15844 VSS.n806 VSS.n802 4.5005
R15845 VSS.n792 VSS.n803 4.57442
R15846 VSS.n799 VSS.n800 0.147342
R15847 VSS.n800 VSS.n801 0.147342
R15848 VSS.n801 VSS.n802 0.147342
R15849 VSS.n803 VSS.n804 2.39784
R15850 VSS.n804 VSS.n805 0.147342
R15851 VSS.n805 VSS.n806 0.147342
R15852 VSS.n806 VSS.t176 3.13212
R15853 VSS.n779 VSS.n784 4.5005
R15854 VSS.n781 VSS.n785 4.5005
R15855 VSS.n782 VSS.n786 4.5005
R15856 VSS.n783 VSS.n787 4.57324
R15857 VSS.n779 VSS.n777 0.147342
R15858 VSS.n780 VSS.n781 0.0732424
R15859 VSS.n781 VSS.n782 0.147342
R15860 VSS.n784 VSS.n788 0.0721009
R15861 VSS.n789 VSS.n785 4.5005
R15862 VSS.n790 VSS.n786 4.5005
R15863 VSS.n791 VSS.n787 4.5005
R15864 VSS.n777 VSS.n788 4.57442
R15865 VSS.n784 VSS.n785 0.147342
R15866 VSS.n785 VSS.n786 0.147342
R15867 VSS.n786 VSS.n787 0.147342
R15868 VSS.n788 VSS.n789 2.39784
R15869 VSS.n789 VSS.n790 0.147342
R15870 VSS.n790 VSS.n791 0.147342
R15871 VSS.n791 VSS.t226 3.13212
R15872 VSS.n764 VSS.n769 4.5005
R15873 VSS.n766 VSS.n770 4.5005
R15874 VSS.n767 VSS.n771 4.5005
R15875 VSS.n768 VSS.n772 4.57324
R15876 VSS.n764 VSS.n762 0.147342
R15877 VSS.n765 VSS.n766 0.0732424
R15878 VSS.n766 VSS.n767 0.147342
R15879 VSS.n769 VSS.n773 0.0721009
R15880 VSS.n774 VSS.n770 4.5005
R15881 VSS.n775 VSS.n771 4.5005
R15882 VSS.n776 VSS.n772 4.5005
R15883 VSS.n762 VSS.n773 4.57442
R15884 VSS.n769 VSS.n770 0.147342
R15885 VSS.n770 VSS.n771 0.147342
R15886 VSS.n771 VSS.n772 0.147342
R15887 VSS.n773 VSS.n774 2.39784
R15888 VSS.n774 VSS.n775 0.147342
R15889 VSS.n775 VSS.n776 0.147342
R15890 VSS.n776 VSS.t303 3.13212
R15891 VSS.n743 VSS.n748 4.5005
R15892 VSS.n745 VSS.n749 4.5005
R15893 VSS.n746 VSS.n750 4.5005
R15894 VSS.n747 VSS.n751 4.57324
R15895 VSS.n743 VSS.n741 0.147342
R15896 VSS.n744 VSS.n745 0.0732424
R15897 VSS.n745 VSS.n746 0.147342
R15898 VSS.n748 VSS.n752 0.0721009
R15899 VSS.n753 VSS.n749 4.5005
R15900 VSS.n754 VSS.n750 4.5005
R15901 VSS.n755 VSS.n751 4.5005
R15902 VSS.n741 VSS.n752 4.57442
R15903 VSS.n748 VSS.n749 0.147342
R15904 VSS.n749 VSS.n750 0.147342
R15905 VSS.n750 VSS.n751 0.147342
R15906 VSS.n752 VSS.n753 2.39784
R15907 VSS.n753 VSS.n754 0.147342
R15908 VSS.n754 VSS.n755 0.147342
R15909 VSS.n755 VSS.t563 3.13212
R15910 VSS.n728 VSS.n733 4.5005
R15911 VSS.n730 VSS.n734 4.5005
R15912 VSS.n731 VSS.n735 4.5005
R15913 VSS.n732 VSS.n736 4.57324
R15914 VSS.n728 VSS.n726 0.147342
R15915 VSS.n729 VSS.n730 0.0732424
R15916 VSS.n730 VSS.n731 0.147342
R15917 VSS.n733 VSS.n737 0.0721009
R15918 VSS.n738 VSS.n734 4.5005
R15919 VSS.n739 VSS.n735 4.5005
R15920 VSS.n740 VSS.n736 4.5005
R15921 VSS.n726 VSS.n737 4.57442
R15922 VSS.n733 VSS.n734 0.147342
R15923 VSS.n734 VSS.n735 0.147342
R15924 VSS.n735 VSS.n736 0.147342
R15925 VSS.n737 VSS.n738 2.39784
R15926 VSS.n738 VSS.n739 0.147342
R15927 VSS.n739 VSS.n740 0.147342
R15928 VSS.n740 VSS.t372 3.13212
R15929 VSS.n713 VSS.n718 4.5005
R15930 VSS.n715 VSS.n719 4.5005
R15931 VSS.n716 VSS.n720 4.5005
R15932 VSS.n717 VSS.n721 4.57324
R15933 VSS.n713 VSS.n711 0.147342
R15934 VSS.n714 VSS.n715 0.0732424
R15935 VSS.n715 VSS.n716 0.147342
R15936 VSS.n718 VSS.n722 0.0721009
R15937 VSS.n723 VSS.n719 4.5005
R15938 VSS.n724 VSS.n720 4.5005
R15939 VSS.n725 VSS.n721 4.5005
R15940 VSS.n711 VSS.n722 4.57442
R15941 VSS.n718 VSS.n719 0.147342
R15942 VSS.n719 VSS.n720 0.147342
R15943 VSS.n720 VSS.n721 0.147342
R15944 VSS.n722 VSS.n723 2.39784
R15945 VSS.n723 VSS.n724 0.147342
R15946 VSS.n724 VSS.n725 0.147342
R15947 VSS.n725 VSS.t593 3.13212
R15948 VSS.n692 VSS.n697 4.5005
R15949 VSS.n694 VSS.n698 4.5005
R15950 VSS.n695 VSS.n699 4.5005
R15951 VSS.n696 VSS.n700 4.57324
R15952 VSS.n692 VSS.n690 0.147342
R15953 VSS.n693 VSS.n694 0.0732424
R15954 VSS.n694 VSS.n695 0.147342
R15955 VSS.n697 VSS.n701 0.0721009
R15956 VSS.n702 VSS.n698 4.5005
R15957 VSS.n703 VSS.n699 4.5005
R15958 VSS.n704 VSS.n700 4.5005
R15959 VSS.n690 VSS.n701 4.57442
R15960 VSS.n697 VSS.n698 0.147342
R15961 VSS.n698 VSS.n699 0.147342
R15962 VSS.n699 VSS.n700 0.147342
R15963 VSS.n701 VSS.n702 2.39784
R15964 VSS.n702 VSS.n703 0.147342
R15965 VSS.n703 VSS.n704 0.147342
R15966 VSS.n704 VSS.t370 3.13212
R15967 VSS.n677 VSS.n682 4.5005
R15968 VSS.n679 VSS.n683 4.5005
R15969 VSS.n680 VSS.n684 4.5005
R15970 VSS.n681 VSS.n685 4.57324
R15971 VSS.n677 VSS.n675 0.147342
R15972 VSS.n678 VSS.n679 0.0732424
R15973 VSS.n679 VSS.n680 0.147342
R15974 VSS.n682 VSS.n686 0.0721009
R15975 VSS.n687 VSS.n683 4.5005
R15976 VSS.n688 VSS.n684 4.5005
R15977 VSS.n689 VSS.n685 4.5005
R15978 VSS.n675 VSS.n686 4.57442
R15979 VSS.n682 VSS.n683 0.147342
R15980 VSS.n683 VSS.n684 0.147342
R15981 VSS.n684 VSS.n685 0.147342
R15982 VSS.n686 VSS.n687 2.39784
R15983 VSS.n687 VSS.n688 0.147342
R15984 VSS.n688 VSS.n689 0.147342
R15985 VSS.n689 VSS.t582 3.13212
R15986 VSS.n662 VSS.n667 4.5005
R15987 VSS.n664 VSS.n668 4.5005
R15988 VSS.n665 VSS.n669 4.5005
R15989 VSS.n666 VSS.n670 4.57324
R15990 VSS.n662 VSS.n660 0.147342
R15991 VSS.n663 VSS.n664 0.0732424
R15992 VSS.n664 VSS.n665 0.147342
R15993 VSS.n667 VSS.n671 0.0721009
R15994 VSS.n672 VSS.n668 4.5005
R15995 VSS.n673 VSS.n669 4.5005
R15996 VSS.n674 VSS.n670 4.5005
R15997 VSS.n660 VSS.n671 4.57442
R15998 VSS.n667 VSS.n668 0.147342
R15999 VSS.n668 VSS.n669 0.147342
R16000 VSS.n669 VSS.n670 0.147342
R16001 VSS.n671 VSS.n672 2.39784
R16002 VSS.n672 VSS.n673 0.147342
R16003 VSS.n673 VSS.n674 0.147342
R16004 VSS.n674 VSS.t404 3.13212
R16005 VSS.n647 VSS.n652 4.5005
R16006 VSS.n649 VSS.n653 4.5005
R16007 VSS.n650 VSS.n654 4.5005
R16008 VSS.n651 VSS.n655 4.57324
R16009 VSS.n647 VSS.n645 0.147342
R16010 VSS.n648 VSS.n649 0.0732424
R16011 VSS.n649 VSS.n650 0.147342
R16012 VSS.n652 VSS.n656 0.0721009
R16013 VSS.n657 VSS.n653 4.5005
R16014 VSS.n658 VSS.n654 4.5005
R16015 VSS.n659 VSS.n655 4.5005
R16016 VSS.n645 VSS.n656 4.57442
R16017 VSS.n652 VSS.n653 0.147342
R16018 VSS.n653 VSS.n654 0.147342
R16019 VSS.n654 VSS.n655 0.147342
R16020 VSS.n656 VSS.n657 2.39784
R16021 VSS.n657 VSS.n658 0.147342
R16022 VSS.n658 VSS.n659 0.147342
R16023 VSS.n659 VSS.t504 3.13212
R16024 VSS.n632 VSS.n637 4.5005
R16025 VSS.n634 VSS.n638 4.5005
R16026 VSS.n635 VSS.n639 4.5005
R16027 VSS.n636 VSS.n640 4.57324
R16028 VSS.n632 VSS.n630 0.147342
R16029 VSS.n633 VSS.n634 0.0732424
R16030 VSS.n634 VSS.n635 0.147342
R16031 VSS.n637 VSS.n641 0.0721009
R16032 VSS.n642 VSS.n638 4.5005
R16033 VSS.n643 VSS.n639 4.5005
R16034 VSS.n644 VSS.n640 4.5005
R16035 VSS.n630 VSS.n641 4.57442
R16036 VSS.n637 VSS.n638 0.147342
R16037 VSS.n638 VSS.n639 0.147342
R16038 VSS.n639 VSS.n640 0.147342
R16039 VSS.n641 VSS.n642 2.39784
R16040 VSS.n642 VSS.n643 0.147342
R16041 VSS.n643 VSS.n644 0.147342
R16042 VSS.n644 VSS.t21 3.13212
R16043 VSS.n617 VSS.n622 4.5005
R16044 VSS.n619 VSS.n623 4.5005
R16045 VSS.n620 VSS.n624 4.5005
R16046 VSS.n621 VSS.n625 4.57324
R16047 VSS.n617 VSS.n615 0.147342
R16048 VSS.n618 VSS.n619 0.0732424
R16049 VSS.n619 VSS.n620 0.147342
R16050 VSS.n622 VSS.n626 0.0721009
R16051 VSS.n627 VSS.n623 4.5005
R16052 VSS.n628 VSS.n624 4.5005
R16053 VSS.n629 VSS.n625 4.5005
R16054 VSS.n615 VSS.n626 4.57442
R16055 VSS.n622 VSS.n623 0.147342
R16056 VSS.n623 VSS.n624 0.147342
R16057 VSS.n624 VSS.n625 0.147342
R16058 VSS.n626 VSS.n627 2.39784
R16059 VSS.n627 VSS.n628 0.147342
R16060 VSS.n628 VSS.n629 0.147342
R16061 VSS.n629 VSS.t397 3.13212
R16062 VSS.n596 VSS.n601 4.5005
R16063 VSS.n598 VSS.n602 4.5005
R16064 VSS.n599 VSS.n603 4.5005
R16065 VSS.n600 VSS.n604 4.57324
R16066 VSS.n596 VSS.n594 0.147342
R16067 VSS.n597 VSS.n598 0.0732424
R16068 VSS.n598 VSS.n599 0.147342
R16069 VSS.n601 VSS.n605 0.0721009
R16070 VSS.n606 VSS.n602 4.5005
R16071 VSS.n607 VSS.n603 4.5005
R16072 VSS.n608 VSS.n604 4.5005
R16073 VSS.n594 VSS.n605 4.57442
R16074 VSS.n601 VSS.n602 0.147342
R16075 VSS.n602 VSS.n603 0.147342
R16076 VSS.n603 VSS.n604 0.147342
R16077 VSS.n605 VSS.n606 2.39784
R16078 VSS.n606 VSS.n607 0.147342
R16079 VSS.n607 VSS.n608 0.147342
R16080 VSS.n608 VSS.t359 3.13212
R16081 VSS.n581 VSS.n586 4.5005
R16082 VSS.n583 VSS.n587 4.5005
R16083 VSS.n584 VSS.n588 4.5005
R16084 VSS.n585 VSS.n589 4.57324
R16085 VSS.n581 VSS.n579 0.147342
R16086 VSS.n582 VSS.n583 0.0732424
R16087 VSS.n583 VSS.n584 0.147342
R16088 VSS.n586 VSS.n590 0.0721009
R16089 VSS.n591 VSS.n587 4.5005
R16090 VSS.n592 VSS.n588 4.5005
R16091 VSS.n593 VSS.n589 4.5005
R16092 VSS.n579 VSS.n590 4.57442
R16093 VSS.n586 VSS.n587 0.147342
R16094 VSS.n587 VSS.n588 0.147342
R16095 VSS.n588 VSS.n589 0.147342
R16096 VSS.n590 VSS.n591 2.39784
R16097 VSS.n591 VSS.n592 0.147342
R16098 VSS.n592 VSS.n593 0.147342
R16099 VSS.n593 VSS.t336 3.13212
R16100 VSS.n566 VSS.n571 4.5005
R16101 VSS.n568 VSS.n572 4.5005
R16102 VSS.n569 VSS.n573 4.5005
R16103 VSS.n570 VSS.n574 4.57324
R16104 VSS.n566 VSS.n564 0.147342
R16105 VSS.n567 VSS.n568 0.0732424
R16106 VSS.n568 VSS.n569 0.147342
R16107 VSS.n571 VSS.n575 0.0721009
R16108 VSS.n576 VSS.n572 4.5005
R16109 VSS.n577 VSS.n573 4.5005
R16110 VSS.n578 VSS.n574 4.5005
R16111 VSS.n564 VSS.n575 4.57442
R16112 VSS.n571 VSS.n572 0.147342
R16113 VSS.n572 VSS.n573 0.147342
R16114 VSS.n573 VSS.n574 0.147342
R16115 VSS.n575 VSS.n576 2.39784
R16116 VSS.n576 VSS.n577 0.147342
R16117 VSS.n577 VSS.n578 0.147342
R16118 VSS.n578 VSS.t322 3.13212
R16119 VSS.n545 VSS.n550 4.5005
R16120 VSS.n547 VSS.n551 4.5005
R16121 VSS.n548 VSS.n552 4.5005
R16122 VSS.n549 VSS.n553 4.57324
R16123 VSS.n545 VSS.n543 0.147342
R16124 VSS.n546 VSS.n547 0.0732424
R16125 VSS.n547 VSS.n548 0.147342
R16126 VSS.n550 VSS.n554 0.0721009
R16127 VSS.n555 VSS.n551 4.5005
R16128 VSS.n556 VSS.n552 4.5005
R16129 VSS.n557 VSS.n553 4.5005
R16130 VSS.n543 VSS.n554 4.57442
R16131 VSS.n550 VSS.n551 0.147342
R16132 VSS.n551 VSS.n552 0.147342
R16133 VSS.n552 VSS.n553 0.147342
R16134 VSS.n554 VSS.n555 2.39784
R16135 VSS.n555 VSS.n556 0.147342
R16136 VSS.n556 VSS.n557 0.147342
R16137 VSS.n557 VSS.t385 3.13212
R16138 VSS.n530 VSS.n535 4.5005
R16139 VSS.n532 VSS.n536 4.5005
R16140 VSS.n533 VSS.n537 4.5005
R16141 VSS.n534 VSS.n538 4.57324
R16142 VSS.n530 VSS.n528 0.147342
R16143 VSS.n531 VSS.n532 0.0732424
R16144 VSS.n532 VSS.n533 0.147342
R16145 VSS.n535 VSS.n539 0.0721009
R16146 VSS.n540 VSS.n536 4.5005
R16147 VSS.n541 VSS.n537 4.5005
R16148 VSS.n542 VSS.n538 4.5005
R16149 VSS.n528 VSS.n539 4.57442
R16150 VSS.n535 VSS.n536 0.147342
R16151 VSS.n536 VSS.n537 0.147342
R16152 VSS.n537 VSS.n538 0.147342
R16153 VSS.n539 VSS.n540 2.39784
R16154 VSS.n540 VSS.n541 0.147342
R16155 VSS.n541 VSS.n542 0.147342
R16156 VSS.n542 VSS.t459 3.13212
R16157 VSS.n515 VSS.n520 4.5005
R16158 VSS.n517 VSS.n521 4.5005
R16159 VSS.n518 VSS.n522 4.5005
R16160 VSS.n519 VSS.n523 4.57324
R16161 VSS.n515 VSS.n513 0.147342
R16162 VSS.n516 VSS.n517 0.0732424
R16163 VSS.n517 VSS.n518 0.147342
R16164 VSS.n520 VSS.n524 0.0721009
R16165 VSS.n525 VSS.n521 4.5005
R16166 VSS.n526 VSS.n522 4.5005
R16167 VSS.n527 VSS.n523 4.5005
R16168 VSS.n513 VSS.n524 4.57442
R16169 VSS.n520 VSS.n521 0.147342
R16170 VSS.n521 VSS.n522 0.147342
R16171 VSS.n522 VSS.n523 0.147342
R16172 VSS.n524 VSS.n525 2.39784
R16173 VSS.n525 VSS.n526 0.147342
R16174 VSS.n526 VSS.n527 0.147342
R16175 VSS.n527 VSS.t227 3.13212
R16176 VSS.n500 VSS.n505 4.5005
R16177 VSS.n502 VSS.n506 4.5005
R16178 VSS.n503 VSS.n507 4.5005
R16179 VSS.n504 VSS.n508 4.57324
R16180 VSS.n500 VSS.n498 0.147342
R16181 VSS.n501 VSS.n502 0.0732424
R16182 VSS.n502 VSS.n503 0.147342
R16183 VSS.n505 VSS.n509 0.0721009
R16184 VSS.n510 VSS.n506 4.5005
R16185 VSS.n511 VSS.n507 4.5005
R16186 VSS.n512 VSS.n508 4.5005
R16187 VSS.n498 VSS.n509 4.57442
R16188 VSS.n505 VSS.n506 0.147342
R16189 VSS.n506 VSS.n507 0.147342
R16190 VSS.n507 VSS.n508 0.147342
R16191 VSS.n509 VSS.n510 2.39784
R16192 VSS.n510 VSS.n511 0.147342
R16193 VSS.n511 VSS.n512 0.147342
R16194 VSS.n512 VSS.t305 3.13212
R16195 VSS.n479 VSS.n484 4.5005
R16196 VSS.n481 VSS.n485 4.5005
R16197 VSS.n482 VSS.n486 4.5005
R16198 VSS.n483 VSS.n487 4.57324
R16199 VSS.n479 VSS.n477 0.147342
R16200 VSS.n480 VSS.n481 0.0732424
R16201 VSS.n481 VSS.n482 0.147342
R16202 VSS.n484 VSS.n488 0.0721009
R16203 VSS.n489 VSS.n485 4.5005
R16204 VSS.n490 VSS.n486 4.5005
R16205 VSS.n491 VSS.n487 4.5005
R16206 VSS.n477 VSS.n488 4.57442
R16207 VSS.n484 VSS.n485 0.147342
R16208 VSS.n485 VSS.n486 0.147342
R16209 VSS.n486 VSS.n487 0.147342
R16210 VSS.n488 VSS.n489 2.39784
R16211 VSS.n489 VSS.n490 0.147342
R16212 VSS.n490 VSS.n491 0.147342
R16213 VSS.n491 VSS.t560 3.13212
R16214 VSS.n464 VSS.n469 4.5005
R16215 VSS.n466 VSS.n470 4.5005
R16216 VSS.n467 VSS.n471 4.5005
R16217 VSS.n468 VSS.n472 4.57324
R16218 VSS.n464 VSS.n462 0.147342
R16219 VSS.n465 VSS.n466 0.0732424
R16220 VSS.n466 VSS.n467 0.147342
R16221 VSS.n469 VSS.n473 0.0721009
R16222 VSS.n474 VSS.n470 4.5005
R16223 VSS.n475 VSS.n471 4.5005
R16224 VSS.n476 VSS.n472 4.5005
R16225 VSS.n462 VSS.n473 4.57442
R16226 VSS.n469 VSS.n470 0.147342
R16227 VSS.n470 VSS.n471 0.147342
R16228 VSS.n471 VSS.n472 0.147342
R16229 VSS.n473 VSS.n474 2.39784
R16230 VSS.n474 VSS.n475 0.147342
R16231 VSS.n475 VSS.n476 0.147342
R16232 VSS.n476 VSS.t375 3.13212
R16233 VSS.n449 VSS.n454 4.5005
R16234 VSS.n451 VSS.n455 4.5005
R16235 VSS.n452 VSS.n456 4.5005
R16236 VSS.n453 VSS.n457 4.57324
R16237 VSS.n449 VSS.n447 0.147342
R16238 VSS.n450 VSS.n451 0.0732424
R16239 VSS.n451 VSS.n452 0.147342
R16240 VSS.n454 VSS.n458 0.0721009
R16241 VSS.n459 VSS.n455 4.5005
R16242 VSS.n460 VSS.n456 4.5005
R16243 VSS.n461 VSS.n457 4.5005
R16244 VSS.n447 VSS.n458 4.57442
R16245 VSS.n454 VSS.n455 0.147342
R16246 VSS.n455 VSS.n456 0.147342
R16247 VSS.n456 VSS.n457 0.147342
R16248 VSS.n458 VSS.n459 2.39784
R16249 VSS.n459 VSS.n460 0.147342
R16250 VSS.n460 VSS.n461 0.147342
R16251 VSS.n461 VSS.t269 3.13212
R16252 VSS.n428 VSS.n433 4.5005
R16253 VSS.n430 VSS.n434 4.5005
R16254 VSS.n431 VSS.n435 4.5005
R16255 VSS.n432 VSS.n436 4.57324
R16256 VSS.n428 VSS.n426 0.147342
R16257 VSS.n429 VSS.n430 0.0732424
R16258 VSS.n430 VSS.n431 0.147342
R16259 VSS.n433 VSS.n437 0.0721009
R16260 VSS.n438 VSS.n434 4.5005
R16261 VSS.n439 VSS.n435 4.5005
R16262 VSS.n440 VSS.n436 4.5005
R16263 VSS.n426 VSS.n437 4.57442
R16264 VSS.n433 VSS.n434 0.147342
R16265 VSS.n434 VSS.n435 0.147342
R16266 VSS.n435 VSS.n436 0.147342
R16267 VSS.n437 VSS.n438 2.39784
R16268 VSS.n438 VSS.n439 0.147342
R16269 VSS.n439 VSS.n440 0.147342
R16270 VSS.n440 VSS.t288 3.13212
R16271 VSS.n413 VSS.n418 4.5005
R16272 VSS.n415 VSS.n419 4.5005
R16273 VSS.n416 VSS.n420 4.5005
R16274 VSS.n417 VSS.n421 4.57324
R16275 VSS.n413 VSS.n411 0.147342
R16276 VSS.n414 VSS.n415 0.0732424
R16277 VSS.n415 VSS.n416 0.147342
R16278 VSS.n418 VSS.n422 0.0721009
R16279 VSS.n423 VSS.n419 4.5005
R16280 VSS.n424 VSS.n420 4.5005
R16281 VSS.n425 VSS.n421 4.5005
R16282 VSS.n411 VSS.n422 4.57442
R16283 VSS.n418 VSS.n419 0.147342
R16284 VSS.n419 VSS.n420 0.147342
R16285 VSS.n420 VSS.n421 0.147342
R16286 VSS.n422 VSS.n423 2.39784
R16287 VSS.n423 VSS.n424 0.147342
R16288 VSS.n424 VSS.n425 0.147342
R16289 VSS.n425 VSS.t583 3.13212
R16290 VSS.n398 VSS.n403 4.5005
R16291 VSS.n400 VSS.n404 4.5005
R16292 VSS.n401 VSS.n405 4.5005
R16293 VSS.n402 VSS.n406 4.57324
R16294 VSS.n398 VSS.n396 0.147342
R16295 VSS.n399 VSS.n400 0.0732424
R16296 VSS.n400 VSS.n401 0.147342
R16297 VSS.n403 VSS.n407 0.0721009
R16298 VSS.n408 VSS.n404 4.5005
R16299 VSS.n409 VSS.n405 4.5005
R16300 VSS.n410 VSS.n406 4.5005
R16301 VSS.n396 VSS.n407 4.57442
R16302 VSS.n403 VSS.n404 0.147342
R16303 VSS.n404 VSS.n405 0.147342
R16304 VSS.n405 VSS.n406 0.147342
R16305 VSS.n407 VSS.n408 2.39784
R16306 VSS.n408 VSS.n409 0.147342
R16307 VSS.n409 VSS.n410 0.147342
R16308 VSS.n410 VSS.t425 3.13212
R16309 VSS.n383 VSS.n388 4.5005
R16310 VSS.n385 VSS.n389 4.5005
R16311 VSS.n386 VSS.n390 4.5005
R16312 VSS.n387 VSS.n391 4.57324
R16313 VSS.n383 VSS.n381 0.147342
R16314 VSS.n384 VSS.n385 0.0732424
R16315 VSS.n385 VSS.n386 0.147342
R16316 VSS.n388 VSS.n392 0.0721009
R16317 VSS.n393 VSS.n389 4.5005
R16318 VSS.n394 VSS.n390 4.5005
R16319 VSS.n395 VSS.n391 4.5005
R16320 VSS.n381 VSS.n392 4.57442
R16321 VSS.n388 VSS.n389 0.147342
R16322 VSS.n389 VSS.n390 0.147342
R16323 VSS.n390 VSS.n391 0.147342
R16324 VSS.n392 VSS.n393 2.39784
R16325 VSS.n393 VSS.n394 0.147342
R16326 VSS.n394 VSS.n395 0.147342
R16327 VSS.n395 VSS.t502 3.13212
R16328 VSS.n368 VSS.n373 4.5005
R16329 VSS.n370 VSS.n374 4.5005
R16330 VSS.n371 VSS.n375 4.5005
R16331 VSS.n372 VSS.n376 4.57324
R16332 VSS.n368 VSS.n366 0.147342
R16333 VSS.n369 VSS.n370 0.0732424
R16334 VSS.n370 VSS.n371 0.147342
R16335 VSS.n373 VSS.n377 0.0721009
R16336 VSS.n378 VSS.n374 4.5005
R16337 VSS.n379 VSS.n375 4.5005
R16338 VSS.n380 VSS.n376 4.5005
R16339 VSS.n366 VSS.n377 4.57442
R16340 VSS.n373 VSS.n374 0.147342
R16341 VSS.n374 VSS.n375 0.147342
R16342 VSS.n375 VSS.n376 0.147342
R16343 VSS.n377 VSS.n378 2.39784
R16344 VSS.n378 VSS.n379 0.147342
R16345 VSS.n379 VSS.n380 0.147342
R16346 VSS.n380 VSS.t27 3.13212
R16347 VSS.n353 VSS.n358 4.5005
R16348 VSS.n355 VSS.n359 4.5005
R16349 VSS.n356 VSS.n360 4.5005
R16350 VSS.n357 VSS.n361 4.57324
R16351 VSS.n353 VSS.n351 0.147342
R16352 VSS.n354 VSS.n355 0.0732424
R16353 VSS.n355 VSS.n356 0.147342
R16354 VSS.n358 VSS.n362 0.0721009
R16355 VSS.n363 VSS.n359 4.5005
R16356 VSS.n364 VSS.n360 4.5005
R16357 VSS.n365 VSS.n361 4.5005
R16358 VSS.n351 VSS.n362 4.57442
R16359 VSS.n358 VSS.n359 0.147342
R16360 VSS.n359 VSS.n360 0.147342
R16361 VSS.n360 VSS.n361 0.147342
R16362 VSS.n362 VSS.n363 2.39784
R16363 VSS.n363 VSS.n364 0.147342
R16364 VSS.n364 VSS.n365 0.147342
R16365 VSS.n365 VSS.t352 3.13212
R16366 VSS.n332 VSS.n337 4.5005
R16367 VSS.n334 VSS.n338 4.5005
R16368 VSS.n335 VSS.n339 4.5005
R16369 VSS.n336 VSS.n340 4.57324
R16370 VSS.n332 VSS.n330 0.147342
R16371 VSS.n333 VSS.n334 0.0732424
R16372 VSS.n334 VSS.n335 0.147342
R16373 VSS.n337 VSS.n341 0.0721009
R16374 VSS.n342 VSS.n338 4.5005
R16375 VSS.n343 VSS.n339 4.5005
R16376 VSS.n344 VSS.n340 4.5005
R16377 VSS.n330 VSS.n341 4.57442
R16378 VSS.n337 VSS.n338 0.147342
R16379 VSS.n338 VSS.n339 0.147342
R16380 VSS.n339 VSS.n340 0.147342
R16381 VSS.n341 VSS.n342 2.39784
R16382 VSS.n342 VSS.n343 0.147342
R16383 VSS.n343 VSS.n344 0.147342
R16384 VSS.n344 VSS.t314 3.13212
R16385 VSS.n317 VSS.n322 4.5005
R16386 VSS.n319 VSS.n323 4.5005
R16387 VSS.n320 VSS.n324 4.5005
R16388 VSS.n321 VSS.n325 4.57324
R16389 VSS.n317 VSS.n315 0.147342
R16390 VSS.n318 VSS.n319 0.0732424
R16391 VSS.n319 VSS.n320 0.147342
R16392 VSS.n322 VSS.n326 0.0721009
R16393 VSS.n327 VSS.n323 4.5005
R16394 VSS.n328 VSS.n324 4.5005
R16395 VSS.n329 VSS.n325 4.5005
R16396 VSS.n315 VSS.n326 4.57442
R16397 VSS.n322 VSS.n323 0.147342
R16398 VSS.n323 VSS.n324 0.147342
R16399 VSS.n324 VSS.n325 0.147342
R16400 VSS.n326 VSS.n327 2.39784
R16401 VSS.n327 VSS.n328 0.147342
R16402 VSS.n328 VSS.n329 0.147342
R16403 VSS.n329 VSS.t339 3.13212
R16404 VSS.n302 VSS.n307 4.5005
R16405 VSS.n304 VSS.n308 4.5005
R16406 VSS.n305 VSS.n309 4.5005
R16407 VSS.n306 VSS.n310 4.57324
R16408 VSS.n302 VSS.n300 0.147342
R16409 VSS.n303 VSS.n304 0.0732424
R16410 VSS.n304 VSS.n305 0.147342
R16411 VSS.n307 VSS.n311 0.0721009
R16412 VSS.n312 VSS.n308 4.5005
R16413 VSS.n313 VSS.n309 4.5005
R16414 VSS.n314 VSS.n310 4.5005
R16415 VSS.n300 VSS.n311 4.57442
R16416 VSS.n307 VSS.n308 0.147342
R16417 VSS.n308 VSS.n309 0.147342
R16418 VSS.n309 VSS.n310 0.147342
R16419 VSS.n311 VSS.n312 2.39784
R16420 VSS.n312 VSS.n313 0.147342
R16421 VSS.n313 VSS.n314 0.147342
R16422 VSS.n314 VSS.t324 3.13212
R16423 VSS.n281 VSS.n286 4.5005
R16424 VSS.n283 VSS.n287 4.5005
R16425 VSS.n284 VSS.n288 4.5005
R16426 VSS.n285 VSS.n289 4.57324
R16427 VSS.n281 VSS.n279 0.147342
R16428 VSS.n282 VSS.n283 0.0732424
R16429 VSS.n283 VSS.n284 0.147342
R16430 VSS.n286 VSS.n290 0.0721009
R16431 VSS.n291 VSS.n287 4.5005
R16432 VSS.n292 VSS.n288 4.5005
R16433 VSS.n293 VSS.n289 4.5005
R16434 VSS.n279 VSS.n290 4.57442
R16435 VSS.n286 VSS.n287 0.147342
R16436 VSS.n287 VSS.n288 0.147342
R16437 VSS.n288 VSS.n289 0.147342
R16438 VSS.n290 VSS.n291 2.39784
R16439 VSS.n291 VSS.n292 0.147342
R16440 VSS.n292 VSS.n293 0.147342
R16441 VSS.n293 VSS.t383 3.13212
R16442 VSS.n266 VSS.n271 4.5005
R16443 VSS.n268 VSS.n272 4.5005
R16444 VSS.n269 VSS.n273 4.5005
R16445 VSS.n270 VSS.n274 4.57324
R16446 VSS.n266 VSS.n264 0.147342
R16447 VSS.n267 VSS.n268 0.0732424
R16448 VSS.n268 VSS.n269 0.147342
R16449 VSS.n271 VSS.n275 0.0721009
R16450 VSS.n276 VSS.n272 4.5005
R16451 VSS.n277 VSS.n273 4.5005
R16452 VSS.n278 VSS.n274 4.5005
R16453 VSS.n264 VSS.n275 4.57442
R16454 VSS.n271 VSS.n272 0.147342
R16455 VSS.n272 VSS.n273 0.147342
R16456 VSS.n273 VSS.n274 0.147342
R16457 VSS.n275 VSS.n276 2.39784
R16458 VSS.n276 VSS.n277 0.147342
R16459 VSS.n277 VSS.n278 0.147342
R16460 VSS.n278 VSS.t175 3.13212
R16461 VSS.n251 VSS.n256 4.5005
R16462 VSS.n253 VSS.n257 4.5005
R16463 VSS.n254 VSS.n258 4.5005
R16464 VSS.n255 VSS.n259 4.57324
R16465 VSS.n251 VSS.n249 0.147342
R16466 VSS.n252 VSS.n253 0.0732424
R16467 VSS.n253 VSS.n254 0.147342
R16468 VSS.n256 VSS.n260 0.0721009
R16469 VSS.n261 VSS.n257 4.5005
R16470 VSS.n262 VSS.n258 4.5005
R16471 VSS.n263 VSS.n259 4.5005
R16472 VSS.n249 VSS.n260 4.57442
R16473 VSS.n256 VSS.n257 0.147342
R16474 VSS.n257 VSS.n258 0.147342
R16475 VSS.n258 VSS.n259 0.147342
R16476 VSS.n260 VSS.n261 2.39784
R16477 VSS.n261 VSS.n262 0.147342
R16478 VSS.n262 VSS.n263 0.147342
R16479 VSS.n263 VSS.t220 3.13212
R16480 VSS.n236 VSS.n241 4.5005
R16481 VSS.n238 VSS.n242 4.5005
R16482 VSS.n239 VSS.n243 4.5005
R16483 VSS.n240 VSS.n244 4.57324
R16484 VSS.n236 VSS.n234 0.147342
R16485 VSS.n237 VSS.n238 0.0732424
R16486 VSS.n238 VSS.n239 0.147342
R16487 VSS.n241 VSS.n245 0.0721009
R16488 VSS.n246 VSS.n242 4.5005
R16489 VSS.n247 VSS.n243 4.5005
R16490 VSS.n248 VSS.n244 4.5005
R16491 VSS.n234 VSS.n245 4.57442
R16492 VSS.n241 VSS.n242 0.147342
R16493 VSS.n242 VSS.n243 0.147342
R16494 VSS.n243 VSS.n244 0.147342
R16495 VSS.n245 VSS.n246 2.39784
R16496 VSS.n246 VSS.n247 0.147342
R16497 VSS.n247 VSS.n248 0.147342
R16498 VSS.n248 VSS.t290 3.13212
R16499 VSS.n215 VSS.n220 4.5005
R16500 VSS.n217 VSS.n221 4.5005
R16501 VSS.n218 VSS.n222 4.5005
R16502 VSS.n219 VSS.n223 4.57324
R16503 VSS.n215 VSS.n213 0.147342
R16504 VSS.n216 VSS.n217 0.0732424
R16505 VSS.n217 VSS.n218 0.147342
R16506 VSS.n220 VSS.n224 0.0721009
R16507 VSS.n225 VSS.n221 4.5005
R16508 VSS.n226 VSS.n222 4.5005
R16509 VSS.n227 VSS.n223 4.5005
R16510 VSS.n213 VSS.n224 4.57442
R16511 VSS.n220 VSS.n221 0.147342
R16512 VSS.n221 VSS.n222 0.147342
R16513 VSS.n222 VSS.n223 0.147342
R16514 VSS.n224 VSS.n225 2.39784
R16515 VSS.n225 VSS.n226 0.147342
R16516 VSS.n226 VSS.n227 0.147342
R16517 VSS.n227 VSS.t564 3.13212
R16518 VSS.n200 VSS.n205 4.5005
R16519 VSS.n202 VSS.n206 4.5005
R16520 VSS.n203 VSS.n207 4.5005
R16521 VSS.n204 VSS.n208 4.57324
R16522 VSS.n200 VSS.n198 0.147342
R16523 VSS.n201 VSS.n202 0.0732424
R16524 VSS.n202 VSS.n203 0.147342
R16525 VSS.n205 VSS.n209 0.0721009
R16526 VSS.n210 VSS.n206 4.5005
R16527 VSS.n211 VSS.n207 4.5005
R16528 VSS.n212 VSS.n208 4.5005
R16529 VSS.n198 VSS.n209 4.57442
R16530 VSS.n205 VSS.n206 0.147342
R16531 VSS.n206 VSS.n207 0.147342
R16532 VSS.n207 VSS.n208 0.147342
R16533 VSS.n209 VSS.n210 2.39784
R16534 VSS.n210 VSS.n211 0.147342
R16535 VSS.n211 VSS.n212 0.147342
R16536 VSS.n212 VSS.t378 3.13212
R16537 VSS.n185 VSS.n190 4.5005
R16538 VSS.n187 VSS.n191 4.5005
R16539 VSS.n188 VSS.n192 4.5005
R16540 VSS.n189 VSS.n193 4.57324
R16541 VSS.n185 VSS.n183 0.147342
R16542 VSS.n186 VSS.n187 0.0732424
R16543 VSS.n187 VSS.n188 0.147342
R16544 VSS.n190 VSS.n194 0.0721009
R16545 VSS.n195 VSS.n191 4.5005
R16546 VSS.n196 VSS.n192 4.5005
R16547 VSS.n197 VSS.n193 4.5005
R16548 VSS.n183 VSS.n194 4.57442
R16549 VSS.n190 VSS.n191 0.147342
R16550 VSS.n191 VSS.n192 0.147342
R16551 VSS.n192 VSS.n193 0.147342
R16552 VSS.n194 VSS.n195 2.39784
R16553 VSS.n195 VSS.n196 0.147342
R16554 VSS.n196 VSS.n197 0.147342
R16555 VSS.n197 VSS.t595 3.13212
R16556 VSS.n164 VSS.n169 4.5005
R16557 VSS.n166 VSS.n170 4.5005
R16558 VSS.n167 VSS.n171 4.5005
R16559 VSS.n168 VSS.n172 4.57324
R16560 VSS.n164 VSS.n162 0.147342
R16561 VSS.n165 VSS.n166 0.0732424
R16562 VSS.n166 VSS.n167 0.147342
R16563 VSS.n169 VSS.n173 0.0721009
R16564 VSS.n174 VSS.n170 4.5005
R16565 VSS.n175 VSS.n171 4.5005
R16566 VSS.n176 VSS.n172 4.5005
R16567 VSS.n162 VSS.n173 4.57442
R16568 VSS.n169 VSS.n170 0.147342
R16569 VSS.n170 VSS.n171 0.147342
R16570 VSS.n171 VSS.n172 0.147342
R16571 VSS.n173 VSS.n174 2.39784
R16572 VSS.n174 VSS.n175 0.147342
R16573 VSS.n175 VSS.n176 0.147342
R16574 VSS.n176 VSS.t366 3.13212
R16575 VSS.n149 VSS.n154 4.5005
R16576 VSS.n151 VSS.n155 4.5005
R16577 VSS.n152 VSS.n156 4.5005
R16578 VSS.n153 VSS.n157 4.57324
R16579 VSS.n149 VSS.n147 0.147342
R16580 VSS.n150 VSS.n151 0.0732424
R16581 VSS.n151 VSS.n152 0.147342
R16582 VSS.n154 VSS.n158 0.0721009
R16583 VSS.n159 VSS.n155 4.5005
R16584 VSS.n160 VSS.n156 4.5005
R16585 VSS.n161 VSS.n157 4.5005
R16586 VSS.n147 VSS.n158 4.57442
R16587 VSS.n154 VSS.n155 0.147342
R16588 VSS.n155 VSS.n156 0.147342
R16589 VSS.n156 VSS.n157 0.147342
R16590 VSS.n158 VSS.n159 2.39784
R16591 VSS.n159 VSS.n160 0.147342
R16592 VSS.n160 VSS.n161 0.147342
R16593 VSS.n161 VSS.t584 3.13212
R16594 VSS.n134 VSS.n139 4.5005
R16595 VSS.n136 VSS.n140 4.5005
R16596 VSS.n137 VSS.n141 4.5005
R16597 VSS.n138 VSS.n142 4.57324
R16598 VSS.n134 VSS.n132 0.147342
R16599 VSS.n135 VSS.n136 0.0732424
R16600 VSS.n136 VSS.n137 0.147342
R16601 VSS.n139 VSS.n143 0.0721009
R16602 VSS.n144 VSS.n140 4.5005
R16603 VSS.n145 VSS.n141 4.5005
R16604 VSS.n146 VSS.n142 4.5005
R16605 VSS.n132 VSS.n143 4.57442
R16606 VSS.n139 VSS.n140 0.147342
R16607 VSS.n140 VSS.n141 0.147342
R16608 VSS.n141 VSS.n142 0.147342
R16609 VSS.n143 VSS.n144 2.39784
R16610 VSS.n144 VSS.n145 0.147342
R16611 VSS.n145 VSS.n146 0.147342
R16612 VSS.n146 VSS.t277 3.13212
R16613 VSS.n119 VSS.n124 4.5005
R16614 VSS.n121 VSS.n125 4.5005
R16615 VSS.n122 VSS.n126 4.5005
R16616 VSS.n123 VSS.n127 4.57324
R16617 VSS.n119 VSS.n117 0.147342
R16618 VSS.n120 VSS.n121 0.0732424
R16619 VSS.n121 VSS.n122 0.147342
R16620 VSS.n124 VSS.n128 0.0721009
R16621 VSS.n129 VSS.n125 4.5005
R16622 VSS.n130 VSS.n126 4.5005
R16623 VSS.n131 VSS.n127 4.5005
R16624 VSS.n117 VSS.n128 4.57442
R16625 VSS.n124 VSS.n125 0.147342
R16626 VSS.n125 VSS.n126 0.147342
R16627 VSS.n126 VSS.n127 0.147342
R16628 VSS.n128 VSS.n129 2.39784
R16629 VSS.n129 VSS.n130 0.147342
R16630 VSS.n130 VSS.n131 0.147342
R16631 VSS.n131 VSS.t82 3.13212
R16632 VSS.n104 VSS.n109 4.5005
R16633 VSS.n106 VSS.n110 4.5005
R16634 VSS.n107 VSS.n111 4.5005
R16635 VSS.n108 VSS.n112 4.57324
R16636 VSS.n104 VSS.n102 0.147342
R16637 VSS.n105 VSS.n106 0.0732424
R16638 VSS.n106 VSS.n107 0.147342
R16639 VSS.n109 VSS.n113 0.0721009
R16640 VSS.n114 VSS.n110 4.5005
R16641 VSS.n115 VSS.n111 4.5005
R16642 VSS.n116 VSS.n112 4.5005
R16643 VSS.n102 VSS.n113 4.57442
R16644 VSS.n109 VSS.n110 0.147342
R16645 VSS.n110 VSS.n111 0.147342
R16646 VSS.n111 VSS.n112 0.147342
R16647 VSS.n113 VSS.n114 2.39784
R16648 VSS.n114 VSS.n115 0.147342
R16649 VSS.n115 VSS.n116 0.147342
R16650 VSS.n116 VSS.t25 3.13212
R16651 VSS.n89 VSS.n94 4.5005
R16652 VSS.n91 VSS.n95 4.5005
R16653 VSS.n92 VSS.n96 4.5005
R16654 VSS.n93 VSS.n97 4.57324
R16655 VSS.n89 VSS.n87 0.147342
R16656 VSS.n90 VSS.n91 0.0732424
R16657 VSS.n91 VSS.n92 0.147342
R16658 VSS.n94 VSS.n98 0.0721009
R16659 VSS.n99 VSS.n95 4.5005
R16660 VSS.n100 VSS.n96 4.5005
R16661 VSS.n101 VSS.n97 4.5005
R16662 VSS.n87 VSS.n98 4.57442
R16663 VSS.n94 VSS.n95 0.147342
R16664 VSS.n95 VSS.n96 0.147342
R16665 VSS.n96 VSS.n97 0.147342
R16666 VSS.n98 VSS.n99 2.39784
R16667 VSS.n99 VSS.n100 0.147342
R16668 VSS.n100 VSS.n101 0.147342
R16669 VSS.n101 VSS.t354 3.13212
R16670 VSS.n68 VSS.n73 4.5005
R16671 VSS.n70 VSS.n74 4.5005
R16672 VSS.n71 VSS.n75 4.5005
R16673 VSS.n72 VSS.n76 4.57324
R16674 VSS.n68 VSS.n66 0.147342
R16675 VSS.n69 VSS.n70 0.0732424
R16676 VSS.n70 VSS.n71 0.147342
R16677 VSS.n73 VSS.n77 0.0721009
R16678 VSS.n78 VSS.n74 4.5005
R16679 VSS.n79 VSS.n75 4.5005
R16680 VSS.n80 VSS.n76 4.5005
R16681 VSS.n66 VSS.n77 4.57442
R16682 VSS.n73 VSS.n74 0.147342
R16683 VSS.n74 VSS.n75 0.147342
R16684 VSS.n75 VSS.n76 0.147342
R16685 VSS.n77 VSS.n78 2.39784
R16686 VSS.n78 VSS.n79 0.147342
R16687 VSS.n79 VSS.n80 0.147342
R16688 VSS.n80 VSS.t315 3.13212
R16689 VSS.n53 VSS.n58 4.5005
R16690 VSS.n55 VSS.n59 4.5005
R16691 VSS.n56 VSS.n60 4.5005
R16692 VSS.n57 VSS.n61 4.57324
R16693 VSS.n53 VSS.n51 0.147342
R16694 VSS.n54 VSS.n55 0.0732424
R16695 VSS.n55 VSS.n56 0.147342
R16696 VSS.n58 VSS.n62 0.0721009
R16697 VSS.n63 VSS.n59 4.5005
R16698 VSS.n64 VSS.n60 4.5005
R16699 VSS.n65 VSS.n61 4.5005
R16700 VSS.n51 VSS.n62 4.57442
R16701 VSS.n58 VSS.n59 0.147342
R16702 VSS.n59 VSS.n60 0.147342
R16703 VSS.n60 VSS.n61 0.147342
R16704 VSS.n62 VSS.n63 2.39784
R16705 VSS.n63 VSS.n64 0.147342
R16706 VSS.n64 VSS.n65 0.147342
R16707 VSS.n65 VSS.t337 3.13212
R16708 VSS.n38 VSS.n43 4.5005
R16709 VSS.n40 VSS.n44 4.5005
R16710 VSS.n41 VSS.n45 4.5005
R16711 VSS.n42 VSS.n46 4.57324
R16712 VSS.n38 VSS.n36 0.147342
R16713 VSS.n39 VSS.n40 0.0732424
R16714 VSS.n40 VSS.n41 0.147342
R16715 VSS.n43 VSS.n47 0.0721009
R16716 VSS.n48 VSS.n44 4.5005
R16717 VSS.n49 VSS.n45 4.5005
R16718 VSS.n50 VSS.n46 4.5005
R16719 VSS.n36 VSS.n47 4.57442
R16720 VSS.n43 VSS.n44 0.147342
R16721 VSS.n44 VSS.n45 0.147342
R16722 VSS.n45 VSS.n46 0.147342
R16723 VSS.n47 VSS.n48 2.39784
R16724 VSS.n48 VSS.n49 0.147342
R16725 VSS.n49 VSS.n50 0.147342
R16726 VSS.n50 VSS.t391 3.13212
R16727 VSS.n17 VSS.n22 4.5005
R16728 VSS.n19 VSS.n23 4.5005
R16729 VSS.n20 VSS.n24 4.5005
R16730 VSS.n21 VSS.n25 4.57324
R16731 VSS.n17 VSS.n15 0.147342
R16732 VSS.n18 VSS.n19 0.0732424
R16733 VSS.n19 VSS.n20 0.147342
R16734 VSS.n22 VSS.n26 0.0721009
R16735 VSS.n27 VSS.n23 4.5005
R16736 VSS.n28 VSS.n24 4.5005
R16737 VSS.n29 VSS.n25 4.5005
R16738 VSS.n15 VSS.n26 4.57442
R16739 VSS.n22 VSS.n23 0.147342
R16740 VSS.n23 VSS.n24 0.147342
R16741 VSS.n24 VSS.n25 0.147342
R16742 VSS.n26 VSS.n27 2.39784
R16743 VSS.n27 VSS.n28 0.147342
R16744 VSS.n28 VSS.n29 0.147342
R16745 VSS.n29 VSS.t386 3.13212
R16746 VSS.n2 VSS.n7 4.5005
R16747 VSS.n4 VSS.n8 4.5005
R16748 VSS.n5 VSS.n9 4.5005
R16749 VSS.n6 VSS.n10 4.57324
R16750 VSS.n2 VSS.n0 0.147342
R16751 VSS.n3 VSS.n4 0.0732424
R16752 VSS.n4 VSS.n5 0.147342
R16753 VSS.n7 VSS.n11 0.0721009
R16754 VSS.n12 VSS.n8 4.5005
R16755 VSS.n13 VSS.n9 4.5005
R16756 VSS.n14 VSS.n10 4.5005
R16757 VSS.n0 VSS.n11 4.57442
R16758 VSS.n7 VSS.n8 0.147342
R16759 VSS.n8 VSS.n9 0.147342
R16760 VSS.n9 VSS.n10 0.147342
R16761 VSS.n11 VSS.n12 2.39784
R16762 VSS.n12 VSS.n13 0.147342
R16763 VSS.n13 VSS.n14 0.147342
R16764 VSS.n14 VSS.t461 3.13212
R16765 BIT_SEL[49].t0 BIT_SEL[49] 116.918
R16766 BIT_SEL[49] BIT_SEL[49].n0 11.2682
R16767 BIT_SEL[49] BIT_SEL[49].n0 1.36014
R16768 BIT_SEL[49] BIT_SEL[49].n1 11.2682
R16769 BIT_SEL[49].n1 BIT_SEL[49] 1.36014
R16770 BIT_SEL[49] BIT_SEL[49].n2 11.2682
R16771 BIT_SEL[49].n2 BIT_SEL[49] 1.36014
R16772 BIT_SEL[49] BIT_SEL[49].n3 11.2682
R16773 BIT_SEL[49].n3 BIT_SEL[49] 1.36014
R16774 BIT_SEL[49] BIT_SEL[49].n4 11.2682
R16775 BIT_SEL[49].n4 BIT_SEL[49] 1.36014
R16776 BIT_SEL[49] BIT_SEL[49].n5 11.2682
R16777 BIT_SEL[49].n5 BIT_SEL[49] 1.36014
R16778 BIT_SEL[49] BIT_SEL[49].n6 11.2682
R16779 BIT_SEL[49].n6 BIT_SEL[49] 1.36014
R16780 BIT_SEL[49].t3 BIT_SEL[49].n6 115.558
R16781 BIT_SEL[49].t6 BIT_SEL[49].n5 115.558
R16782 BIT_SEL[49].t2 BIT_SEL[49].n4 115.558
R16783 BIT_SEL[49].t4 BIT_SEL[49].n3 115.558
R16784 BIT_SEL[49].t1 BIT_SEL[49].n2 115.558
R16785 BIT_SEL[49].n1 BIT_SEL[49].t7 115.558
R16786 BIT_SEL[49].n0 BIT_SEL[49].t5 115.558
R16787 a_20810_3154.t0 a_20810_3154.t1 6.02155
R16788 a_638_27395.t0 a_638_27395.n0 7.71211
R16789 a_638_27395.n2 a_638_27395.t9 7.71211
R16790 a_638_27395.n3 a_638_27395.t13 7.71211
R16791 a_638_27395.n4 a_638_27395.t51 7.71211
R16792 a_638_27395.n5 a_638_27395.t56 7.71211
R16793 a_638_27395.n6 a_638_27395.t36 7.71211
R16794 a_638_27395.n7 a_638_27395.t55 7.71211
R16795 a_638_27395.n8 a_638_27395.t38 7.71211
R16796 a_638_27395.n9 a_638_27395.t12 7.71211
R16797 a_638_27395.n10 a_638_27395.t15 7.71211
R16798 a_638_27395.n11 a_638_27395.t41 7.71211
R16799 a_638_27395.n12 a_638_27395.t61 7.71211
R16800 a_638_27395.n13 a_638_27395.t67 7.71211
R16801 a_638_27395.n14 a_638_27395.t33 7.71211
R16802 a_638_27395.n15 a_638_27395.t47 7.71211
R16803 a_638_27395.n16 a_638_27395.t27 7.71211
R16804 a_638_27395.n17 a_638_27395.t11 7.71211
R16805 a_638_27395.n18 a_638_27395.t48 7.71211
R16806 a_638_27395.n19 a_638_27395.t45 7.71211
R16807 a_638_27395.n20 a_638_27395.t37 7.71211
R16808 a_638_27395.n21 a_638_27395.t66 7.71211
R16809 a_638_27395.n22 a_638_27395.t53 7.71211
R16810 a_638_27395.n23 a_638_27395.t3 7.71211
R16811 a_638_27395.n24 a_638_27395.t26 7.71211
R16812 a_638_27395.n25 a_638_27395.t8 7.71211
R16813 a_638_27395.n26 a_638_27395.t31 7.71211
R16814 a_638_27395.n27 a_638_27395.t58 7.71211
R16815 a_638_27395.n28 a_638_27395.t21 7.71211
R16816 a_638_27395.n29 a_638_27395.t1 7.71211
R16817 a_638_27395.n30 a_638_27395.t18 7.71211
R16818 a_638_27395.n31 a_638_27395.t16 7.71211
R16819 a_638_27395.n32 a_638_27395.t17 7.71211
R16820 a_638_27395.n3 a_638_27395.n2 0.427167
R16821 a_638_27395.n4 a_638_27395.n3 0.427167
R16822 a_638_27395.n5 a_638_27395.n4 0.427167
R16823 a_638_27395.n6 a_638_27395.n5 0.427167
R16824 a_638_27395.n7 a_638_27395.n6 0.427167
R16825 a_638_27395.n8 a_638_27395.n7 0.427167
R16826 a_638_27395.n9 a_638_27395.n8 0.427167
R16827 a_638_27395.n10 a_638_27395.n9 0.619389
R16828 a_638_27395.n11 a_638_27395.n10 0.427167
R16829 a_638_27395.n12 a_638_27395.n11 0.427167
R16830 a_638_27395.n13 a_638_27395.n12 0.427167
R16831 a_638_27395.n14 a_638_27395.n13 0.427167
R16832 a_638_27395.n15 a_638_27395.n14 0.427167
R16833 a_638_27395.n16 a_638_27395.n15 0.427167
R16834 a_638_27395.n17 a_638_27395.n16 0.427167
R16835 a_638_27395.n18 a_638_27395.n17 0.619389
R16836 a_638_27395.n19 a_638_27395.n18 0.427167
R16837 a_638_27395.n0 a_638_27395.n19 0.427167
R16838 a_638_27395.n0 a_638_27395.n20 0.427167
R16839 a_638_27395.n20 a_638_27395.n21 0.427167
R16840 a_638_27395.n21 a_638_27395.n22 0.427167
R16841 a_638_27395.n22 a_638_27395.n23 0.427167
R16842 a_638_27395.n23 a_638_27395.n24 0.427167
R16843 a_638_27395.n24 a_638_27395.n25 0.619389
R16844 a_638_27395.n25 a_638_27395.n26 0.427167
R16845 a_638_27395.n26 a_638_27395.n27 0.427167
R16846 a_638_27395.n27 a_638_27395.n28 0.427167
R16847 a_638_27395.n28 a_638_27395.n29 0.427167
R16848 a_638_27395.n29 a_638_27395.n30 0.427167
R16849 a_638_27395.n30 a_638_27395.n31 0.427167
R16850 a_638_27395.n31 a_638_27395.n32 0.427167
R16851 a_638_27395.n32 a_638_27395.n1 0.334944
R16852 a_638_27395.n1 a_638_27395.n33 0.227167
R16853 a_638_27395.n34 a_638_27395.n35 0.466493
R16854 a_638_27395.n2 a_638_27395.n34 0.69448
R16855 a_638_27395.n35 a_638_27395.t5 7.71211
R16856 a_638_27395.n36 a_638_27395.t39 7.71211
R16857 a_638_27395.n37 a_638_27395.t4 7.71211
R16858 a_638_27395.n38 a_638_27395.t42 7.71211
R16859 a_638_27395.n39 a_638_27395.t57 7.71211
R16860 a_638_27395.n40 a_638_27395.t44 7.71211
R16861 a_638_27395.n41 a_638_27395.t65 7.71211
R16862 a_638_27395.n42 a_638_27395.t60 7.71211
R16863 a_638_27395.n43 a_638_27395.t52 7.71211
R16864 a_638_27395.n44 a_638_27395.t46 7.71211
R16865 a_638_27395.n45 a_638_27395.t50 7.71211
R16866 a_638_27395.n46 a_638_27395.t7 7.71211
R16867 a_638_27395.n47 a_638_27395.t2 7.71211
R16868 a_638_27395.n48 a_638_27395.t6 7.71211
R16869 a_638_27395.n49 a_638_27395.t32 7.71211
R16870 a_638_27395.n50 a_638_27395.t30 7.71211
R16871 a_638_27395.n51 a_638_27395.t35 7.71211
R16872 a_638_27395.n52 a_638_27395.t10 7.71211
R16873 a_638_27395.n53 a_638_27395.t63 7.71211
R16874 a_638_27395.n54 a_638_27395.t64 7.71211
R16875 a_638_27395.n55 a_638_27395.t24 7.71211
R16876 a_638_27395.n56 a_638_27395.t62 7.71211
R16877 a_638_27395.n57 a_638_27395.t68 7.71211
R16878 a_638_27395.n58 a_638_27395.t14 7.71211
R16879 a_638_27395.n59 a_638_27395.t43 7.71211
R16880 a_638_27395.n60 a_638_27395.t22 7.71211
R16881 a_638_27395.n61 a_638_27395.t34 7.71211
R16882 a_638_27395.n62 a_638_27395.t40 7.71211
R16883 a_638_27395.n63 a_638_27395.t54 7.71211
R16884 a_638_27395.n64 a_638_27395.t49 7.71211
R16885 a_638_27395.n65 a_638_27395.t59 7.71211
R16886 a_638_27395.n66 a_638_27395.t28 7.71211
R16887 a_638_27395.n35 a_638_27395.n36 0.427167
R16888 a_638_27395.n36 a_638_27395.n37 0.427167
R16889 a_638_27395.n37 a_638_27395.n38 0.427167
R16890 a_638_27395.n38 a_638_27395.n39 0.427167
R16891 a_638_27395.n39 a_638_27395.n40 0.427167
R16892 a_638_27395.n40 a_638_27395.n41 0.427167
R16893 a_638_27395.n41 a_638_27395.n42 0.427167
R16894 a_638_27395.n42 a_638_27395.n43 0.619389
R16895 a_638_27395.n43 a_638_27395.n44 0.427167
R16896 a_638_27395.n44 a_638_27395.n45 0.427167
R16897 a_638_27395.n45 a_638_27395.n46 0.427167
R16898 a_638_27395.n46 a_638_27395.n47 0.427167
R16899 a_638_27395.n47 a_638_27395.n48 0.427167
R16900 a_638_27395.n48 a_638_27395.n49 0.427167
R16901 a_638_27395.n49 a_638_27395.n50 0.427167
R16902 a_638_27395.n50 a_638_27395.n51 0.619389
R16903 a_638_27395.n51 a_638_27395.n52 0.427167
R16904 a_638_27395.n52 a_638_27395.n53 0.427167
R16905 a_638_27395.n53 a_638_27395.n54 0.427167
R16906 a_638_27395.n54 a_638_27395.n55 0.427167
R16907 a_638_27395.n55 a_638_27395.n56 0.427167
R16908 a_638_27395.n56 a_638_27395.n57 0.427167
R16909 a_638_27395.n57 a_638_27395.n58 0.427167
R16910 a_638_27395.n58 a_638_27395.n59 0.619389
R16911 a_638_27395.n60 a_638_27395.n59 0.427167
R16912 a_638_27395.n61 a_638_27395.n60 0.427167
R16913 a_638_27395.n62 a_638_27395.n61 0.427167
R16914 a_638_27395.n63 a_638_27395.n62 0.427167
R16915 a_638_27395.n64 a_638_27395.n63 0.427167
R16916 a_638_27395.n65 a_638_27395.n64 0.427167
R16917 a_638_27395.n66 a_638_27395.n65 0.427167
R16918 a_638_27395.n71 a_638_27395.n66 0.548278
R16919 a_638_27395.n71 a_638_27395.n68 0.227167
R16920 a_638_27395.n72 a_638_27395.n71 4.74618
R16921 a_638_27395.n1 a_638_27395.n72 4.60509
R16922 a_638_27395.n72 a_638_27395.t29 0.113082
R16923 a_638_27395.n70 a_638_27395.n69 0.0655
R16924 a_638_27395.n70 a_638_27395.n68 4.74618
R16925 a_638_27395.n33 a_638_27395.n70 4.60509
R16926 a_638_27395.n69 a_638_27395.t19 0.0480817
R16927 a_638_27395.n69 a_638_27395.t25 0.0480817
R16928 a_638_27395.n68 a_638_27395.n67 4.96756
R16929 a_638_27395.n33 a_638_27395.n67 4.83019
R16930 a_638_27395.n67 a_638_27395.t20 0.113082
R16931 a_638_27395.n34 a_638_27395.t23 9.85476
R16932 a_1340_25152.t0 a_1340_25152.t1 6.39548
R16933 a_110_52624.t0 a_110_52624.t1 19.5535
R16934 a_154_52536.t0 a_154_52536.t1 13.9628
R16935 VDD.n1 VDD.n20 13.5005
R16936 VDD.n2 VDD.n19 13.5005
R16937 VDD.n3 VDD.n18 13.5005
R16938 VDD.n4 VDD.n17 13.5005
R16939 VDD.n5 VDD.n16 13.5005
R16940 VDD.n6 VDD.n13 13.5005
R16941 VDD.n7 VDD.n12 13.5005
R16942 VDD.n8 VDD.n11 13.5005
R16943 VDD.n9 VDD.n10 13.5005
R16944 VDD.n1 VDD.n32 13.5005
R16945 VDD.n2 VDD.n31 13.5005
R16946 VDD.n3 VDD.n30 13.5005
R16947 VDD.n4 VDD.n29 13.5005
R16948 VDD.n5 VDD.n28 13.5005
R16949 VDD.n6 VDD.n25 13.5005
R16950 VDD.n7 VDD.n24 13.5005
R16951 VDD.n8 VDD.n23 13.5005
R16952 VDD.n9 VDD.n22 13.5005
R16953 VDD.n266 VDD.n1 0.0319875
R16954 VDD.n267 VDD.n2 13.5005
R16955 VDD.n268 VDD.n3 13.5005
R16956 VDD.n269 VDD.n4 13.5005
R16957 VDD.n270 VDD.n5 13.5005
R16958 VDD.n271 VDD.n6 13.5005
R16959 VDD.n272 VDD.n7 13.5005
R16960 VDD.n273 VDD.n8 13.5005
R16961 VDD.n274 VDD.n9 0.0319875
R16962 VDD.n34 VDD.n53 13.5005
R16963 VDD.n35 VDD.n52 13.5005
R16964 VDD.n36 VDD.n51 13.5005
R16965 VDD.n37 VDD.n50 13.5005
R16966 VDD.n38 VDD.n49 13.5005
R16967 VDD.n39 VDD.n46 13.5005
R16968 VDD.n40 VDD.n45 13.5005
R16969 VDD.n41 VDD.n44 13.5005
R16970 VDD.n42 VDD.n43 13.5005
R16971 VDD.n34 VDD.n65 13.5005
R16972 VDD.n35 VDD.n64 13.5005
R16973 VDD.n36 VDD.n63 13.5005
R16974 VDD.n37 VDD.n62 13.5005
R16975 VDD.n38 VDD.n61 13.5005
R16976 VDD.n39 VDD.n58 13.5005
R16977 VDD.n40 VDD.n57 13.5005
R16978 VDD.n41 VDD.n56 13.5005
R16979 VDD.n42 VDD.n55 13.5005
R16980 VDD.n276 VDD.n34 0.0319875
R16981 VDD.n277 VDD.n35 13.5005
R16982 VDD.n278 VDD.n36 13.5005
R16983 VDD.n279 VDD.n37 13.5005
R16984 VDD.n280 VDD.n38 13.5005
R16985 VDD.n281 VDD.n39 13.5005
R16986 VDD.n282 VDD.n40 13.5005
R16987 VDD.n283 VDD.n41 13.5005
R16988 VDD.n284 VDD.n42 0.0319875
R16989 VDD.n67 VDD.n86 13.5005
R16990 VDD.n68 VDD.n85 13.5005
R16991 VDD.n69 VDD.n84 13.5005
R16992 VDD.n70 VDD.n83 13.5005
R16993 VDD.n71 VDD.n82 13.5005
R16994 VDD.n72 VDD.n79 13.5005
R16995 VDD.n73 VDD.n78 13.5005
R16996 VDD.n74 VDD.n77 13.5005
R16997 VDD.n75 VDD.n76 13.5005
R16998 VDD.n67 VDD.n98 13.5005
R16999 VDD.n68 VDD.n97 13.5005
R17000 VDD.n69 VDD.n96 13.5005
R17001 VDD.n70 VDD.n95 13.5005
R17002 VDD.n71 VDD.n94 13.5005
R17003 VDD.n72 VDD.n91 13.5005
R17004 VDD.n73 VDD.n90 13.5005
R17005 VDD.n74 VDD.n89 13.5005
R17006 VDD.n75 VDD.n88 13.5005
R17007 VDD.n286 VDD.n67 0.0319875
R17008 VDD.n287 VDD.n68 13.5005
R17009 VDD.n288 VDD.n69 13.5005
R17010 VDD.n289 VDD.n70 13.5005
R17011 VDD.n290 VDD.n71 13.5005
R17012 VDD.n291 VDD.n72 13.5005
R17013 VDD.n292 VDD.n73 13.5005
R17014 VDD.n293 VDD.n74 13.5005
R17015 VDD.n294 VDD.n75 0.0319875
R17016 VDD.n100 VDD.n119 13.5005
R17017 VDD.n101 VDD.n118 13.5005
R17018 VDD.n102 VDD.n117 13.5005
R17019 VDD.n103 VDD.n116 13.5005
R17020 VDD.n104 VDD.n115 13.5005
R17021 VDD.n105 VDD.n112 13.5005
R17022 VDD.n106 VDD.n111 13.5005
R17023 VDD.n107 VDD.n110 13.5005
R17024 VDD.n108 VDD.n109 13.5005
R17025 VDD.n100 VDD.n131 13.5005
R17026 VDD.n101 VDD.n130 13.5005
R17027 VDD.n102 VDD.n129 13.5005
R17028 VDD.n103 VDD.n128 13.5005
R17029 VDD.n104 VDD.n127 13.5005
R17030 VDD.n105 VDD.n124 13.5005
R17031 VDD.n106 VDD.n123 13.5005
R17032 VDD.n107 VDD.n122 13.5005
R17033 VDD.n108 VDD.n121 13.5005
R17034 VDD.n296 VDD.n100 0.0319875
R17035 VDD.n297 VDD.n101 13.5005
R17036 VDD.n298 VDD.n102 13.5005
R17037 VDD.n299 VDD.n103 13.5005
R17038 VDD.n300 VDD.n104 13.5005
R17039 VDD.n301 VDD.n105 13.5005
R17040 VDD.n302 VDD.n106 13.5005
R17041 VDD.n303 VDD.n107 13.5005
R17042 VDD.n304 VDD.n108 0.0319875
R17043 VDD.n133 VDD.n152 13.5005
R17044 VDD.n134 VDD.n151 13.5005
R17045 VDD.n135 VDD.n150 13.5005
R17046 VDD.n136 VDD.n149 13.5005
R17047 VDD.n137 VDD.n148 13.5005
R17048 VDD.n138 VDD.n145 13.5005
R17049 VDD.n139 VDD.n144 13.5005
R17050 VDD.n140 VDD.n143 13.5005
R17051 VDD.n141 VDD.n142 13.5005
R17052 VDD.n133 VDD.n164 13.5005
R17053 VDD.n134 VDD.n163 13.5005
R17054 VDD.n135 VDD.n162 13.5005
R17055 VDD.n136 VDD.n161 13.5005
R17056 VDD.n137 VDD.n160 13.5005
R17057 VDD.n138 VDD.n157 13.5005
R17058 VDD.n139 VDD.n156 13.5005
R17059 VDD.n140 VDD.n155 13.5005
R17060 VDD.n141 VDD.n154 13.5005
R17061 VDD.n306 VDD.n133 0.0319875
R17062 VDD.n307 VDD.n134 13.5005
R17063 VDD.n308 VDD.n135 13.5005
R17064 VDD.n309 VDD.n136 13.5005
R17065 VDD.n310 VDD.n137 13.5005
R17066 VDD.n311 VDD.n138 13.5005
R17067 VDD.n312 VDD.n139 13.5005
R17068 VDD.n313 VDD.n140 13.5005
R17069 VDD.n314 VDD.n141 0.0319875
R17070 VDD.n166 VDD.n185 13.5005
R17071 VDD.n167 VDD.n184 13.5005
R17072 VDD.n168 VDD.n183 13.5005
R17073 VDD.n169 VDD.n182 13.5005
R17074 VDD.n170 VDD.n181 13.5005
R17075 VDD.n178 VDD.n171 13.5005
R17076 VDD.n177 VDD.n172 13.5005
R17077 VDD.n176 VDD.n173 13.5005
R17078 VDD.n175 VDD.n174 13.5005
R17079 VDD.n166 VDD.n197 13.5005
R17080 VDD.n167 VDD.n196 13.5005
R17081 VDD.n168 VDD.n195 13.5005
R17082 VDD.n169 VDD.n194 13.5005
R17083 VDD.n170 VDD.n193 13.5005
R17084 VDD.n190 VDD.n171 13.5005
R17085 VDD.n189 VDD.n172 13.5005
R17086 VDD.n188 VDD.n173 13.5005
R17087 VDD.n187 VDD.n174 13.5005
R17088 VDD.n316 VDD.n166 0.0319875
R17089 VDD.n317 VDD.n167 13.5005
R17090 VDD.n318 VDD.n168 13.5005
R17091 VDD.n319 VDD.n169 13.5005
R17092 VDD.n320 VDD.n170 13.5005
R17093 VDD.n321 VDD.n171 13.5005
R17094 VDD.n322 VDD.n172 13.5005
R17095 VDD.n323 VDD.n173 13.5005
R17096 VDD.n324 VDD.n174 0.0319875
R17097 VDD.n199 VDD.n218 13.5005
R17098 VDD.n200 VDD.n217 13.5005
R17099 VDD.n201 VDD.n216 13.5005
R17100 VDD.n202 VDD.n215 13.5005
R17101 VDD.n203 VDD.n214 13.5005
R17102 VDD.n204 VDD.n211 13.5005
R17103 VDD.n205 VDD.n210 13.5005
R17104 VDD.n206 VDD.n209 13.5005
R17105 VDD.n207 VDD.n208 13.5005
R17106 VDD.n199 VDD.n230 13.5005
R17107 VDD.n200 VDD.n229 13.5005
R17108 VDD.n201 VDD.n228 13.5005
R17109 VDD.n202 VDD.n227 13.5005
R17110 VDD.n203 VDD.n226 13.5005
R17111 VDD.n204 VDD.n223 13.5005
R17112 VDD.n205 VDD.n222 13.5005
R17113 VDD.n206 VDD.n221 13.5005
R17114 VDD.n207 VDD.n220 13.5005
R17115 VDD.n199 VDD.n326 0.0319875
R17116 VDD.n327 VDD.n200 13.5005
R17117 VDD.n328 VDD.n201 13.5005
R17118 VDD.n329 VDD.n202 13.5005
R17119 VDD.n330 VDD.n203 13.5005
R17120 VDD.n331 VDD.n204 13.5005
R17121 VDD.n332 VDD.n205 13.5005
R17122 VDD.n333 VDD.n206 13.5005
R17123 VDD.n207 VDD.n334 0.0319875
R17124 VDD.n251 VDD.n232 13.5005
R17125 VDD.n250 VDD.n233 13.5005
R17126 VDD.n249 VDD.n234 13.5005
R17127 VDD.n248 VDD.n235 13.5005
R17128 VDD.n247 VDD.n236 13.5005
R17129 VDD.n237 VDD.n244 13.5005
R17130 VDD.n238 VDD.n243 13.5005
R17131 VDD.n239 VDD.n242 13.5005
R17132 VDD.n240 VDD.n241 13.5005
R17133 VDD.n263 VDD.n232 13.5005
R17134 VDD.n262 VDD.n233 13.5005
R17135 VDD.n261 VDD.n234 13.5005
R17136 VDD.n260 VDD.n235 13.5005
R17137 VDD.n259 VDD.n236 13.5005
R17138 VDD.n237 VDD.n256 13.5005
R17139 VDD.n238 VDD.n255 13.5005
R17140 VDD.n239 VDD.n254 13.5005
R17141 VDD.n240 VDD.n253 13.5005
R17142 VDD.n337 VDD.n232 0.0319875
R17143 VDD.n338 VDD.n233 13.5005
R17144 VDD.n339 VDD.n234 13.5005
R17145 VDD.n340 VDD.n235 13.5005
R17146 VDD.n341 VDD.n236 13.5005
R17147 VDD.n342 VDD.n237 13.5005
R17148 VDD.n343 VDD.n238 13.5005
R17149 VDD.n344 VDD.n239 13.5005
R17150 VDD.n264 VDD.n240 0.0319875
R17151 VDD.n337 VDD.n231 0.0333961
R17152 VDD.n232 VDD.n233 0.0640294
R17153 VDD.n233 VDD.n234 0.0640294
R17154 VDD.n234 VDD.n235 0.0640294
R17155 VDD.n235 VDD.n236 0.0640294
R17156 VDD.n236 VDD 0.0574647
R17157 VDD VDD.n237 0.0705941
R17158 VDD.n238 VDD.n237 0.0640294
R17159 VDD.n239 VDD.n238 0.0640294
R17160 VDD.n240 VDD.n239 0.0640294
R17161 VDD.n252 VDD.n264 0.0333961
R17162 VDD.n198 VDD.n252 0.135712
R17163 VDD.n326 VDD.n198 0.0333961
R17164 VDD.n200 VDD.n199 0.0640294
R17165 VDD.n201 VDD.n200 0.0640294
R17166 VDD.n202 VDD.n201 0.0640294
R17167 VDD.n203 VDD.n202 0.0640294
R17168 VDD VDD.n203 0.0574647
R17169 VDD VDD.n204 0.0705941
R17170 VDD.n204 VDD.n205 0.0640294
R17171 VDD.n205 VDD.n206 0.0640294
R17172 VDD.n206 VDD.n207 0.0640294
R17173 VDD.n334 VDD.n219 0.0333961
R17174 VDD.n219 VDD.n165 0.135712
R17175 VDD.n165 VDD.n316 0.0333961
R17176 VDD.n166 VDD.n167 0.0640294
R17177 VDD.n167 VDD.n168 0.0640294
R17178 VDD.n168 VDD.n169 0.0640294
R17179 VDD.n169 VDD.n170 0.0640294
R17180 VDD.n170 VDD 0.0574647
R17181 VDD VDD.n171 0.0705941
R17182 VDD.n172 VDD.n171 0.0640294
R17183 VDD.n173 VDD.n172 0.0640294
R17184 VDD.n174 VDD.n173 0.0640294
R17185 VDD.n324 VDD.n186 0.0333961
R17186 VDD.n186 VDD.n132 0.135712
R17187 VDD.n132 VDD.n306 0.0333961
R17188 VDD.n133 VDD.n134 0.0640294
R17189 VDD.n134 VDD.n135 0.0640294
R17190 VDD.n135 VDD.n136 0.0640294
R17191 VDD.n136 VDD.n137 0.0640294
R17192 VDD.n137 VDD 0.0574647
R17193 VDD VDD.n138 0.0705941
R17194 VDD.n139 VDD.n138 0.0640294
R17195 VDD.n140 VDD.n139 0.0640294
R17196 VDD.n141 VDD.n140 0.0640294
R17197 VDD.n314 VDD.n153 0.0333961
R17198 VDD.n153 VDD.n99 0.135712
R17199 VDD.n99 VDD.n296 0.0333961
R17200 VDD.n100 VDD.n101 0.0640294
R17201 VDD.n101 VDD.n102 0.0640294
R17202 VDD.n102 VDD.n103 0.0640294
R17203 VDD.n103 VDD.n104 0.0640294
R17204 VDD.n104 VDD 0.0574647
R17205 VDD VDD.n105 0.0705941
R17206 VDD.n106 VDD.n105 0.0640294
R17207 VDD.n107 VDD.n106 0.0640294
R17208 VDD.n108 VDD.n107 0.0640294
R17209 VDD.n304 VDD.n120 0.0333961
R17210 VDD.n120 VDD.n66 0.135712
R17211 VDD.n66 VDD.n286 0.0333961
R17212 VDD.n67 VDD.n68 0.0640294
R17213 VDD.n68 VDD.n69 0.0640294
R17214 VDD.n69 VDD.n70 0.0640294
R17215 VDD.n70 VDD.n71 0.0640294
R17216 VDD.n71 VDD 0.0574647
R17217 VDD VDD.n72 0.0705941
R17218 VDD.n73 VDD.n72 0.0640294
R17219 VDD.n74 VDD.n73 0.0640294
R17220 VDD.n75 VDD.n74 0.0640294
R17221 VDD.n294 VDD.n87 0.0333961
R17222 VDD.n87 VDD.n33 0.135712
R17223 VDD.n33 VDD.n276 0.0333961
R17224 VDD.n34 VDD.n35 0.0640294
R17225 VDD.n35 VDD.n36 0.0640294
R17226 VDD.n36 VDD.n37 0.0640294
R17227 VDD.n37 VDD.n38 0.0640294
R17228 VDD.n38 VDD 0.0574647
R17229 VDD VDD.n39 0.0705941
R17230 VDD.n40 VDD.n39 0.0640294
R17231 VDD.n41 VDD.n40 0.0640294
R17232 VDD.n42 VDD.n41 0.0640294
R17233 VDD.n284 VDD.n54 0.0333961
R17234 VDD.n54 VDD.n0 0.135712
R17235 VDD.n0 VDD.n266 0.0333961
R17236 VDD.n1 VDD.n2 0.0640294
R17237 VDD.n2 VDD.n3 0.0640294
R17238 VDD.n3 VDD.n4 0.0640294
R17239 VDD.n4 VDD.n5 0.0640294
R17240 VDD.n5 VDD 0.0574647
R17241 VDD VDD.n6 0.0705941
R17242 VDD.n7 VDD.n6 0.0640294
R17243 VDD.n8 VDD.n7 0.0640294
R17244 VDD.n9 VDD.n8 0.0640294
R17245 VDD.n274 VDD.n21 0.0333961
R17246 VDD.n265 VDD.n336 0.158
R17247 VDD.n338 VDD.n337 7.4988
R17248 VDD.n339 VDD.n338 0.614136
R17249 VDD.n340 VDD.n339 0.614136
R17250 VDD.n341 VDD.n340 0.614136
R17251 VDD.n336 VDD.n341 0.550727
R17252 VDD.n342 VDD.n336 0.677545
R17253 VDD.n343 VDD.n342 0.614136
R17254 VDD.n344 VDD.n343 0.614136
R17255 VDD.n264 VDD.n344 7.4988
R17256 VDD.n265 VDD.n275 0.158
R17257 VDD.n265 VDD.n285 0.158
R17258 VDD.n265 VDD.n295 0.158
R17259 VDD.n265 VDD.n305 0.158
R17260 VDD.n265 VDD.n315 0.158
R17261 VDD.n265 VDD.n325 0.158
R17262 VDD.n335 VDD.n265 0.158
R17263 VDD.t76 VDD.t6 3.23711
R17264 VDD.t86 VDD.t76 3.23711
R17265 VDD.t2 VDD.t86 3.23711
R17266 VDD.n265 VDD.t2 4.03039
R17267 VDD.n326 VDD.n327 7.4988
R17268 VDD.n327 VDD.n328 0.614136
R17269 VDD.n328 VDD.n329 0.614136
R17270 VDD.n329 VDD.n330 0.614136
R17271 VDD.n330 VDD.n335 0.550727
R17272 VDD.n331 VDD.n335 0.677545
R17273 VDD.n332 VDD.n331 0.614136
R17274 VDD.n333 VDD.n332 0.614136
R17275 VDD.n334 VDD.n333 7.4988
R17276 VDD.n316 VDD.n317 7.4988
R17277 VDD.n317 VDD.n318 0.614136
R17278 VDD.n318 VDD.n319 0.614136
R17279 VDD.n319 VDD.n320 0.614136
R17280 VDD.n320 VDD.n325 0.550727
R17281 VDD.n325 VDD.n321 0.677545
R17282 VDD.n321 VDD.n322 0.614136
R17283 VDD.n322 VDD.n323 0.614136
R17284 VDD.n323 VDD.n324 7.4988
R17285 VDD.n306 VDD.n307 7.4988
R17286 VDD.n308 VDD.n307 0.614136
R17287 VDD.n309 VDD.n308 0.614136
R17288 VDD.n310 VDD.n309 0.614136
R17289 VDD.n315 VDD.n310 0.550727
R17290 VDD.n315 VDD.n311 0.677545
R17291 VDD.n311 VDD.n312 0.614136
R17292 VDD.n312 VDD.n313 0.614136
R17293 VDD.n313 VDD.n314 7.4988
R17294 VDD.n296 VDD.n297 7.4988
R17295 VDD.n298 VDD.n297 0.614136
R17296 VDD.n299 VDD.n298 0.614136
R17297 VDD.n300 VDD.n299 0.614136
R17298 VDD.n305 VDD.n300 0.550727
R17299 VDD.n305 VDD.n301 0.677545
R17300 VDD.n301 VDD.n302 0.614136
R17301 VDD.n302 VDD.n303 0.614136
R17302 VDD.n303 VDD.n304 7.4988
R17303 VDD.n286 VDD.n287 7.4988
R17304 VDD.n288 VDD.n287 0.614136
R17305 VDD.n289 VDD.n288 0.614136
R17306 VDD.n290 VDD.n289 0.614136
R17307 VDD.n295 VDD.n290 0.550727
R17308 VDD.n295 VDD.n291 0.677545
R17309 VDD.n291 VDD.n292 0.614136
R17310 VDD.n292 VDD.n293 0.614136
R17311 VDD.n293 VDD.n294 7.4988
R17312 VDD.n276 VDD.n277 7.4988
R17313 VDD.n278 VDD.n277 0.614136
R17314 VDD.n279 VDD.n278 0.614136
R17315 VDD.n280 VDD.n279 0.614136
R17316 VDD.n285 VDD.n280 0.550727
R17317 VDD.n285 VDD.n281 0.677545
R17318 VDD.n281 VDD.n282 0.614136
R17319 VDD.n282 VDD.n283 0.614136
R17320 VDD.n283 VDD.n284 7.4988
R17321 VDD.n266 VDD.n267 7.4988
R17322 VDD.n268 VDD.n267 0.614136
R17323 VDD.n269 VDD.n268 0.614136
R17324 VDD.n270 VDD.n269 0.614136
R17325 VDD.n275 VDD.n270 0.550727
R17326 VDD.n275 VDD.n271 0.677545
R17327 VDD.n271 VDD.n272 0.614136
R17328 VDD.n272 VDD.n273 0.614136
R17329 VDD.n273 VDD.n274 7.4988
R17330 VDD.n253 VDD.n252 14.2278
R17331 VDD.n254 VDD.n253 0.727797
R17332 VDD.n255 VDD.n254 0.727797
R17333 VDD.n256 VDD.n255 0.727797
R17334 VDD.n258 VDD.n257 0.0655
R17335 VDD.n256 VDD.n258 0.804419
R17336 VDD.n258 VDD.n259 0.653608
R17337 VDD.n259 VDD.n260 0.727797
R17338 VDD.n260 VDD.n261 0.727797
R17339 VDD.n261 VDD.n262 0.727797
R17340 VDD.n262 VDD.n263 0.727797
R17341 VDD.n231 VDD.n263 14.2278
R17342 VDD.n257 VDD.t111 0.0480817
R17343 VDD.n257 VDD.t75 0.0480817
R17344 VDD.n241 VDD.n252 14.2278
R17345 VDD.n242 VDD.n241 0.727797
R17346 VDD.n243 VDD.n242 0.727797
R17347 VDD.n244 VDD.n243 0.727797
R17348 VDD.n246 VDD.n245 0.0655
R17349 VDD.n244 VDD.n246 0.804419
R17350 VDD.n246 VDD.n247 0.653608
R17351 VDD.n247 VDD.n248 0.727797
R17352 VDD.n248 VDD.n249 0.727797
R17353 VDD.n249 VDD.n250 0.727797
R17354 VDD.n250 VDD.n251 0.727797
R17355 VDD.n231 VDD.n251 14.2278
R17356 VDD.n245 VDD.t46 0.0480817
R17357 VDD.n245 VDD.t77 0.0480817
R17358 VDD.n220 VDD.n219 14.2278
R17359 VDD.n221 VDD.n220 0.727797
R17360 VDD.n222 VDD.n221 0.727797
R17361 VDD.n223 VDD.n222 0.727797
R17362 VDD.n225 VDD.n224 0.0655
R17363 VDD.n225 VDD.n223 0.804419
R17364 VDD.n226 VDD.n225 0.653608
R17365 VDD.n227 VDD.n226 0.727797
R17366 VDD.n228 VDD.n227 0.727797
R17367 VDD.n229 VDD.n228 0.727797
R17368 VDD.n230 VDD.n229 0.727797
R17369 VDD.n198 VDD.n230 14.2278
R17370 VDD.n224 VDD.t121 0.0480817
R17371 VDD.n224 VDD.t282 0.0480817
R17372 VDD.n208 VDD.n219 14.2278
R17373 VDD.n209 VDD.n208 0.727797
R17374 VDD.n210 VDD.n209 0.727797
R17375 VDD.n211 VDD.n210 0.727797
R17376 VDD.n213 VDD.n212 0.0655
R17377 VDD.n213 VDD.n211 0.804419
R17378 VDD.n214 VDD.n213 0.653608
R17379 VDD.n215 VDD.n214 0.727797
R17380 VDD.n216 VDD.n215 0.727797
R17381 VDD.n217 VDD.n216 0.727797
R17382 VDD.n218 VDD.n217 0.727797
R17383 VDD.n198 VDD.n218 14.2278
R17384 VDD.n212 VDD.t120 0.0480817
R17385 VDD.n212 VDD.t289 0.0480817
R17386 VDD.n187 VDD.n186 14.2278
R17387 VDD.n188 VDD.n187 0.727797
R17388 VDD.n189 VDD.n188 0.727797
R17389 VDD.n190 VDD.n189 0.727797
R17390 VDD.n192 VDD.n191 0.0655
R17391 VDD.n192 VDD.n190 0.804419
R17392 VDD.n193 VDD.n192 0.653608
R17393 VDD.n194 VDD.n193 0.727797
R17394 VDD.n195 VDD.n194 0.727797
R17395 VDD.n196 VDD.n195 0.727797
R17396 VDD.n197 VDD.n196 0.727797
R17397 VDD.n165 VDD.n197 14.2278
R17398 VDD.n191 VDD.t261 0.0480817
R17399 VDD.n191 VDD.t262 0.0480817
R17400 VDD.n175 VDD.n186 14.2278
R17401 VDD.n176 VDD.n175 0.727797
R17402 VDD.n177 VDD.n176 0.727797
R17403 VDD.n178 VDD.n177 0.727797
R17404 VDD.n180 VDD.n179 0.0655
R17405 VDD.n180 VDD.n178 0.804419
R17406 VDD.n181 VDD.n180 0.653608
R17407 VDD.n182 VDD.n181 0.727797
R17408 VDD.n183 VDD.n182 0.727797
R17409 VDD.n184 VDD.n183 0.727797
R17410 VDD.n185 VDD.n184 0.727797
R17411 VDD.n165 VDD.n185 14.2278
R17412 VDD.n179 VDD.t247 0.0480817
R17413 VDD.n179 VDD.t263 0.0480817
R17414 VDD.n154 VDD.n153 14.2278
R17415 VDD.n155 VDD.n154 0.727797
R17416 VDD.n156 VDD.n155 0.727797
R17417 VDD.n157 VDD.n156 0.727797
R17418 VDD.n159 VDD.n158 0.0655
R17419 VDD.n157 VDD.n159 0.804419
R17420 VDD.n160 VDD.n159 0.653608
R17421 VDD.n161 VDD.n160 0.727797
R17422 VDD.n162 VDD.n161 0.727797
R17423 VDD.n163 VDD.n162 0.727797
R17424 VDD.n164 VDD.n163 0.727797
R17425 VDD.n132 VDD.n164 14.2278
R17426 VDD.n158 VDD.t140 0.0480817
R17427 VDD.n158 VDD.t125 0.0480817
R17428 VDD.n142 VDD.n153 14.2278
R17429 VDD.n143 VDD.n142 0.727797
R17430 VDD.n144 VDD.n143 0.727797
R17431 VDD.n145 VDD.n144 0.727797
R17432 VDD.n147 VDD.n146 0.0655
R17433 VDD.n145 VDD.n147 0.804419
R17434 VDD.n148 VDD.n147 0.653608
R17435 VDD.n149 VDD.n148 0.727797
R17436 VDD.n150 VDD.n149 0.727797
R17437 VDD.n151 VDD.n150 0.727797
R17438 VDD.n152 VDD.n151 0.727797
R17439 VDD.n132 VDD.n152 14.2278
R17440 VDD.n146 VDD.t167 0.0480817
R17441 VDD.n146 VDD.t124 0.0480817
R17442 VDD.n121 VDD.n120 14.2278
R17443 VDD.n122 VDD.n121 0.727797
R17444 VDD.n123 VDD.n122 0.727797
R17445 VDD.n124 VDD.n123 0.727797
R17446 VDD.n126 VDD.n125 0.0655
R17447 VDD.n124 VDD.n126 0.804419
R17448 VDD.n127 VDD.n126 0.653608
R17449 VDD.n128 VDD.n127 0.727797
R17450 VDD.n129 VDD.n128 0.727797
R17451 VDD.n130 VDD.n129 0.727797
R17452 VDD.n131 VDD.n130 0.727797
R17453 VDD.n99 VDD.n131 14.2278
R17454 VDD.n125 VDD.t209 0.0480817
R17455 VDD.n125 VDD.t3 0.0480817
R17456 VDD.n109 VDD.n120 14.2278
R17457 VDD.n110 VDD.n109 0.727797
R17458 VDD.n111 VDD.n110 0.727797
R17459 VDD.n112 VDD.n111 0.727797
R17460 VDD.n114 VDD.n113 0.0655
R17461 VDD.n112 VDD.n114 0.804419
R17462 VDD.n115 VDD.n114 0.653608
R17463 VDD.n116 VDD.n115 0.727797
R17464 VDD.n117 VDD.n116 0.727797
R17465 VDD.n118 VDD.n117 0.727797
R17466 VDD.n119 VDD.n118 0.727797
R17467 VDD.n99 VDD.n119 14.2278
R17468 VDD.n113 VDD.t7 0.0480817
R17469 VDD.n113 VDD.t208 0.0480817
R17470 VDD.n88 VDD.n87 14.2278
R17471 VDD.n89 VDD.n88 0.727797
R17472 VDD.n90 VDD.n89 0.727797
R17473 VDD.n91 VDD.n90 0.727797
R17474 VDD.n93 VDD.n92 0.0655
R17475 VDD.n91 VDD.n93 0.804419
R17476 VDD.n94 VDD.n93 0.653608
R17477 VDD.n95 VDD.n94 0.727797
R17478 VDD.n96 VDD.n95 0.727797
R17479 VDD.n97 VDD.n96 0.727797
R17480 VDD.n98 VDD.n97 0.727797
R17481 VDD.n66 VDD.n98 14.2278
R17482 VDD.n92 VDD.t166 0.0480817
R17483 VDD.n92 VDD.t141 0.0480817
R17484 VDD.n76 VDD.n87 14.2278
R17485 VDD.n77 VDD.n76 0.727797
R17486 VDD.n78 VDD.n77 0.727797
R17487 VDD.n79 VDD.n78 0.727797
R17488 VDD.n81 VDD.n80 0.0655
R17489 VDD.n79 VDD.n81 0.804419
R17490 VDD.n82 VDD.n81 0.653608
R17491 VDD.n83 VDD.n82 0.727797
R17492 VDD.n84 VDD.n83 0.727797
R17493 VDD.n85 VDD.n84 0.727797
R17494 VDD.n86 VDD.n85 0.727797
R17495 VDD.n66 VDD.n86 14.2278
R17496 VDD.n80 VDD.t123 0.0480817
R17497 VDD.n80 VDD.t122 0.0480817
R17498 VDD.n55 VDD.n54 14.2278
R17499 VDD.n56 VDD.n55 0.727797
R17500 VDD.n57 VDD.n56 0.727797
R17501 VDD.n58 VDD.n57 0.727797
R17502 VDD.n60 VDD.n59 0.0655
R17503 VDD.n58 VDD.n60 0.804419
R17504 VDD.n61 VDD.n60 0.653608
R17505 VDD.n62 VDD.n61 0.727797
R17506 VDD.n63 VDD.n62 0.727797
R17507 VDD.n64 VDD.n63 0.727797
R17508 VDD.n65 VDD.n64 0.727797
R17509 VDD.n33 VDD.n65 14.2278
R17510 VDD.n59 VDD.t254 0.0480817
R17511 VDD.n59 VDD.t252 0.0480817
R17512 VDD.n43 VDD.n54 14.2278
R17513 VDD.n44 VDD.n43 0.727797
R17514 VDD.n45 VDD.n44 0.727797
R17515 VDD.n46 VDD.n45 0.727797
R17516 VDD.n48 VDD.n47 0.0655
R17517 VDD.n46 VDD.n48 0.804419
R17518 VDD.n49 VDD.n48 0.653608
R17519 VDD.n50 VDD.n49 0.727797
R17520 VDD.n51 VDD.n50 0.727797
R17521 VDD.n52 VDD.n51 0.727797
R17522 VDD.n53 VDD.n52 0.727797
R17523 VDD.n33 VDD.n53 14.2278
R17524 VDD.n47 VDD.t246 0.0480817
R17525 VDD.n47 VDD.t253 0.0480817
R17526 VDD.n22 VDD.n21 14.2278
R17527 VDD.n23 VDD.n22 0.727797
R17528 VDD.n24 VDD.n23 0.727797
R17529 VDD.n25 VDD.n24 0.727797
R17530 VDD.n27 VDD.n26 0.0655
R17531 VDD.n25 VDD.n27 0.804419
R17532 VDD.n28 VDD.n27 0.653608
R17533 VDD.n29 VDD.n28 0.727797
R17534 VDD.n30 VDD.n29 0.727797
R17535 VDD.n31 VDD.n30 0.727797
R17536 VDD.n32 VDD.n31 0.727797
R17537 VDD.n0 VDD.n32 14.2278
R17538 VDD.n26 VDD.t87 0.0480817
R17539 VDD.n26 VDD.t89 0.0480817
R17540 VDD.n10 VDD.n21 14.2278
R17541 VDD.n11 VDD.n10 0.727797
R17542 VDD.n12 VDD.n11 0.727797
R17543 VDD.n13 VDD.n12 0.727797
R17544 VDD.n15 VDD.n14 0.0655
R17545 VDD.n13 VDD.n15 0.804419
R17546 VDD.n16 VDD.n15 0.653608
R17547 VDD.n17 VDD.n16 0.727797
R17548 VDD.n18 VDD.n17 0.727797
R17549 VDD.n19 VDD.n18 0.727797
R17550 VDD.n20 VDD.n19 0.727797
R17551 VDD.n0 VDD.n20 14.2278
R17552 VDD.n14 VDD.t88 0.0480817
R17553 VDD.n14 VDD.t90 0.0480817
R17554 a_638_35272.t0 a_638_35272.n0 7.71211
R17555 a_638_35272.n1 a_638_35272.t68 7.71211
R17556 a_638_35272.n2 a_638_35272.t56 7.71211
R17557 a_638_35272.n3 a_638_35272.t63 7.71211
R17558 a_638_35272.n4 a_638_35272.t38 7.71211
R17559 a_638_35272.n5 a_638_35272.t60 7.71211
R17560 a_638_35272.n6 a_638_35272.t14 7.71211
R17561 a_638_35272.n7 a_638_35272.t52 7.71211
R17562 a_638_35272.n8 a_638_35272.t34 7.71211
R17563 a_638_35272.n9 a_638_35272.t33 7.71211
R17564 a_638_35272.n10 a_638_35272.t15 7.71211
R17565 a_638_35272.n11 a_638_35272.t47 7.71211
R17566 a_638_35272.n12 a_638_35272.t6 7.71211
R17567 a_638_35272.n13 a_638_35272.t24 7.71211
R17568 a_638_35272.n14 a_638_35272.t1 7.71211
R17569 a_638_35272.n15 a_638_35272.t62 7.71211
R17570 a_638_35272.n16 a_638_35272.t30 7.71211
R17571 a_638_35272.n17 a_638_35272.t8 7.71211
R17572 a_638_35272.n18 a_638_35272.t11 7.71211
R17573 a_638_35272.n19 a_638_35272.t43 7.71211
R17574 a_638_35272.n20 a_638_35272.t37 7.71211
R17575 a_638_35272.n21 a_638_35272.t49 7.71211
R17576 a_638_35272.n22 a_638_35272.t39 7.71211
R17577 a_638_35272.n23 a_638_35272.t46 7.71211
R17578 a_638_35272.n24 a_638_35272.t50 7.71211
R17579 a_638_35272.n25 a_638_35272.t48 7.71211
R17580 a_638_35272.n26 a_638_35272.t5 7.71211
R17581 a_638_35272.n27 a_638_35272.t67 7.71211
R17582 a_638_35272.n28 a_638_35272.t57 7.71211
R17583 a_638_35272.n29 a_638_35272.t40 7.71211
R17584 a_638_35272.n30 a_638_35272.t12 7.71211
R17585 a_638_35272.n31 a_638_35272.t29 7.71211
R17586 a_638_35272.n2 a_638_35272.n1 0.427167
R17587 a_638_35272.n3 a_638_35272.n2 0.427167
R17588 a_638_35272.n4 a_638_35272.n3 0.427167
R17589 a_638_35272.n5 a_638_35272.n4 0.427167
R17590 a_638_35272.n6 a_638_35272.n5 0.427167
R17591 a_638_35272.n7 a_638_35272.n6 0.427167
R17592 a_638_35272.n8 a_638_35272.n7 0.427167
R17593 a_638_35272.n9 a_638_35272.n8 0.619389
R17594 a_638_35272.n10 a_638_35272.n9 0.427167
R17595 a_638_35272.n11 a_638_35272.n10 0.427167
R17596 a_638_35272.n12 a_638_35272.n11 0.427167
R17597 a_638_35272.n13 a_638_35272.n12 0.427167
R17598 a_638_35272.n14 a_638_35272.n13 0.427167
R17599 a_638_35272.n15 a_638_35272.n14 0.427167
R17600 a_638_35272.n0 a_638_35272.n15 0.427167
R17601 a_638_35272.n0 a_638_35272.n16 0.619389
R17602 a_638_35272.n16 a_638_35272.n17 0.427167
R17603 a_638_35272.n17 a_638_35272.n18 0.427167
R17604 a_638_35272.n18 a_638_35272.n19 0.427167
R17605 a_638_35272.n19 a_638_35272.n20 0.427167
R17606 a_638_35272.n20 a_638_35272.n21 0.427167
R17607 a_638_35272.n21 a_638_35272.n22 0.427167
R17608 a_638_35272.n22 a_638_35272.n23 0.427167
R17609 a_638_35272.n23 a_638_35272.n24 0.619389
R17610 a_638_35272.n24 a_638_35272.n25 0.427167
R17611 a_638_35272.n25 a_638_35272.n26 0.427167
R17612 a_638_35272.n26 a_638_35272.n27 0.427167
R17613 a_638_35272.n27 a_638_35272.n28 0.427167
R17614 a_638_35272.n28 a_638_35272.n29 0.427167
R17615 a_638_35272.n29 a_638_35272.n30 0.427167
R17616 a_638_35272.n30 a_638_35272.n31 0.427167
R17617 a_638_35272.n31 a_638_35272.n34 0.548278
R17618 a_638_35272.n34 a_638_35272.n70 0.227167
R17619 a_638_35272.n1 a_638_35272.n32 0.466493
R17620 a_638_35272.n36 a_638_35272.t19 7.71211
R17621 a_638_35272.n37 a_638_35272.t54 7.71211
R17622 a_638_35272.n38 a_638_35272.t26 7.71211
R17623 a_638_35272.n39 a_638_35272.t18 7.71211
R17624 a_638_35272.n40 a_638_35272.t31 7.71211
R17625 a_638_35272.n41 a_638_35272.t13 7.71211
R17626 a_638_35272.n42 a_638_35272.t45 7.71211
R17627 a_638_35272.n43 a_638_35272.t35 7.71211
R17628 a_638_35272.n44 a_638_35272.t61 7.71211
R17629 a_638_35272.n45 a_638_35272.t36 7.71211
R17630 a_638_35272.n46 a_638_35272.t55 7.71211
R17631 a_638_35272.n47 a_638_35272.t17 7.71211
R17632 a_638_35272.n48 a_638_35272.t64 7.71211
R17633 a_638_35272.n49 a_638_35272.t65 7.71211
R17634 a_638_35272.n50 a_638_35272.t41 7.71211
R17635 a_638_35272.n51 a_638_35272.t7 7.71211
R17636 a_638_35272.n52 a_638_35272.t22 7.71211
R17637 a_638_35272.n53 a_638_35272.t25 7.71211
R17638 a_638_35272.n54 a_638_35272.t42 7.71211
R17639 a_638_35272.n55 a_638_35272.t53 7.71211
R17640 a_638_35272.n56 a_638_35272.t20 7.71211
R17641 a_638_35272.n57 a_638_35272.t4 7.71211
R17642 a_638_35272.n58 a_638_35272.t66 7.71211
R17643 a_638_35272.n59 a_638_35272.t44 7.71211
R17644 a_638_35272.n60 a_638_35272.t9 7.71211
R17645 a_638_35272.n61 a_638_35272.t51 7.71211
R17646 a_638_35272.n62 a_638_35272.t27 7.71211
R17647 a_638_35272.n63 a_638_35272.t21 7.71211
R17648 a_638_35272.n64 a_638_35272.t28 7.71211
R17649 a_638_35272.n65 a_638_35272.t16 7.71211
R17650 a_638_35272.n66 a_638_35272.t10 7.71211
R17651 a_638_35272.n67 a_638_35272.t23 7.71211
R17652 a_638_35272.n32 a_638_35272.n36 0.69448
R17653 a_638_35272.n36 a_638_35272.n37 0.427167
R17654 a_638_35272.n37 a_638_35272.n38 0.427167
R17655 a_638_35272.n38 a_638_35272.n39 0.427167
R17656 a_638_35272.n39 a_638_35272.n40 0.427167
R17657 a_638_35272.n40 a_638_35272.n41 0.427167
R17658 a_638_35272.n41 a_638_35272.n42 0.427167
R17659 a_638_35272.n42 a_638_35272.n43 0.427167
R17660 a_638_35272.n43 a_638_35272.n44 0.619389
R17661 a_638_35272.n44 a_638_35272.n45 0.427167
R17662 a_638_35272.n45 a_638_35272.n46 0.427167
R17663 a_638_35272.n46 a_638_35272.n47 0.427167
R17664 a_638_35272.n47 a_638_35272.n48 0.427167
R17665 a_638_35272.n48 a_638_35272.n49 0.427167
R17666 a_638_35272.n49 a_638_35272.n50 0.427167
R17667 a_638_35272.n50 a_638_35272.n51 0.427167
R17668 a_638_35272.n51 a_638_35272.n52 0.619389
R17669 a_638_35272.n52 a_638_35272.n53 0.427167
R17670 a_638_35272.n53 a_638_35272.n54 0.427167
R17671 a_638_35272.n54 a_638_35272.n55 0.427167
R17672 a_638_35272.n55 a_638_35272.n56 0.427167
R17673 a_638_35272.n56 a_638_35272.n57 0.427167
R17674 a_638_35272.n57 a_638_35272.n58 0.427167
R17675 a_638_35272.n58 a_638_35272.n59 0.427167
R17676 a_638_35272.n59 a_638_35272.n60 0.619389
R17677 a_638_35272.n60 a_638_35272.n61 0.427167
R17678 a_638_35272.n61 a_638_35272.n62 0.427167
R17679 a_638_35272.n62 a_638_35272.n63 0.427167
R17680 a_638_35272.n64 a_638_35272.n63 0.427167
R17681 a_638_35272.n65 a_638_35272.n64 0.427167
R17682 a_638_35272.n66 a_638_35272.n65 0.427167
R17683 a_638_35272.n67 a_638_35272.n66 0.427167
R17684 a_638_35272.n35 a_638_35272.n67 0.334944
R17685 a_638_35272.n35 a_638_35272.n71 0.227167
R17686 a_638_35272.n70 a_638_35272.n72 4.96756
R17687 a_638_35272.n72 a_638_35272.n71 4.83019
R17688 a_638_35272.n72 a_638_35272.t2 0.113082
R17689 a_638_35272.n69 a_638_35272.n68 0.0655
R17690 a_638_35272.n69 a_638_35272.n71 4.60509
R17691 a_638_35272.n70 a_638_35272.n69 4.74618
R17692 a_638_35272.n68 a_638_35272.t58 0.0480817
R17693 a_638_35272.n68 a_638_35272.t59 0.0480817
R17694 a_638_35272.n33 a_638_35272.n35 4.60509
R17695 a_638_35272.n34 a_638_35272.n33 4.74618
R17696 a_638_35272.n33 a_638_35272.t3 0.113082
R17697 a_638_35272.n32 a_638_35272.t32 9.85476
R17698 a_1340_32660.t0 a_1340_32660.t1 7.42556
R17699 BIT_SEL[39].t1 BIT_SEL[39] 120.195
R17700 BIT_SEL[39] BIT_SEL[39].n0 9.23514
R17701 BIT_SEL[39] BIT_SEL[39].n0 3.39318
R17702 BIT_SEL[39] BIT_SEL[39].n1 9.23514
R17703 BIT_SEL[39].n1 BIT_SEL[39] 3.39318
R17704 BIT_SEL[39] BIT_SEL[39].n2 9.23514
R17705 BIT_SEL[39].n2 BIT_SEL[39] 3.39318
R17706 BIT_SEL[39] BIT_SEL[39].n3 9.23514
R17707 BIT_SEL[39].n3 BIT_SEL[39] 3.39318
R17708 BIT_SEL[39] BIT_SEL[39].n4 9.23514
R17709 BIT_SEL[39].n4 BIT_SEL[39] 3.39318
R17710 BIT_SEL[39] BIT_SEL[39].n5 9.23514
R17711 BIT_SEL[39].n5 BIT_SEL[39] 3.39318
R17712 BIT_SEL[39] BIT_SEL[39].n6 9.23514
R17713 BIT_SEL[39].n6 BIT_SEL[39] 3.39318
R17714 BIT_SEL[39].t2 BIT_SEL[39].n6 116.802
R17715 BIT_SEL[39].t4 BIT_SEL[39].n5 116.802
R17716 BIT_SEL[39].t0 BIT_SEL[39].n4 116.802
R17717 BIT_SEL[39].t6 BIT_SEL[39].n3 116.802
R17718 BIT_SEL[39].t5 BIT_SEL[39].n2 116.802
R17719 BIT_SEL[39].n1 BIT_SEL[39].t3 116.802
R17720 BIT_SEL[39].n0 BIT_SEL[39].t7 116.802
R17721 a_14320_41274.t0 a_14320_41274.t1 5.92075
R17722 a_638_43149.t0 a_638_43149.n0 7.71211
R17723 a_638_43149.n1 a_638_43149.t6 7.71211
R17724 a_638_43149.n2 a_638_43149.t20 7.71211
R17725 a_638_43149.n3 a_638_43149.t10 7.71211
R17726 a_638_43149.n4 a_638_43149.t60 7.71211
R17727 a_638_43149.n5 a_638_43149.t9 7.71211
R17728 a_638_43149.n6 a_638_43149.t26 7.71211
R17729 a_638_43149.n7 a_638_43149.t54 7.71211
R17730 a_638_43149.n8 a_638_43149.t1 7.71211
R17731 a_638_43149.n9 a_638_43149.t59 7.71211
R17732 a_638_43149.n10 a_638_43149.t62 7.71211
R17733 a_638_43149.n11 a_638_43149.t66 7.71211
R17734 a_638_43149.n12 a_638_43149.t63 7.71211
R17735 a_638_43149.n13 a_638_43149.t18 7.71211
R17736 a_638_43149.n14 a_638_43149.t65 7.71211
R17737 a_638_43149.n15 a_638_43149.t38 7.71211
R17738 a_638_43149.n16 a_638_43149.t15 7.71211
R17739 a_638_43149.n17 a_638_43149.t67 7.71211
R17740 a_638_43149.n18 a_638_43149.t61 7.71211
R17741 a_638_43149.n19 a_638_43149.t53 7.71211
R17742 a_638_43149.n20 a_638_43149.t22 7.71211
R17743 a_638_43149.n21 a_638_43149.t45 7.71211
R17744 a_638_43149.n22 a_638_43149.t46 7.71211
R17745 a_638_43149.n23 a_638_43149.t19 7.71211
R17746 a_638_43149.n24 a_638_43149.t34 7.71211
R17747 a_638_43149.n25 a_638_43149.t56 7.71211
R17748 a_638_43149.n26 a_638_43149.t44 7.71211
R17749 a_638_43149.n27 a_638_43149.t23 7.71211
R17750 a_638_43149.n28 a_638_43149.t21 7.71211
R17751 a_638_43149.n29 a_638_43149.t36 7.71211
R17752 a_638_43149.n30 a_638_43149.t57 7.71211
R17753 a_638_43149.n31 a_638_43149.t47 7.71211
R17754 a_638_43149.n2 a_638_43149.n1 0.427167
R17755 a_638_43149.n3 a_638_43149.n2 0.427167
R17756 a_638_43149.n4 a_638_43149.n3 0.427167
R17757 a_638_43149.n5 a_638_43149.n4 0.427167
R17758 a_638_43149.n6 a_638_43149.n5 0.427167
R17759 a_638_43149.n7 a_638_43149.n6 0.427167
R17760 a_638_43149.n8 a_638_43149.n7 0.427167
R17761 a_638_43149.n9 a_638_43149.n8 0.619389
R17762 a_638_43149.n10 a_638_43149.n9 0.427167
R17763 a_638_43149.n11 a_638_43149.n10 0.427167
R17764 a_638_43149.n12 a_638_43149.n11 0.427167
R17765 a_638_43149.n13 a_638_43149.n12 0.427167
R17766 a_638_43149.n14 a_638_43149.n13 0.427167
R17767 a_638_43149.n15 a_638_43149.n14 0.427167
R17768 a_638_43149.n16 a_638_43149.n15 0.427167
R17769 a_638_43149.n17 a_638_43149.n16 0.619389
R17770 a_638_43149.n18 a_638_43149.n17 0.427167
R17771 a_638_43149.n19 a_638_43149.n18 0.427167
R17772 a_638_43149.n20 a_638_43149.n19 0.427167
R17773 a_638_43149.n21 a_638_43149.n20 0.427167
R17774 a_638_43149.n22 a_638_43149.n21 0.427167
R17775 a_638_43149.n0 a_638_43149.n22 0.427167
R17776 a_638_43149.n0 a_638_43149.n23 0.427167
R17777 a_638_43149.n23 a_638_43149.n24 0.619389
R17778 a_638_43149.n24 a_638_43149.n25 0.427167
R17779 a_638_43149.n25 a_638_43149.n26 0.427167
R17780 a_638_43149.n26 a_638_43149.n27 0.427167
R17781 a_638_43149.n27 a_638_43149.n28 0.427167
R17782 a_638_43149.n28 a_638_43149.n29 0.427167
R17783 a_638_43149.n29 a_638_43149.n30 0.427167
R17784 a_638_43149.n30 a_638_43149.n31 0.427167
R17785 a_638_43149.n31 a_638_43149.n34 0.548278
R17786 a_638_43149.n34 a_638_43149.n70 0.227167
R17787 a_638_43149.n1 a_638_43149.n32 0.466493
R17788 a_638_43149.n36 a_638_43149.t4 7.71211
R17789 a_638_43149.n37 a_638_43149.t51 7.71211
R17790 a_638_43149.n38 a_638_43149.t39 7.71211
R17791 a_638_43149.n39 a_638_43149.t14 7.71211
R17792 a_638_43149.n40 a_638_43149.t5 7.71211
R17793 a_638_43149.n41 a_638_43149.t50 7.71211
R17794 a_638_43149.n42 a_638_43149.t12 7.71211
R17795 a_638_43149.n43 a_638_43149.t13 7.71211
R17796 a_638_43149.n44 a_638_43149.t16 7.71211
R17797 a_638_43149.n45 a_638_43149.t49 7.71211
R17798 a_638_43149.n46 a_638_43149.t40 7.71211
R17799 a_638_43149.n47 a_638_43149.t3 7.71211
R17800 a_638_43149.n48 a_638_43149.t31 7.71211
R17801 a_638_43149.n49 a_638_43149.t27 7.71211
R17802 a_638_43149.n50 a_638_43149.t41 7.71211
R17803 a_638_43149.n51 a_638_43149.t11 7.71211
R17804 a_638_43149.n52 a_638_43149.t52 7.71211
R17805 a_638_43149.n53 a_638_43149.t55 7.71211
R17806 a_638_43149.n54 a_638_43149.t8 7.71211
R17807 a_638_43149.n55 a_638_43149.t43 7.71211
R17808 a_638_43149.n56 a_638_43149.t29 7.71211
R17809 a_638_43149.n57 a_638_43149.t25 7.71211
R17810 a_638_43149.n58 a_638_43149.t48 7.71211
R17811 a_638_43149.n59 a_638_43149.t64 7.71211
R17812 a_638_43149.n60 a_638_43149.t7 7.71211
R17813 a_638_43149.n61 a_638_43149.t42 7.71211
R17814 a_638_43149.n62 a_638_43149.t2 7.71211
R17815 a_638_43149.n63 a_638_43149.t33 7.71211
R17816 a_638_43149.n64 a_638_43149.t17 7.71211
R17817 a_638_43149.n65 a_638_43149.t37 7.71211
R17818 a_638_43149.n66 a_638_43149.t58 7.71211
R17819 a_638_43149.n67 a_638_43149.t68 7.71211
R17820 a_638_43149.n32 a_638_43149.n36 0.69448
R17821 a_638_43149.n36 a_638_43149.n37 0.427167
R17822 a_638_43149.n37 a_638_43149.n38 0.427167
R17823 a_638_43149.n38 a_638_43149.n39 0.427167
R17824 a_638_43149.n39 a_638_43149.n40 0.427167
R17825 a_638_43149.n40 a_638_43149.n41 0.427167
R17826 a_638_43149.n41 a_638_43149.n42 0.427167
R17827 a_638_43149.n42 a_638_43149.n43 0.427167
R17828 a_638_43149.n43 a_638_43149.n44 0.619389
R17829 a_638_43149.n44 a_638_43149.n45 0.427167
R17830 a_638_43149.n45 a_638_43149.n46 0.427167
R17831 a_638_43149.n46 a_638_43149.n47 0.427167
R17832 a_638_43149.n47 a_638_43149.n48 0.427167
R17833 a_638_43149.n48 a_638_43149.n49 0.427167
R17834 a_638_43149.n49 a_638_43149.n50 0.427167
R17835 a_638_43149.n50 a_638_43149.n51 0.427167
R17836 a_638_43149.n51 a_638_43149.n52 0.619389
R17837 a_638_43149.n52 a_638_43149.n53 0.427167
R17838 a_638_43149.n53 a_638_43149.n54 0.427167
R17839 a_638_43149.n54 a_638_43149.n55 0.427167
R17840 a_638_43149.n55 a_638_43149.n56 0.427167
R17841 a_638_43149.n57 a_638_43149.n56 0.427167
R17842 a_638_43149.n58 a_638_43149.n57 0.427167
R17843 a_638_43149.n59 a_638_43149.n58 0.427167
R17844 a_638_43149.n60 a_638_43149.n59 0.619389
R17845 a_638_43149.n61 a_638_43149.n60 0.427167
R17846 a_638_43149.n62 a_638_43149.n61 0.427167
R17847 a_638_43149.n63 a_638_43149.n62 0.427167
R17848 a_638_43149.n64 a_638_43149.n63 0.427167
R17849 a_638_43149.n65 a_638_43149.n64 0.427167
R17850 a_638_43149.n66 a_638_43149.n65 0.427167
R17851 a_638_43149.n67 a_638_43149.n66 0.427167
R17852 a_638_43149.n35 a_638_43149.n67 0.334944
R17853 a_638_43149.n35 a_638_43149.n71 0.227167
R17854 a_638_43149.n70 a_638_43149.n72 4.96756
R17855 a_638_43149.n72 a_638_43149.n71 4.83019
R17856 a_638_43149.n72 a_638_43149.t32 0.113082
R17857 a_638_43149.n69 a_638_43149.n68 0.0655
R17858 a_638_43149.n69 a_638_43149.n71 4.60509
R17859 a_638_43149.n70 a_638_43149.n69 4.74618
R17860 a_638_43149.n68 a_638_43149.t24 0.0480817
R17861 a_638_43149.n68 a_638_43149.t35 0.0480817
R17862 a_638_43149.n33 a_638_43149.n35 4.60509
R17863 a_638_43149.n34 a_638_43149.n33 4.74618
R17864 a_638_43149.n33 a_638_43149.t28 0.113082
R17865 a_638_43149.n32 a_638_43149.t30 9.85476
R17866 a_1340_40906.t0 a_1340_40906.t1 6.39662
R17867 a_7738_27712.t0 a_7738_27712.t1 6.66648
R17868 BIT_SEL[11].n6 BIT_SEL[11] 4.57764
R17869 BIT_SEL[11] BIT_SEL[11].n6 8.05068
R17870 BIT_SEL[11] BIT_SEL[11].t2 122.203
R17871 BIT_SEL[11].n6 BIT_SEL[11].t0 117.626
R17872 BIT_SEL[11] BIT_SEL[11].n0 8.05068
R17873 BIT_SEL[11].n0 BIT_SEL[11] 4.57764
R17874 BIT_SEL[11] BIT_SEL[11].n1 8.05068
R17875 BIT_SEL[11].n1 BIT_SEL[11] 4.57764
R17876 BIT_SEL[11] BIT_SEL[11].n2 8.05068
R17877 BIT_SEL[11].n2 BIT_SEL[11] 4.57764
R17878 BIT_SEL[11] BIT_SEL[11].n3 8.05068
R17879 BIT_SEL[11].n3 BIT_SEL[11] 4.57764
R17880 BIT_SEL[11] BIT_SEL[11].n4 8.05068
R17881 BIT_SEL[11].n4 BIT_SEL[11] 4.57764
R17882 BIT_SEL[11] BIT_SEL[11].n5 8.05068
R17883 BIT_SEL[11].n5 BIT_SEL[11] 4.57764
R17884 BIT_SEL[11].t7 BIT_SEL[11].n5 117.626
R17885 BIT_SEL[11].t4 BIT_SEL[11].n4 117.626
R17886 BIT_SEL[11].t6 BIT_SEL[11].n3 117.626
R17887 BIT_SEL[11].t1 BIT_SEL[11].n2 117.626
R17888 BIT_SEL[11].t5 BIT_SEL[11].n1 117.626
R17889 BIT_SEL[11].t3 BIT_SEL[11].n0 117.626
R17890 a_1340_9029.t0 a_1340_9029.t1 7.42556
R17891 a_638_11641.t0 a_638_11641.n0 7.71211
R17892 a_638_11641.n2 a_638_11641.t29 7.71211
R17893 a_638_11641.n3 a_638_11641.t25 7.71211
R17894 a_638_11641.n4 a_638_11641.t50 7.71211
R17895 a_638_11641.n5 a_638_11641.t13 7.71211
R17896 a_638_11641.n6 a_638_11641.t37 7.71211
R17897 a_638_11641.n7 a_638_11641.t16 7.71211
R17898 a_638_11641.n8 a_638_11641.t52 7.71211
R17899 a_638_11641.n9 a_638_11641.t64 7.71211
R17900 a_638_11641.n10 a_638_11641.t56 7.71211
R17901 a_638_11641.n11 a_638_11641.t35 7.71211
R17902 a_638_11641.n12 a_638_11641.t28 7.71211
R17903 a_638_11641.n13 a_638_11641.t24 7.71211
R17904 a_638_11641.n14 a_638_11641.t33 7.71211
R17905 a_638_11641.n15 a_638_11641.t22 7.71211
R17906 a_638_11641.n16 a_638_11641.t57 7.71211
R17907 a_638_11641.n17 a_638_11641.t10 7.71211
R17908 a_638_11641.n18 a_638_11641.t27 7.71211
R17909 a_638_11641.n19 a_638_11641.t11 7.71211
R17910 a_638_11641.n20 a_638_11641.t7 7.71211
R17911 a_638_11641.n21 a_638_11641.t2 7.71211
R17912 a_638_11641.n22 a_638_11641.t44 7.71211
R17913 a_638_11641.n23 a_638_11641.t54 7.71211
R17914 a_638_11641.n24 a_638_11641.t59 7.71211
R17915 a_638_11641.n25 a_638_11641.t18 7.71211
R17916 a_638_11641.n26 a_638_11641.t12 7.71211
R17917 a_638_11641.n27 a_638_11641.t17 7.71211
R17918 a_638_11641.n28 a_638_11641.t51 7.71211
R17919 a_638_11641.n29 a_638_11641.t66 7.71211
R17920 a_638_11641.n30 a_638_11641.t48 7.71211
R17921 a_638_11641.n31 a_638_11641.t8 7.71211
R17922 a_638_11641.n32 a_638_11641.t41 7.71211
R17923 a_638_11641.n3 a_638_11641.n2 0.427167
R17924 a_638_11641.n4 a_638_11641.n3 0.427167
R17925 a_638_11641.n5 a_638_11641.n4 0.427167
R17926 a_638_11641.n6 a_638_11641.n5 0.427167
R17927 a_638_11641.n0 a_638_11641.n6 0.427167
R17928 a_638_11641.n0 a_638_11641.n7 0.427167
R17929 a_638_11641.n7 a_638_11641.n8 0.427167
R17930 a_638_11641.n8 a_638_11641.n9 0.619389
R17931 a_638_11641.n9 a_638_11641.n10 0.427167
R17932 a_638_11641.n10 a_638_11641.n11 0.427167
R17933 a_638_11641.n11 a_638_11641.n12 0.427167
R17934 a_638_11641.n12 a_638_11641.n13 0.427167
R17935 a_638_11641.n13 a_638_11641.n14 0.427167
R17936 a_638_11641.n14 a_638_11641.n15 0.427167
R17937 a_638_11641.n15 a_638_11641.n16 0.427167
R17938 a_638_11641.n16 a_638_11641.n17 0.619389
R17939 a_638_11641.n17 a_638_11641.n18 0.427167
R17940 a_638_11641.n18 a_638_11641.n19 0.427167
R17941 a_638_11641.n19 a_638_11641.n20 0.427167
R17942 a_638_11641.n20 a_638_11641.n21 0.427167
R17943 a_638_11641.n21 a_638_11641.n22 0.427167
R17944 a_638_11641.n22 a_638_11641.n23 0.427167
R17945 a_638_11641.n23 a_638_11641.n24 0.427167
R17946 a_638_11641.n24 a_638_11641.n25 0.619389
R17947 a_638_11641.n25 a_638_11641.n26 0.427167
R17948 a_638_11641.n26 a_638_11641.n27 0.427167
R17949 a_638_11641.n27 a_638_11641.n28 0.427167
R17950 a_638_11641.n28 a_638_11641.n29 0.427167
R17951 a_638_11641.n29 a_638_11641.n30 0.427167
R17952 a_638_11641.n30 a_638_11641.n31 0.427167
R17953 a_638_11641.n31 a_638_11641.n32 0.427167
R17954 a_638_11641.n32 a_638_11641.n1 0.334944
R17955 a_638_11641.n1 a_638_11641.n33 0.227167
R17956 a_638_11641.n34 a_638_11641.n35 0.466493
R17957 a_638_11641.n2 a_638_11641.n34 0.69448
R17958 a_638_11641.n35 a_638_11641.t1 7.71211
R17959 a_638_11641.n36 a_638_11641.t42 7.71211
R17960 a_638_11641.n37 a_638_11641.t23 7.71211
R17961 a_638_11641.n38 a_638_11641.t63 7.71211
R17962 a_638_11641.n39 a_638_11641.t65 7.71211
R17963 a_638_11641.n40 a_638_11641.t53 7.71211
R17964 a_638_11641.n41 a_638_11641.t55 7.71211
R17965 a_638_11641.n42 a_638_11641.t30 7.71211
R17966 a_638_11641.n43 a_638_11641.t40 7.71211
R17967 a_638_11641.n44 a_638_11641.t19 7.71211
R17968 a_638_11641.n45 a_638_11641.t36 7.71211
R17969 a_638_11641.n46 a_638_11641.t9 7.71211
R17970 a_638_11641.n47 a_638_11641.t5 7.71211
R17971 a_638_11641.n48 a_638_11641.t4 7.71211
R17972 a_638_11641.n49 a_638_11641.t46 7.71211
R17973 a_638_11641.n50 a_638_11641.t14 7.71211
R17974 a_638_11641.n51 a_638_11641.t39 7.71211
R17975 a_638_11641.n52 a_638_11641.t3 7.71211
R17976 a_638_11641.n53 a_638_11641.t58 7.71211
R17977 a_638_11641.n54 a_638_11641.t60 7.71211
R17978 a_638_11641.n55 a_638_11641.t45 7.71211
R17979 a_638_11641.n56 a_638_11641.t43 7.71211
R17980 a_638_11641.n57 a_638_11641.t6 7.71211
R17981 a_638_11641.n58 a_638_11641.t31 7.71211
R17982 a_638_11641.n59 a_638_11641.t47 7.71211
R17983 a_638_11641.n60 a_638_11641.t38 7.71211
R17984 a_638_11641.n61 a_638_11641.t32 7.71211
R17985 a_638_11641.n62 a_638_11641.t62 7.71211
R17986 a_638_11641.n63 a_638_11641.t15 7.71211
R17987 a_638_11641.n64 a_638_11641.t61 7.71211
R17988 a_638_11641.n65 a_638_11641.t49 7.71211
R17989 a_638_11641.n66 a_638_11641.t34 7.71211
R17990 a_638_11641.n35 a_638_11641.n36 0.427167
R17991 a_638_11641.n36 a_638_11641.n37 0.427167
R17992 a_638_11641.n37 a_638_11641.n38 0.427167
R17993 a_638_11641.n38 a_638_11641.n39 0.427167
R17994 a_638_11641.n39 a_638_11641.n40 0.427167
R17995 a_638_11641.n40 a_638_11641.n41 0.427167
R17996 a_638_11641.n41 a_638_11641.n42 0.427167
R17997 a_638_11641.n42 a_638_11641.n43 0.619389
R17998 a_638_11641.n43 a_638_11641.n44 0.427167
R17999 a_638_11641.n44 a_638_11641.n45 0.427167
R18000 a_638_11641.n45 a_638_11641.n46 0.427167
R18001 a_638_11641.n46 a_638_11641.n47 0.427167
R18002 a_638_11641.n47 a_638_11641.n48 0.427167
R18003 a_638_11641.n48 a_638_11641.n49 0.427167
R18004 a_638_11641.n49 a_638_11641.n50 0.427167
R18005 a_638_11641.n50 a_638_11641.n51 0.619389
R18006 a_638_11641.n51 a_638_11641.n52 0.427167
R18007 a_638_11641.n52 a_638_11641.n53 0.427167
R18008 a_638_11641.n53 a_638_11641.n54 0.427167
R18009 a_638_11641.n54 a_638_11641.n55 0.427167
R18010 a_638_11641.n55 a_638_11641.n56 0.427167
R18011 a_638_11641.n56 a_638_11641.n57 0.427167
R18012 a_638_11641.n57 a_638_11641.n58 0.427167
R18013 a_638_11641.n58 a_638_11641.n59 0.619389
R18014 a_638_11641.n59 a_638_11641.n60 0.427167
R18015 a_638_11641.n60 a_638_11641.n61 0.427167
R18016 a_638_11641.n61 a_638_11641.n62 0.427167
R18017 a_638_11641.n62 a_638_11641.n63 0.427167
R18018 a_638_11641.n63 a_638_11641.n64 0.427167
R18019 a_638_11641.n64 a_638_11641.n65 0.427167
R18020 a_638_11641.n65 a_638_11641.n66 0.427167
R18021 a_638_11641.n66 a_638_11641.n71 0.548278
R18022 a_638_11641.n71 a_638_11641.n68 0.227167
R18023 a_638_11641.n71 a_638_11641.n72 4.74618
R18024 a_638_11641.n1 a_638_11641.n72 4.60509
R18025 a_638_11641.n72 a_638_11641.t20 0.113082
R18026 a_638_11641.n70 a_638_11641.n69 0.0655
R18027 a_638_11641.n68 a_638_11641.n70 4.74618
R18028 a_638_11641.n33 a_638_11641.n70 4.60509
R18029 a_638_11641.n69 a_638_11641.t68 0.0480817
R18030 a_638_11641.n69 a_638_11641.t21 0.0480817
R18031 a_638_11641.n68 a_638_11641.n67 4.96756
R18032 a_638_11641.n33 a_638_11641.n67 4.83019
R18033 a_638_11641.n67 a_638_11641.t67 0.113082
R18034 a_638_11641.n34 a_638_11641.t26 9.85476
R18035 a_20810_9398.t0 a_20810_9398.t1 6.39548
R18036 a_154_29353.t0 a_154_29353.t1 13.9628
R18037 a_110_29441.t0 a_110_29441.t1 19.5535
R18038 BIT_SEL[25].n6 BIT_SEL[25] 3.98461
R18039 BIT_SEL[25] BIT_SEL[25].n6 8.64371
R18040 BIT_SEL[25] BIT_SEL[25].t3 121.198
R18041 BIT_SEL[25].n6 BIT_SEL[25].t1 117.215
R18042 BIT_SEL[25] BIT_SEL[25].n0 8.64371
R18043 BIT_SEL[25].n0 BIT_SEL[25] 3.98461
R18044 BIT_SEL[25] BIT_SEL[25].n1 8.64371
R18045 BIT_SEL[25].n1 BIT_SEL[25] 3.98461
R18046 BIT_SEL[25] BIT_SEL[25].n2 8.64371
R18047 BIT_SEL[25].n2 BIT_SEL[25] 3.98461
R18048 BIT_SEL[25] BIT_SEL[25].n3 8.64371
R18049 BIT_SEL[25].n3 BIT_SEL[25] 3.98461
R18050 BIT_SEL[25] BIT_SEL[25].n4 8.64371
R18051 BIT_SEL[25].n4 BIT_SEL[25] 3.98461
R18052 BIT_SEL[25] BIT_SEL[25].n5 8.64371
R18053 BIT_SEL[25].n5 BIT_SEL[25] 3.98461
R18054 BIT_SEL[25].t7 BIT_SEL[25].n5 117.215
R18055 BIT_SEL[25].t5 BIT_SEL[25].n4 117.215
R18056 BIT_SEL[25].t2 BIT_SEL[25].n3 117.215
R18057 BIT_SEL[25].t4 BIT_SEL[25].n2 117.215
R18058 BIT_SEL[25].t0 BIT_SEL[25].n1 117.215
R18059 BIT_SEL[25].t6 BIT_SEL[25].n0 117.215
R18060 a_7830_25152.t0 a_7830_25152.t1 6.39548
R18061 a_110_6258.t0 a_110_6258.t1 19.5535
R18062 a_154_6170.t0 a_154_6170.t1 13.9628
R18063 a_110_61397.t0 a_110_61397.t1 19.5535
R18064 a_154_61309.t0 a_154_61309.t1 13.9628
R18065 a_110_49568.t0 a_110_49568.n0 8.34715
R18066 a_110_49568.n0 a_110_49568.n3 0.1805
R18067 a_110_49568.n3 a_110_49568.n2 4.47779
R18068 a_110_49568.n2 a_110_49568.t3 12.3497
R18069 a_110_49568.n2 a_110_49568.t5 17.192
R18070 a_110_49568.n0 a_110_49568.n1 14.1624
R18071 a_110_49568.n1 a_110_49568.t4 12.3497
R18072 a_110_49568.n1 a_110_49568.t2 17.192
R18073 a_110_49568.n3 a_110_49568.t1 4.44412
R18074 OUT[6] OUT[6].n0 9.0005
R18075 OUT[6].n0 OUT[6].t1 8.56064
R18076 OUT[6].n0 OUT[6].t0 4.38216
R18077 a_7738_43466.t0 a_7738_43466.t1 6.66648
R18078 BIT_SEL[52] BIT_SEL[52].n0 2.54461
R18079 BIT_SEL[52] BIT_SEL[52].n0 10.0837
R18080 BIT_SEL[52] BIT_SEL[52].n1 2.54461
R18081 BIT_SEL[52].n1 BIT_SEL[52] 10.0837
R18082 BIT_SEL[52] BIT_SEL[52].n2 2.54461
R18083 BIT_SEL[52].n2 BIT_SEL[52] 10.0837
R18084 BIT_SEL[52] BIT_SEL[52].n3 2.54461
R18085 BIT_SEL[52].n3 BIT_SEL[52] 10.0837
R18086 BIT_SEL[52] BIT_SEL[52].n4 2.54461
R18087 BIT_SEL[52].n4 BIT_SEL[52] 10.0837
R18088 BIT_SEL[52] BIT_SEL[52].n5 2.54461
R18089 BIT_SEL[52].n5 BIT_SEL[52] 10.0837
R18090 BIT_SEL[52] BIT_SEL[52].n6 2.54461
R18091 BIT_SEL[52].n6 BIT_SEL[52] 10.0837
R18092 BIT_SEL[52].t3 BIT_SEL[52] 118.73
R18093 BIT_SEL[52].t1 BIT_SEL[52].n6 116.186
R18094 BIT_SEL[52].t7 BIT_SEL[52].n5 116.186
R18095 BIT_SEL[52].t0 BIT_SEL[52].n4 116.186
R18096 BIT_SEL[52].t5 BIT_SEL[52].n3 116.186
R18097 BIT_SEL[52].t2 BIT_SEL[52].n2 116.186
R18098 BIT_SEL[52].n1 BIT_SEL[52].t4 116.186
R18099 BIT_SEL[52].n0 BIT_SEL[52].t6 116.186
R18100 a_20810_36903.t0 a_20810_36903.t1 7.18213
R18101 a_1340_11031.t0 a_1340_11031.t1 6.02155
R18102 a_154_16100.t0 a_154_16100.t1 13.9628
R18103 a_110_16188.t0 a_110_16188.t1 19.5535
R18104 a_20810_52289.t0 a_20810_52289.t1 8.02269
R18105 BIT_SEL[38] BIT_SEL[38].n0 3.39479
R18106 BIT_SEL[38] BIT_SEL[38].n0 9.23354
R18107 BIT_SEL[38] BIT_SEL[38].n1 3.39479
R18108 BIT_SEL[38].n1 BIT_SEL[38] 9.23354
R18109 BIT_SEL[38] BIT_SEL[38].n2 3.39479
R18110 BIT_SEL[38].n2 BIT_SEL[38] 9.23354
R18111 BIT_SEL[38] BIT_SEL[38].n3 3.39479
R18112 BIT_SEL[38].n3 BIT_SEL[38] 9.23354
R18113 BIT_SEL[38] BIT_SEL[38].n4 3.39479
R18114 BIT_SEL[38].n4 BIT_SEL[38] 9.23354
R18115 BIT_SEL[38] BIT_SEL[38].n5 3.39479
R18116 BIT_SEL[38].n5 BIT_SEL[38] 9.23354
R18117 BIT_SEL[38] BIT_SEL[38].n6 3.39479
R18118 BIT_SEL[38].n6 BIT_SEL[38] 9.23354
R18119 BIT_SEL[38].t4 BIT_SEL[38] 119.992
R18120 BIT_SEL[38].t3 BIT_SEL[38].n6 116.597
R18121 BIT_SEL[38].t1 BIT_SEL[38].n5 116.597
R18122 BIT_SEL[38].t7 BIT_SEL[38].n4 116.597
R18123 BIT_SEL[38].t6 BIT_SEL[38].n3 116.597
R18124 BIT_SEL[38].t2 BIT_SEL[38].n2 116.597
R18125 BIT_SEL[38].n1 BIT_SEL[38].t0 116.597
R18126 BIT_SEL[38].n0 BIT_SEL[38].t5 116.597
R18127 a_14320_13801.t0 a_14320_13801.t1 6.38524
R18128 a_20810_25152.t0 a_20810_25152.t1 6.39662
R18129 BIT_SEL[23].n6 BIT_SEL[23] 3.39318
R18130 BIT_SEL[23] BIT_SEL[23].n6 9.23514
R18131 BIT_SEL[23] BIT_SEL[23].t4 120.195
R18132 BIT_SEL[23].n6 BIT_SEL[23].t2 116.802
R18133 BIT_SEL[23] BIT_SEL[23].n0 9.23514
R18134 BIT_SEL[23].n0 BIT_SEL[23] 3.39318
R18135 BIT_SEL[23] BIT_SEL[23].n1 9.23514
R18136 BIT_SEL[23].n1 BIT_SEL[23] 3.39318
R18137 BIT_SEL[23] BIT_SEL[23].n2 9.23514
R18138 BIT_SEL[23].n2 BIT_SEL[23] 3.39318
R18139 BIT_SEL[23] BIT_SEL[23].n3 9.23514
R18140 BIT_SEL[23].n3 BIT_SEL[23] 3.39318
R18141 BIT_SEL[23] BIT_SEL[23].n4 9.23514
R18142 BIT_SEL[23].n4 BIT_SEL[23] 3.39318
R18143 BIT_SEL[23] BIT_SEL[23].n5 9.23514
R18144 BIT_SEL[23].n5 BIT_SEL[23] 3.39318
R18145 BIT_SEL[23].t5 BIT_SEL[23].n5 116.802
R18146 BIT_SEL[23].t7 BIT_SEL[23].n4 116.802
R18147 BIT_SEL[23].t3 BIT_SEL[23].n3 116.802
R18148 BIT_SEL[23].t1 BIT_SEL[23].n2 116.802
R18149 BIT_SEL[23].t0 BIT_SEL[23].n1 116.802
R18150 BIT_SEL[23].t6 BIT_SEL[23].n0 116.802
R18151 a_7830_25520.t0 a_7830_25520.t1 5.92075
R18152 a_20810_7557.t0 a_20810_7557.t1 9.05337
R18153 a_638_3764.t0 a_638_3764.n0 7.71211
R18154 a_638_3764.n1 a_638_3764.t64 7.71211
R18155 a_638_3764.n2 a_638_3764.t32 7.71211
R18156 a_638_3764.n3 a_638_3764.t23 7.71211
R18157 a_638_3764.n4 a_638_3764.t19 7.71211
R18158 a_638_3764.n5 a_638_3764.t38 7.71211
R18159 a_638_3764.n6 a_638_3764.t42 7.71211
R18160 a_638_3764.n7 a_638_3764.t55 7.71211
R18161 a_638_3764.n8 a_638_3764.t28 7.71211
R18162 a_638_3764.n9 a_638_3764.t61 7.71211
R18163 a_638_3764.n10 a_638_3764.t35 7.71211
R18164 a_638_3764.n11 a_638_3764.t26 7.71211
R18165 a_638_3764.n12 a_638_3764.t41 7.71211
R18166 a_638_3764.n13 a_638_3764.t16 7.71211
R18167 a_638_3764.n14 a_638_3764.t11 7.71211
R18168 a_638_3764.n15 a_638_3764.t68 7.71211
R18169 a_638_3764.n16 a_638_3764.t15 7.71211
R18170 a_638_3764.n17 a_638_3764.t53 7.71211
R18171 a_638_3764.n18 a_638_3764.t62 7.71211
R18172 a_638_3764.n19 a_638_3764.t18 7.71211
R18173 a_638_3764.n20 a_638_3764.t51 7.71211
R18174 a_638_3764.n21 a_638_3764.t31 7.71211
R18175 a_638_3764.n22 a_638_3764.t58 7.71211
R18176 a_638_3764.n23 a_638_3764.t2 7.71211
R18177 a_638_3764.n24 a_638_3764.t54 7.71211
R18178 a_638_3764.n25 a_638_3764.t30 7.71211
R18179 a_638_3764.n26 a_638_3764.t59 7.71211
R18180 a_638_3764.n27 a_638_3764.t1 7.71211
R18181 a_638_3764.n28 a_638_3764.t52 7.71211
R18182 a_638_3764.n29 a_638_3764.t14 7.71211
R18183 a_638_3764.n30 a_638_3764.t4 7.71211
R18184 a_638_3764.n31 a_638_3764.t57 7.71211
R18185 a_638_3764.n2 a_638_3764.n1 0.427167
R18186 a_638_3764.n3 a_638_3764.n2 0.427167
R18187 a_638_3764.n4 a_638_3764.n3 0.427167
R18188 a_638_3764.n5 a_638_3764.n4 0.427167
R18189 a_638_3764.n6 a_638_3764.n5 0.427167
R18190 a_638_3764.n7 a_638_3764.n6 0.427167
R18191 a_638_3764.n8 a_638_3764.n7 0.427167
R18192 a_638_3764.n9 a_638_3764.n8 0.619389
R18193 a_638_3764.n10 a_638_3764.n9 0.427167
R18194 a_638_3764.n11 a_638_3764.n10 0.427167
R18195 a_638_3764.n12 a_638_3764.n11 0.427167
R18196 a_638_3764.n13 a_638_3764.n12 0.427167
R18197 a_638_3764.n14 a_638_3764.n13 0.427167
R18198 a_638_3764.n15 a_638_3764.n14 0.427167
R18199 a_638_3764.n16 a_638_3764.n15 0.427167
R18200 a_638_3764.n0 a_638_3764.n16 0.619389
R18201 a_638_3764.n0 a_638_3764.n17 0.427167
R18202 a_638_3764.n17 a_638_3764.n18 0.427167
R18203 a_638_3764.n18 a_638_3764.n19 0.427167
R18204 a_638_3764.n19 a_638_3764.n20 0.427167
R18205 a_638_3764.n20 a_638_3764.n21 0.427167
R18206 a_638_3764.n21 a_638_3764.n22 0.427167
R18207 a_638_3764.n22 a_638_3764.n23 0.427167
R18208 a_638_3764.n23 a_638_3764.n24 0.619389
R18209 a_638_3764.n24 a_638_3764.n25 0.427167
R18210 a_638_3764.n25 a_638_3764.n26 0.427167
R18211 a_638_3764.n26 a_638_3764.n27 0.427167
R18212 a_638_3764.n27 a_638_3764.n28 0.427167
R18213 a_638_3764.n28 a_638_3764.n29 0.427167
R18214 a_638_3764.n29 a_638_3764.n30 0.427167
R18215 a_638_3764.n30 a_638_3764.n31 0.427167
R18216 a_638_3764.n31 a_638_3764.n34 0.548278
R18217 a_638_3764.n34 a_638_3764.n70 0.227167
R18218 a_638_3764.n1 a_638_3764.n32 0.466493
R18219 a_638_3764.n36 a_638_3764.t40 7.71211
R18220 a_638_3764.n37 a_638_3764.t13 7.71211
R18221 a_638_3764.n38 a_638_3764.t12 7.71211
R18222 a_638_3764.n39 a_638_3764.t9 7.71211
R18223 a_638_3764.n40 a_638_3764.t48 7.71211
R18224 a_638_3764.n41 a_638_3764.t60 7.71211
R18225 a_638_3764.n42 a_638_3764.t10 7.71211
R18226 a_638_3764.n43 a_638_3764.t36 7.71211
R18227 a_638_3764.n44 a_638_3764.t49 7.71211
R18228 a_638_3764.n45 a_638_3764.t25 7.71211
R18229 a_638_3764.n46 a_638_3764.t50 7.71211
R18230 a_638_3764.n47 a_638_3764.t44 7.71211
R18231 a_638_3764.n48 a_638_3764.t17 7.71211
R18232 a_638_3764.n49 a_638_3764.t66 7.71211
R18233 a_638_3764.n50 a_638_3764.t22 7.71211
R18234 a_638_3764.n51 a_638_3764.t8 7.71211
R18235 a_638_3764.n52 a_638_3764.t43 7.71211
R18236 a_638_3764.n53 a_638_3764.t63 7.71211
R18237 a_638_3764.n54 a_638_3764.t34 7.71211
R18238 a_638_3764.n55 a_638_3764.t24 7.71211
R18239 a_638_3764.n56 a_638_3764.t56 7.71211
R18240 a_638_3764.n57 a_638_3764.t46 7.71211
R18241 a_638_3764.n58 a_638_3764.t3 7.71211
R18242 a_638_3764.n59 a_638_3764.t21 7.71211
R18243 a_638_3764.n60 a_638_3764.t45 7.71211
R18244 a_638_3764.n61 a_638_3764.t65 7.71211
R18245 a_638_3764.n62 a_638_3764.t47 7.71211
R18246 a_638_3764.n63 a_638_3764.t39 7.71211
R18247 a_638_3764.n64 a_638_3764.t67 7.71211
R18248 a_638_3764.n65 a_638_3764.t37 7.71211
R18249 a_638_3764.n66 a_638_3764.t20 7.71211
R18250 a_638_3764.n67 a_638_3764.t27 7.71211
R18251 a_638_3764.n32 a_638_3764.n36 0.69448
R18252 a_638_3764.n36 a_638_3764.n37 0.427167
R18253 a_638_3764.n37 a_638_3764.n38 0.427167
R18254 a_638_3764.n38 a_638_3764.n39 0.427167
R18255 a_638_3764.n39 a_638_3764.n40 0.427167
R18256 a_638_3764.n40 a_638_3764.n41 0.427167
R18257 a_638_3764.n41 a_638_3764.n42 0.427167
R18258 a_638_3764.n42 a_638_3764.n43 0.427167
R18259 a_638_3764.n43 a_638_3764.n44 0.619389
R18260 a_638_3764.n44 a_638_3764.n45 0.427167
R18261 a_638_3764.n45 a_638_3764.n46 0.427167
R18262 a_638_3764.n46 a_638_3764.n47 0.427167
R18263 a_638_3764.n47 a_638_3764.n48 0.427167
R18264 a_638_3764.n48 a_638_3764.n49 0.427167
R18265 a_638_3764.n49 a_638_3764.n50 0.427167
R18266 a_638_3764.n50 a_638_3764.n51 0.427167
R18267 a_638_3764.n51 a_638_3764.n52 0.619389
R18268 a_638_3764.n52 a_638_3764.n53 0.427167
R18269 a_638_3764.n53 a_638_3764.n54 0.427167
R18270 a_638_3764.n54 a_638_3764.n55 0.427167
R18271 a_638_3764.n55 a_638_3764.n56 0.427167
R18272 a_638_3764.n56 a_638_3764.n57 0.427167
R18273 a_638_3764.n57 a_638_3764.n58 0.427167
R18274 a_638_3764.n58 a_638_3764.n59 0.427167
R18275 a_638_3764.n59 a_638_3764.n60 0.619389
R18276 a_638_3764.n60 a_638_3764.n61 0.427167
R18277 a_638_3764.n62 a_638_3764.n61 0.427167
R18278 a_638_3764.n63 a_638_3764.n62 0.427167
R18279 a_638_3764.n64 a_638_3764.n63 0.427167
R18280 a_638_3764.n65 a_638_3764.n64 0.427167
R18281 a_638_3764.n66 a_638_3764.n65 0.427167
R18282 a_638_3764.n67 a_638_3764.n66 0.427167
R18283 a_638_3764.n35 a_638_3764.n67 0.334944
R18284 a_638_3764.n35 a_638_3764.n71 0.227167
R18285 a_638_3764.n70 a_638_3764.n72 4.96756
R18286 a_638_3764.n72 a_638_3764.n71 4.83019
R18287 a_638_3764.n72 a_638_3764.t6 0.113082
R18288 a_638_3764.n69 a_638_3764.n68 0.0655
R18289 a_638_3764.n69 a_638_3764.n71 4.60509
R18290 a_638_3764.n70 a_638_3764.n69 4.74618
R18291 a_638_3764.n68 a_638_3764.t7 0.0480817
R18292 a_638_3764.n68 a_638_3764.t29 0.0480817
R18293 a_638_3764.n33 a_638_3764.n35 4.60509
R18294 a_638_3764.n34 a_638_3764.n33 4.74618
R18295 a_638_3764.n33 a_638_3764.t5 0.113082
R18296 a_638_3764.n32 a_638_3764.t33 9.85476
R18297 a_110_434.t0 a_110_434.t1 19.5535
R18298 a_154_346.t0 a_154_346.t1 13.9628
R18299 a_14320_62328.t0 a_14320_62328.t1 8.02468
R18300 BIT_SEL[54].n6 BIT_SEL[54] 9.23354
R18301 BIT_SEL[54] BIT_SEL[54].n6 3.39479
R18302 BIT_SEL[54].n6 BIT_SEL[54].t6 116.597
R18303 BIT_SEL[54] BIT_SEL[54].n0 3.39479
R18304 BIT_SEL[54].n0 BIT_SEL[54] 9.23354
R18305 BIT_SEL[54] BIT_SEL[54].n1 3.39479
R18306 BIT_SEL[54].n1 BIT_SEL[54] 9.23354
R18307 BIT_SEL[54] BIT_SEL[54].n2 3.39479
R18308 BIT_SEL[54].n2 BIT_SEL[54] 9.23354
R18309 BIT_SEL[54] BIT_SEL[54].n3 3.39479
R18310 BIT_SEL[54].n3 BIT_SEL[54] 9.23354
R18311 BIT_SEL[54] BIT_SEL[54].n4 3.39479
R18312 BIT_SEL[54].n4 BIT_SEL[54] 9.23354
R18313 BIT_SEL[54] BIT_SEL[54].n5 3.39479
R18314 BIT_SEL[54].n5 BIT_SEL[54] 9.23354
R18315 BIT_SEL[54].t5 BIT_SEL[54] 119.992
R18316 BIT_SEL[54].t4 BIT_SEL[54].n5 116.597
R18317 BIT_SEL[54].t2 BIT_SEL[54].n4 116.597
R18318 BIT_SEL[54].t0 BIT_SEL[54].n3 116.597
R18319 BIT_SEL[54].t7 BIT_SEL[54].n2 116.597
R18320 BIT_SEL[54].t3 BIT_SEL[54].n1 116.597
R18321 BIT_SEL[54].t1 BIT_SEL[54].n0 116.597
R18322 a_20810_37432.t0 a_20810_37432.t1 6.38524
R18323 a_110_34710.t0 a_110_34710.n4 4.88081
R18324 a_110_34710.n4 a_110_34710.n5 2.6905
R18325 a_110_34710.n5 a_110_34710.t2 2.06607
R18326 a_110_34710.n5 a_110_34710.t1 2.2382
R18327 a_110_34710.n4 a_110_34710.n0 0.766047
R18328 a_110_34710.n0 a_110_34710.t5 8.68401
R18329 a_110_34710.n2 a_110_34710.n3 5.21793
R18330 a_110_34710.n0 a_110_34710.n2 4.76793
R18331 a_110_34710.n3 a_110_34710.t3 8.51897
R18332 a_110_34710.n3 a_110_34710.t4 4.4523
R18333 a_110_34710.n2 a_110_34710.n1 8.53373
R18334 a_110_34710.n1 a_110_34710.t6 12.3497
R18335 a_110_34710.n1 a_110_34710.t7 17.192
R18336 a_110_33814.t0 a_110_33814.n3 4.44412
R18337 a_110_33814.n3 a_110_33814.n0 0.1805
R18338 a_110_33814.n3 a_110_33814.n2 4.47779
R18339 a_110_33814.n2 a_110_33814.t4 12.3497
R18340 a_110_33814.n2 a_110_33814.t5 17.192
R18341 a_110_33814.n0 a_110_33814.n1 14.1624
R18342 a_110_33814.n1 a_110_33814.t2 12.3497
R18343 a_110_33814.n1 a_110_33814.t3 17.192
R18344 a_110_33814.n0 a_110_33814.t1 8.34715
R18345 a_20810_52657.t0 a_20810_52657.t1 7.18213
R18346 a_1248_59220.t0 a_1248_59220.t1 6.66648
R18347 a_1340_26785.t0 a_1340_26785.t1 6.02155
R18348 a_1340_7557.t0 a_1340_7557.t1 9.05295
R18349 a_20810_40906.t0 a_20810_40906.t1 6.39662
R18350 BIT_SEL[57].n6 BIT_SEL[57] 3.98461
R18351 BIT_SEL[57] BIT_SEL[57].n6 8.64371
R18352 BIT_SEL[57] BIT_SEL[57].t5 121.198
R18353 BIT_SEL[57].n6 BIT_SEL[57].t1 117.215
R18354 BIT_SEL[57] BIT_SEL[57].n0 8.64371
R18355 BIT_SEL[57].n0 BIT_SEL[57] 3.98461
R18356 BIT_SEL[57] BIT_SEL[57].n1 8.64371
R18357 BIT_SEL[57].n1 BIT_SEL[57] 3.98461
R18358 BIT_SEL[57] BIT_SEL[57].n2 8.64371
R18359 BIT_SEL[57].n2 BIT_SEL[57] 3.98461
R18360 BIT_SEL[57] BIT_SEL[57].n3 8.64371
R18361 BIT_SEL[57].n3 BIT_SEL[57] 3.98461
R18362 BIT_SEL[57] BIT_SEL[57].n4 8.64371
R18363 BIT_SEL[57].n4 BIT_SEL[57] 3.98461
R18364 BIT_SEL[57] BIT_SEL[57].n5 8.64371
R18365 BIT_SEL[57].n5 BIT_SEL[57] 3.98461
R18366 BIT_SEL[57].t6 BIT_SEL[57].n5 117.215
R18367 BIT_SEL[57].t3 BIT_SEL[57].n4 117.215
R18368 BIT_SEL[57].t0 BIT_SEL[57].n3 117.215
R18369 BIT_SEL[57].t2 BIT_SEL[57].n2 117.215
R18370 BIT_SEL[57].t7 BIT_SEL[57].n1 117.215
R18371 BIT_SEL[57].t4 BIT_SEL[57].n0 117.215
R18372 BIT_SEL[60].n6 BIT_SEL[60] 7.2005
R18373 BIT_SEL[60] BIT_SEL[60].n6 5.42782
R18374 BIT_SEL[60].n6 BIT_SEL[60].t0 117.832
R18375 BIT_SEL[60] BIT_SEL[60].n0 5.42782
R18376 BIT_SEL[60].n0 BIT_SEL[60] 7.2005
R18377 BIT_SEL[60] BIT_SEL[60].n1 5.42782
R18378 BIT_SEL[60].n1 BIT_SEL[60] 7.2005
R18379 BIT_SEL[60] BIT_SEL[60].n2 5.42782
R18380 BIT_SEL[60].n2 BIT_SEL[60] 7.2005
R18381 BIT_SEL[60] BIT_SEL[60].n3 5.42782
R18382 BIT_SEL[60].n3 BIT_SEL[60] 7.2005
R18383 BIT_SEL[60] BIT_SEL[60].n4 5.42782
R18384 BIT_SEL[60].n4 BIT_SEL[60] 7.2005
R18385 BIT_SEL[60] BIT_SEL[60].n5 5.42782
R18386 BIT_SEL[60].n5 BIT_SEL[60] 7.2005
R18387 BIT_SEL[60].t5 BIT_SEL[60] 123.258
R18388 BIT_SEL[60].t2 BIT_SEL[60].n5 117.832
R18389 BIT_SEL[60].t4 BIT_SEL[60].n4 117.832
R18390 BIT_SEL[60].t1 BIT_SEL[60].n3 117.832
R18391 BIT_SEL[60].t3 BIT_SEL[60].n2 117.832
R18392 BIT_SEL[60].t7 BIT_SEL[60].n1 117.832
R18393 BIT_SEL[60].t6 BIT_SEL[60].n0 117.832
R18394 a_20810_7189.t0 a_20810_7189.t1 8.02427
R18395 a_20810_55763.t0 a_20810_55763.t1 8.49425
R18396 BIT_SEL[58].n6 BIT_SEL[58] 8.05068
R18397 BIT_SEL[58] BIT_SEL[58].n6 4.57764
R18398 BIT_SEL[58].n6 BIT_SEL[58].t7 117.419
R18399 BIT_SEL[58] BIT_SEL[58].n0 4.57764
R18400 BIT_SEL[58].n0 BIT_SEL[58] 8.05068
R18401 BIT_SEL[58] BIT_SEL[58].n1 4.57764
R18402 BIT_SEL[58].n1 BIT_SEL[58] 8.05068
R18403 BIT_SEL[58] BIT_SEL[58].n2 4.57764
R18404 BIT_SEL[58].n2 BIT_SEL[58] 8.05068
R18405 BIT_SEL[58] BIT_SEL[58].n3 4.57764
R18406 BIT_SEL[58].n3 BIT_SEL[58] 8.05068
R18407 BIT_SEL[58] BIT_SEL[58].n4 4.57764
R18408 BIT_SEL[58].n4 BIT_SEL[58] 8.05068
R18409 BIT_SEL[58] BIT_SEL[58].n5 4.57764
R18410 BIT_SEL[58].n5 BIT_SEL[58] 8.05068
R18411 BIT_SEL[58].t5 BIT_SEL[58] 121.998
R18412 BIT_SEL[58].t4 BIT_SEL[58].n5 117.419
R18413 BIT_SEL[58].t2 BIT_SEL[58].n4 117.419
R18414 BIT_SEL[58].t0 BIT_SEL[58].n3 117.419
R18415 BIT_SEL[58].t6 BIT_SEL[58].n2 117.419
R18416 BIT_SEL[58].t3 BIT_SEL[58].n1 117.419
R18417 BIT_SEL[58].t1 BIT_SEL[58].n0 117.419
R18418 a_20810_38168.t0 a_20810_38168.t1 6.9546
R18419 a_154_24873.t0 a_154_24873.t1 13.9628
R18420 a_110_24961.t0 a_110_24961.t1 19.5535
R18421 a_110_21116.t0 a_110_21116.t1 19.5535
R18422 a_154_21028.t0 a_154_21028.t1 13.9628
R18423 BIT_SEL[7].t0 BIT_SEL[7] 120.195
R18424 BIT_SEL[7] BIT_SEL[7].n0 9.23514
R18425 BIT_SEL[7] BIT_SEL[7].n0 3.39318
R18426 BIT_SEL[7] BIT_SEL[7].n1 9.23514
R18427 BIT_SEL[7].n1 BIT_SEL[7] 3.39318
R18428 BIT_SEL[7] BIT_SEL[7].n2 9.23514
R18429 BIT_SEL[7].n2 BIT_SEL[7] 3.39318
R18430 BIT_SEL[7] BIT_SEL[7].n3 9.23514
R18431 BIT_SEL[7].n3 BIT_SEL[7] 3.39318
R18432 BIT_SEL[7] BIT_SEL[7].n4 9.23514
R18433 BIT_SEL[7].n4 BIT_SEL[7] 3.39318
R18434 BIT_SEL[7] BIT_SEL[7].n5 9.23514
R18435 BIT_SEL[7].n5 BIT_SEL[7] 3.39318
R18436 BIT_SEL[7] BIT_SEL[7].n6 9.23514
R18437 BIT_SEL[7].n6 BIT_SEL[7] 3.39318
R18438 BIT_SEL[7].t1 BIT_SEL[7].n6 116.802
R18439 BIT_SEL[7].t3 BIT_SEL[7].n5 116.802
R18440 BIT_SEL[7].t6 BIT_SEL[7].n4 116.802
R18441 BIT_SEL[7].t5 BIT_SEL[7].n3 116.802
R18442 BIT_SEL[7].t4 BIT_SEL[7].n2 116.802
R18443 BIT_SEL[7].n1 BIT_SEL[7].t2 116.802
R18444 BIT_SEL[7].n0 BIT_SEL[7].t7 116.802
R18445 a_1340_1889.t0 a_1340_1889.t1 5.92075
R18446 BIT_SEL[51].t7 BIT_SEL[51] 117.93
R18447 BIT_SEL[51] BIT_SEL[51].n0 10.6768
R18448 BIT_SEL[51] BIT_SEL[51].n0 1.95157
R18449 BIT_SEL[51] BIT_SEL[51].n1 10.6768
R18450 BIT_SEL[51].n1 BIT_SEL[51] 1.95157
R18451 BIT_SEL[51] BIT_SEL[51].n2 10.6768
R18452 BIT_SEL[51].n2 BIT_SEL[51] 1.95157
R18453 BIT_SEL[51] BIT_SEL[51].n3 10.6768
R18454 BIT_SEL[51].n3 BIT_SEL[51] 1.95157
R18455 BIT_SEL[51] BIT_SEL[51].n4 10.6768
R18456 BIT_SEL[51].n4 BIT_SEL[51] 1.95157
R18457 BIT_SEL[51] BIT_SEL[51].n5 10.6768
R18458 BIT_SEL[51].n5 BIT_SEL[51] 1.95157
R18459 BIT_SEL[51] BIT_SEL[51].n6 10.6768
R18460 BIT_SEL[51].n6 BIT_SEL[51] 1.95157
R18461 BIT_SEL[51].t5 BIT_SEL[51].n6 115.98
R18462 BIT_SEL[51].t4 BIT_SEL[51].n5 115.98
R18463 BIT_SEL[51].t3 BIT_SEL[51].n4 115.98
R18464 BIT_SEL[51].t1 BIT_SEL[51].n3 115.98
R18465 BIT_SEL[51].t0 BIT_SEL[51].n2 115.98
R18466 BIT_SEL[51].n1 BIT_SEL[51].t6 115.98
R18467 BIT_SEL[51].n0 BIT_SEL[51].t2 115.98
R18468 a_20810_26417.t0 a_20810_26417.t1 7.5582
R18469 a_110_2306.t0 a_110_2306.n3 4.44412
R18470 a_110_2306.n3 a_110_2306.n0 0.1805
R18471 a_110_2306.n3 a_110_2306.n2 4.47779
R18472 a_110_2306.n2 a_110_2306.t4 12.3497
R18473 a_110_2306.n2 a_110_2306.t3 17.192
R18474 a_110_2306.n0 a_110_2306.n1 14.1624
R18475 a_110_2306.n1 a_110_2306.t2 12.3497
R18476 a_110_2306.n1 a_110_2306.t5 17.192
R18477 a_110_2306.n0 a_110_2306.t1 8.34715
R18478 OUT[0] OUT[0].n0 9.0005
R18479 OUT[0].n0 OUT[0].t1 8.56064
R18480 OUT[0].n0 OUT[0].t0 4.38216
R18481 a_14320_45309.t0 a_14320_45309.t1 6.38524
R18482 a_1340_42539.t0 a_1340_42539.t1 6.02155
R18483 BIT_SEL[62] BIT_SEL[62].n0 6.01925
R18484 BIT_SEL[62] BIT_SEL[62].n0 6.60907
R18485 BIT_SEL[62] BIT_SEL[62].n1 6.01925
R18486 BIT_SEL[62].n1 BIT_SEL[62] 6.60907
R18487 BIT_SEL[62] BIT_SEL[62].n2 6.01925
R18488 BIT_SEL[62].n2 BIT_SEL[62] 6.60907
R18489 BIT_SEL[62] BIT_SEL[62].n3 6.01925
R18490 BIT_SEL[62].n3 BIT_SEL[62] 6.60907
R18491 BIT_SEL[62] BIT_SEL[62].n4 6.01925
R18492 BIT_SEL[62].n4 BIT_SEL[62] 6.60907
R18493 BIT_SEL[62] BIT_SEL[62].n5 6.01925
R18494 BIT_SEL[62].n5 BIT_SEL[62] 6.60907
R18495 BIT_SEL[62] BIT_SEL[62].n6 6.01925
R18496 BIT_SEL[62].n6 BIT_SEL[62] 6.60907
R18497 BIT_SEL[62].t6 BIT_SEL[62] 124.261
R18498 BIT_SEL[62].t1 BIT_SEL[62].n6 118.243
R18499 BIT_SEL[62].t4 BIT_SEL[62].n5 118.243
R18500 BIT_SEL[62].t2 BIT_SEL[62].n4 118.243
R18501 BIT_SEL[62].t7 BIT_SEL[62].n3 118.243
R18502 BIT_SEL[62].t5 BIT_SEL[62].n2 118.243
R18503 BIT_SEL[62].n1 BIT_SEL[62].t3 118.243
R18504 BIT_SEL[62].n0 BIT_SEL[62].t0 118.243
R18505 a_110_10183.t0 a_110_10183.n3 4.44412
R18506 a_110_10183.n3 a_110_10183.n0 0.1805
R18507 a_110_10183.n3 a_110_10183.n2 4.47779
R18508 a_110_10183.n2 a_110_10183.t5 12.3497
R18509 a_110_10183.n2 a_110_10183.t2 17.192
R18510 a_110_10183.n0 a_110_10183.n1 14.1624
R18511 a_110_10183.n1 a_110_10183.t3 12.3497
R18512 a_110_10183.n1 a_110_10183.t4 17.192
R18513 a_110_10183.n0 a_110_10183.t1 8.34715
R18514 a_110_11079.t0 a_110_11079.n4 4.88081
R18515 a_110_11079.n4 a_110_11079.n5 2.6905
R18516 a_110_11079.n5 a_110_11079.t2 2.06607
R18517 a_110_11079.n5 a_110_11079.t1 2.2382
R18518 a_110_11079.n4 a_110_11079.n0 0.766047
R18519 a_110_11079.n0 a_110_11079.t5 8.68401
R18520 a_110_11079.n2 a_110_11079.n3 5.21793
R18521 a_110_11079.n0 a_110_11079.n2 4.76793
R18522 a_110_11079.n3 a_110_11079.t4 8.51897
R18523 a_110_11079.n3 a_110_11079.t3 4.4523
R18524 a_110_11079.n2 a_110_11079.n1 8.53373
R18525 a_110_11079.n1 a_110_11079.t6 12.3497
R18526 a_110_11079.n1 a_110_11079.t7 17.192
R18527 a_1340_57028.t0 a_1340_57028.t1 5.92117
R18528 a_14320_9398.t0 a_14320_9398.t1 6.39662
R18529 a_154_40627.t0 a_154_40627.t1 13.9628
R18530 a_110_40715.t0 a_110_40715.t1 19.5535
R18531 BIT_SEL[14].n6 BIT_SEL[14] 6.60907
R18532 BIT_SEL[14] BIT_SEL[14].n6 6.01925
R18533 BIT_SEL[14].n6 BIT_SEL[14].t3 118.243
R18534 BIT_SEL[14] BIT_SEL[14].n0 6.01925
R18535 BIT_SEL[14].n0 BIT_SEL[14] 6.60907
R18536 BIT_SEL[14] BIT_SEL[14].n1 6.01925
R18537 BIT_SEL[14].n1 BIT_SEL[14] 6.60907
R18538 BIT_SEL[14] BIT_SEL[14].n2 6.01925
R18539 BIT_SEL[14].n2 BIT_SEL[14] 6.60907
R18540 BIT_SEL[14] BIT_SEL[14].n3 6.01925
R18541 BIT_SEL[14].n3 BIT_SEL[14] 6.60907
R18542 BIT_SEL[14] BIT_SEL[14].n4 6.01925
R18543 BIT_SEL[14].n4 BIT_SEL[14] 6.60907
R18544 BIT_SEL[14] BIT_SEL[14].n5 6.01925
R18545 BIT_SEL[14].n5 BIT_SEL[14] 6.60907
R18546 BIT_SEL[14].t1 BIT_SEL[14] 124.261
R18547 BIT_SEL[14].t4 BIT_SEL[14].n5 118.243
R18548 BIT_SEL[14].t7 BIT_SEL[14].n4 118.243
R18549 BIT_SEL[14].t5 BIT_SEL[14].n3 118.243
R18550 BIT_SEL[14].t2 BIT_SEL[14].n2 118.243
R18551 BIT_SEL[14].t0 BIT_SEL[14].n1 118.243
R18552 BIT_SEL[14].t6 BIT_SEL[14].n0 118.243
R18553 a_1340_23311.t0 a_1340_23311.t1 9.05337
R18554 a_154_5722.t0 a_154_5722.t1 13.9628
R18555 a_110_5810.t0 a_110_5810.t1 19.5535
R18556 a_7830_52657.t0 a_7830_52657.t1 7.18327
R18557 a_638_51026.t0 a_638_51026.n0 7.71211
R18558 a_638_51026.n2 a_638_51026.t59 7.71211
R18559 a_638_51026.n3 a_638_51026.t3 7.71211
R18560 a_638_51026.n4 a_638_51026.t5 7.71211
R18561 a_638_51026.n5 a_638_51026.t58 7.71211
R18562 a_638_51026.n6 a_638_51026.t22 7.71211
R18563 a_638_51026.n7 a_638_51026.t10 7.71211
R18564 a_638_51026.n8 a_638_51026.t20 7.71211
R18565 a_638_51026.n9 a_638_51026.t27 7.71211
R18566 a_638_51026.n10 a_638_51026.t40 7.71211
R18567 a_638_51026.n11 a_638_51026.t55 7.71211
R18568 a_638_51026.n12 a_638_51026.t52 7.71211
R18569 a_638_51026.n13 a_638_51026.t42 7.71211
R18570 a_638_51026.n14 a_638_51026.t6 7.71211
R18571 a_638_51026.n15 a_638_51026.t66 7.71211
R18572 a_638_51026.n16 a_638_51026.t67 7.71211
R18573 a_638_51026.n17 a_638_51026.t32 7.71211
R18574 a_638_51026.n18 a_638_51026.t36 7.71211
R18575 a_638_51026.n19 a_638_51026.t56 7.71211
R18576 a_638_51026.n20 a_638_51026.t2 7.71211
R18577 a_638_51026.n21 a_638_51026.t28 7.71211
R18578 a_638_51026.n22 a_638_51026.t45 7.71211
R18579 a_638_51026.n23 a_638_51026.t65 7.71211
R18580 a_638_51026.n24 a_638_51026.t26 7.71211
R18581 a_638_51026.n25 a_638_51026.t50 7.71211
R18582 a_638_51026.n26 a_638_51026.t54 7.71211
R18583 a_638_51026.n27 a_638_51026.t29 7.71211
R18584 a_638_51026.n28 a_638_51026.t57 7.71211
R18585 a_638_51026.n29 a_638_51026.t46 7.71211
R18586 a_638_51026.n30 a_638_51026.t41 7.71211
R18587 a_638_51026.n31 a_638_51026.t39 7.71211
R18588 a_638_51026.n32 a_638_51026.t64 7.71211
R18589 a_638_51026.n3 a_638_51026.n2 0.427167
R18590 a_638_51026.n4 a_638_51026.n3 0.427167
R18591 a_638_51026.n5 a_638_51026.n4 0.427167
R18592 a_638_51026.n6 a_638_51026.n5 0.427167
R18593 a_638_51026.n7 a_638_51026.n6 0.427167
R18594 a_638_51026.n8 a_638_51026.n7 0.427167
R18595 a_638_51026.n9 a_638_51026.n8 0.427167
R18596 a_638_51026.n10 a_638_51026.n9 0.619389
R18597 a_638_51026.n11 a_638_51026.n10 0.427167
R18598 a_638_51026.n12 a_638_51026.n11 0.427167
R18599 a_638_51026.n13 a_638_51026.n12 0.427167
R18600 a_638_51026.n14 a_638_51026.n13 0.427167
R18601 a_638_51026.n15 a_638_51026.n14 0.427167
R18602 a_638_51026.n16 a_638_51026.n15 0.427167
R18603 a_638_51026.n17 a_638_51026.n16 0.427167
R18604 a_638_51026.n18 a_638_51026.n17 0.619389
R18605 a_638_51026.n0 a_638_51026.n18 0.427167
R18606 a_638_51026.n0 a_638_51026.n19 0.427167
R18607 a_638_51026.n19 a_638_51026.n20 0.427167
R18608 a_638_51026.n20 a_638_51026.n21 0.427167
R18609 a_638_51026.n21 a_638_51026.n22 0.427167
R18610 a_638_51026.n22 a_638_51026.n23 0.427167
R18611 a_638_51026.n23 a_638_51026.n24 0.427167
R18612 a_638_51026.n24 a_638_51026.n25 0.619389
R18613 a_638_51026.n25 a_638_51026.n26 0.427167
R18614 a_638_51026.n26 a_638_51026.n27 0.427167
R18615 a_638_51026.n27 a_638_51026.n28 0.427167
R18616 a_638_51026.n28 a_638_51026.n29 0.427167
R18617 a_638_51026.n29 a_638_51026.n30 0.427167
R18618 a_638_51026.n30 a_638_51026.n31 0.427167
R18619 a_638_51026.n31 a_638_51026.n32 0.427167
R18620 a_638_51026.n32 a_638_51026.n1 0.334944
R18621 a_638_51026.n1 a_638_51026.n33 0.227167
R18622 a_638_51026.n34 a_638_51026.n35 0.466493
R18623 a_638_51026.n2 a_638_51026.n34 0.69448
R18624 a_638_51026.n35 a_638_51026.t43 7.71211
R18625 a_638_51026.n36 a_638_51026.t1 7.71211
R18626 a_638_51026.n37 a_638_51026.t44 7.71211
R18627 a_638_51026.n38 a_638_51026.t34 7.71211
R18628 a_638_51026.n39 a_638_51026.t9 7.71211
R18629 a_638_51026.n40 a_638_51026.t68 7.71211
R18630 a_638_51026.n41 a_638_51026.t12 7.71211
R18631 a_638_51026.n42 a_638_51026.t53 7.71211
R18632 a_638_51026.n43 a_638_51026.t21 7.71211
R18633 a_638_51026.n44 a_638_51026.t18 7.71211
R18634 a_638_51026.n45 a_638_51026.t15 7.71211
R18635 a_638_51026.n46 a_638_51026.t30 7.71211
R18636 a_638_51026.n47 a_638_51026.t48 7.71211
R18637 a_638_51026.n48 a_638_51026.t49 7.71211
R18638 a_638_51026.n49 a_638_51026.t7 7.71211
R18639 a_638_51026.n50 a_638_51026.t25 7.71211
R18640 a_638_51026.n51 a_638_51026.t33 7.71211
R18641 a_638_51026.n52 a_638_51026.t17 7.71211
R18642 a_638_51026.n53 a_638_51026.t47 7.71211
R18643 a_638_51026.n54 a_638_51026.t14 7.71211
R18644 a_638_51026.n55 a_638_51026.t16 7.71211
R18645 a_638_51026.n56 a_638_51026.t4 7.71211
R18646 a_638_51026.n57 a_638_51026.t51 7.71211
R18647 a_638_51026.n58 a_638_51026.t24 7.71211
R18648 a_638_51026.n59 a_638_51026.t23 7.71211
R18649 a_638_51026.n60 a_638_51026.t8 7.71211
R18650 a_638_51026.n61 a_638_51026.t37 7.71211
R18651 a_638_51026.n62 a_638_51026.t19 7.71211
R18652 a_638_51026.n63 a_638_51026.t38 7.71211
R18653 a_638_51026.n64 a_638_51026.t13 7.71211
R18654 a_638_51026.n65 a_638_51026.t35 7.71211
R18655 a_638_51026.n66 a_638_51026.t11 7.71211
R18656 a_638_51026.n35 a_638_51026.n36 0.427167
R18657 a_638_51026.n36 a_638_51026.n37 0.427167
R18658 a_638_51026.n37 a_638_51026.n38 0.427167
R18659 a_638_51026.n38 a_638_51026.n39 0.427167
R18660 a_638_51026.n39 a_638_51026.n40 0.427167
R18661 a_638_51026.n40 a_638_51026.n41 0.427167
R18662 a_638_51026.n41 a_638_51026.n42 0.427167
R18663 a_638_51026.n42 a_638_51026.n43 0.619389
R18664 a_638_51026.n43 a_638_51026.n44 0.427167
R18665 a_638_51026.n44 a_638_51026.n45 0.427167
R18666 a_638_51026.n45 a_638_51026.n46 0.427167
R18667 a_638_51026.n46 a_638_51026.n47 0.427167
R18668 a_638_51026.n47 a_638_51026.n48 0.427167
R18669 a_638_51026.n48 a_638_51026.n49 0.427167
R18670 a_638_51026.n49 a_638_51026.n50 0.427167
R18671 a_638_51026.n50 a_638_51026.n51 0.619389
R18672 a_638_51026.n51 a_638_51026.n52 0.427167
R18673 a_638_51026.n52 a_638_51026.n53 0.427167
R18674 a_638_51026.n53 a_638_51026.n54 0.427167
R18675 a_638_51026.n54 a_638_51026.n55 0.427167
R18676 a_638_51026.n55 a_638_51026.n56 0.427167
R18677 a_638_51026.n56 a_638_51026.n57 0.427167
R18678 a_638_51026.n57 a_638_51026.n58 0.427167
R18679 a_638_51026.n58 a_638_51026.n59 0.619389
R18680 a_638_51026.n60 a_638_51026.n59 0.427167
R18681 a_638_51026.n61 a_638_51026.n60 0.427167
R18682 a_638_51026.n62 a_638_51026.n61 0.427167
R18683 a_638_51026.n63 a_638_51026.n62 0.427167
R18684 a_638_51026.n64 a_638_51026.n63 0.427167
R18685 a_638_51026.n65 a_638_51026.n64 0.427167
R18686 a_638_51026.n66 a_638_51026.n65 0.427167
R18687 a_638_51026.n71 a_638_51026.n66 0.548278
R18688 a_638_51026.n71 a_638_51026.n68 0.227167
R18689 a_638_51026.n72 a_638_51026.n71 4.74618
R18690 a_638_51026.n1 a_638_51026.n72 4.60509
R18691 a_638_51026.n72 a_638_51026.t60 0.113082
R18692 a_638_51026.n70 a_638_51026.n69 0.0655
R18693 a_638_51026.n70 a_638_51026.n68 4.74618
R18694 a_638_51026.n33 a_638_51026.n70 4.60509
R18695 a_638_51026.n69 a_638_51026.t62 0.0480817
R18696 a_638_51026.n69 a_638_51026.t63 0.0480817
R18697 a_638_51026.n68 a_638_51026.n67 4.96756
R18698 a_638_51026.n33 a_638_51026.n67 4.83019
R18699 a_638_51026.n67 a_638_51026.t61 0.113082
R18700 a_638_51026.n34 a_638_51026.t31 9.85476
R18701 a_20810_26785.t0 a_20810_26785.t1 6.02155
R18702 a_14320_1521.t0 a_14320_1521.t1 6.39548
R18703 a_1340_55395.t0 a_1340_55395.t1 9.52407
R18704 BIT_SEL[40] BIT_SEL[40].n0 3.98621
R18705 BIT_SEL[40] BIT_SEL[40].n0 8.64211
R18706 BIT_SEL[40] BIT_SEL[40].n1 3.98621
R18707 BIT_SEL[40].n1 BIT_SEL[40] 8.64211
R18708 BIT_SEL[40] BIT_SEL[40].n2 3.98621
R18709 BIT_SEL[40].n2 BIT_SEL[40] 8.64211
R18710 BIT_SEL[40] BIT_SEL[40].n3 3.98621
R18711 BIT_SEL[40].n3 BIT_SEL[40] 8.64211
R18712 BIT_SEL[40] BIT_SEL[40].n4 3.98621
R18713 BIT_SEL[40].n4 BIT_SEL[40] 8.64211
R18714 BIT_SEL[40] BIT_SEL[40].n5 3.98621
R18715 BIT_SEL[40].n5 BIT_SEL[40] 8.64211
R18716 BIT_SEL[40] BIT_SEL[40].n6 3.98621
R18717 BIT_SEL[40].n6 BIT_SEL[40] 8.64211
R18718 BIT_SEL[40].t1 BIT_SEL[40] 120.995
R18719 BIT_SEL[40].t3 BIT_SEL[40].n6 117.008
R18720 BIT_SEL[40].t0 BIT_SEL[40].n5 117.008
R18721 BIT_SEL[40].t7 BIT_SEL[40].n4 117.008
R18722 BIT_SEL[40].t5 BIT_SEL[40].n3 117.008
R18723 BIT_SEL[40].t4 BIT_SEL[40].n2 117.008
R18724 BIT_SEL[40].n1 BIT_SEL[40].t2 117.008
R18725 BIT_SEL[40].n0 BIT_SEL[40].t6 117.008
R18726 a_14320_45677.t0 a_14320_45677.t1 5.92611
R18727 BIT_SEL[48] BIT_SEL[48].n0 1.36175
R18728 BIT_SEL[48] BIT_SEL[48].n0 11.2666
R18729 BIT_SEL[48] BIT_SEL[48].n1 1.36175
R18730 BIT_SEL[48].n1 BIT_SEL[48] 11.2666
R18731 BIT_SEL[48] BIT_SEL[48].n2 1.36175
R18732 BIT_SEL[48].n2 BIT_SEL[48] 11.2666
R18733 BIT_SEL[48] BIT_SEL[48].n3 1.36175
R18734 BIT_SEL[48].n3 BIT_SEL[48] 11.2666
R18735 BIT_SEL[48] BIT_SEL[48].n4 1.36175
R18736 BIT_SEL[48].n4 BIT_SEL[48] 11.2666
R18737 BIT_SEL[48] BIT_SEL[48].n5 1.36175
R18738 BIT_SEL[48].n5 BIT_SEL[48] 11.2666
R18739 BIT_SEL[48] BIT_SEL[48].n6 1.36175
R18740 BIT_SEL[48].n6 BIT_SEL[48] 11.2666
R18741 BIT_SEL[48].t2 BIT_SEL[48] 116.835
R18742 BIT_SEL[48].t5 BIT_SEL[48].n6 115.474
R18743 BIT_SEL[48].t7 BIT_SEL[48].n5 115.474
R18744 BIT_SEL[48].t4 BIT_SEL[48].n4 115.474
R18745 BIT_SEL[48].t3 BIT_SEL[48].n3 115.474
R18746 BIT_SEL[48].t0 BIT_SEL[48].n2 115.474
R18747 BIT_SEL[48].n1 BIT_SEL[48].t6 115.474
R18748 BIT_SEL[48].n0 BIT_SEL[48].t1 115.474
R18749 a_20718_19835.t0 a_20718_19835.t1 6.66648
R18750 COL_PROG_N[0] COL_PROG_N[0].n0 0.0965
R18751 COL_PROG_N[0].n0 COL_PROG_N[0].n1 0.3065
R18752 COL_PROG_N[0].n1 COL_PROG_N[0].n2 0.3065
R18753 COL_PROG_N[0].n2 COL_PROG_N[0].t2 292.788
R18754 COL_PROG_N[0].n2 COL_PROG_N[0].t1 292.481
R18755 COL_PROG_N[0].n1 COL_PROG_N[0].t0 292.481
R18756 COL_PROG_N[0].n0 COL_PROG_N[0].t3 292.481
R18757 a_154_62653.t0 a_154_62653.t1 13.9628
R18758 a_110_62741.t0 a_110_62741.t1 19.5535
R18759 BIT_SEL[15].n6 BIT_SEL[15] 6.01764
R18760 BIT_SEL[15] BIT_SEL[15].n6 6.61068
R18761 BIT_SEL[15] BIT_SEL[15].t5 124.466
R18762 BIT_SEL[15].n6 BIT_SEL[15].t4 118.448
R18763 BIT_SEL[15] BIT_SEL[15].n0 6.61068
R18764 BIT_SEL[15].n0 BIT_SEL[15] 6.01764
R18765 BIT_SEL[15] BIT_SEL[15].n1 6.61068
R18766 BIT_SEL[15].n1 BIT_SEL[15] 6.01764
R18767 BIT_SEL[15] BIT_SEL[15].n2 6.61068
R18768 BIT_SEL[15].n2 BIT_SEL[15] 6.01764
R18769 BIT_SEL[15] BIT_SEL[15].n3 6.61068
R18770 BIT_SEL[15].n3 BIT_SEL[15] 6.01764
R18771 BIT_SEL[15] BIT_SEL[15].n4 6.61068
R18772 BIT_SEL[15].n4 BIT_SEL[15] 6.01764
R18773 BIT_SEL[15] BIT_SEL[15].n5 6.61068
R18774 BIT_SEL[15].n5 BIT_SEL[15] 6.01764
R18775 BIT_SEL[15].t1 BIT_SEL[15].n5 118.448
R18776 BIT_SEL[15].t7 BIT_SEL[15].n4 118.448
R18777 BIT_SEL[15].t6 BIT_SEL[15].n3 118.448
R18778 BIT_SEL[15].t3 BIT_SEL[15].n2 118.448
R18779 BIT_SEL[15].t0 BIT_SEL[15].n1 118.448
R18780 BIT_SEL[15].t2 BIT_SEL[15].n0 118.448
R18781 a_1340_23887.t0 a_1340_23887.t1 9.52293
R18782 a_20810_42539.t0 a_20810_42539.t1 6.02155
R18783 a_14320_25152.t0 a_14320_25152.t1 6.39548
R18784 a_7830_14169.t0 a_7830_14169.t1 5.92569
R18785 a_14320_61431.t0 a_14320_61431.t1 5.92569
R18786 BIT_SEL[22] BIT_SEL[22].n0 3.39479
R18787 BIT_SEL[22] BIT_SEL[22].n0 9.23354
R18788 BIT_SEL[22] BIT_SEL[22].n1 3.39479
R18789 BIT_SEL[22].n1 BIT_SEL[22] 9.23354
R18790 BIT_SEL[22] BIT_SEL[22].n2 3.39479
R18791 BIT_SEL[22].n2 BIT_SEL[22] 9.23354
R18792 BIT_SEL[22] BIT_SEL[22].n3 3.39479
R18793 BIT_SEL[22].n3 BIT_SEL[22] 9.23354
R18794 BIT_SEL[22] BIT_SEL[22].n4 3.39479
R18795 BIT_SEL[22].n4 BIT_SEL[22] 9.23354
R18796 BIT_SEL[22] BIT_SEL[22].n5 3.39479
R18797 BIT_SEL[22].n5 BIT_SEL[22] 9.23354
R18798 BIT_SEL[22] BIT_SEL[22].n6 3.39479
R18799 BIT_SEL[22].n6 BIT_SEL[22] 9.23354
R18800 BIT_SEL[22].t6 BIT_SEL[22] 119.992
R18801 BIT_SEL[22].t5 BIT_SEL[22].n6 116.597
R18802 BIT_SEL[22].t3 BIT_SEL[22].n5 116.597
R18803 BIT_SEL[22].t1 BIT_SEL[22].n4 116.597
R18804 BIT_SEL[22].t0 BIT_SEL[22].n3 116.597
R18805 BIT_SEL[22].t4 BIT_SEL[22].n2 116.597
R18806 BIT_SEL[22].n1 BIT_SEL[22].t2 116.597
R18807 BIT_SEL[22].n0 BIT_SEL[22].t7 116.597
R18808 a_7830_29555.t0 a_7830_29555.t1 6.38411
R18809 BIT_SEL[20] BIT_SEL[20].n0 2.54461
R18810 BIT_SEL[20] BIT_SEL[20].n0 10.0837
R18811 BIT_SEL[20] BIT_SEL[20].n1 2.54461
R18812 BIT_SEL[20].n1 BIT_SEL[20] 10.0837
R18813 BIT_SEL[20] BIT_SEL[20].n2 2.54461
R18814 BIT_SEL[20].n2 BIT_SEL[20] 10.0837
R18815 BIT_SEL[20] BIT_SEL[20].n3 2.54461
R18816 BIT_SEL[20].n3 BIT_SEL[20] 10.0837
R18817 BIT_SEL[20] BIT_SEL[20].n4 2.54461
R18818 BIT_SEL[20].n4 BIT_SEL[20] 10.0837
R18819 BIT_SEL[20] BIT_SEL[20].n5 2.54461
R18820 BIT_SEL[20].n5 BIT_SEL[20] 10.0837
R18821 BIT_SEL[20] BIT_SEL[20].n6 2.54461
R18822 BIT_SEL[20].n6 BIT_SEL[20] 10.0837
R18823 BIT_SEL[20].t4 BIT_SEL[20] 118.73
R18824 BIT_SEL[20].t2 BIT_SEL[20].n6 116.186
R18825 BIT_SEL[20].t0 BIT_SEL[20].n5 116.186
R18826 BIT_SEL[20].t1 BIT_SEL[20].n4 116.186
R18827 BIT_SEL[20].t7 BIT_SEL[20].n3 116.186
R18828 BIT_SEL[20].t3 BIT_SEL[20].n2 116.186
R18829 BIT_SEL[20].n1 BIT_SEL[20].t5 116.186
R18830 BIT_SEL[20].n0 BIT_SEL[20].t6 116.186
R18831 a_7830_44780.t0 a_7830_44780.t1 7.18327
R18832 a_20810_21149.t0 a_20810_21149.t1 7.18327
R18833 a_20810_57556.t0 a_20810_57556.t1 6.71945
R18834 a_14228_4081.t0 a_14228_4081.t1 6.66648
R18835 a_20810_58293.t0 a_20810_58293.t1 6.02155
R18836 a_14320_40906.t0 a_14320_40906.t1 6.39548
R18837 a_110_37318.t0 a_110_37318.t1 19.5535
R18838 a_154_37230.t0 a_154_37230.t1 13.9628
R18839 BIT_SEL[34] BIT_SEL[34].n0 1.95318
R18840 BIT_SEL[34] BIT_SEL[34].n0 10.6751
R18841 BIT_SEL[34] BIT_SEL[34].n1 1.95318
R18842 BIT_SEL[34].n1 BIT_SEL[34] 10.6751
R18843 BIT_SEL[34] BIT_SEL[34].n2 1.95318
R18844 BIT_SEL[34].n2 BIT_SEL[34] 10.6751
R18845 BIT_SEL[34] BIT_SEL[34].n3 1.95318
R18846 BIT_SEL[34].n3 BIT_SEL[34] 10.6751
R18847 BIT_SEL[34] BIT_SEL[34].n4 1.95318
R18848 BIT_SEL[34].n4 BIT_SEL[34] 10.6751
R18849 BIT_SEL[34] BIT_SEL[34].n5 1.95318
R18850 BIT_SEL[34].n5 BIT_SEL[34] 10.6751
R18851 BIT_SEL[34] BIT_SEL[34].n6 1.95318
R18852 BIT_SEL[34].n6 BIT_SEL[34] 10.6751
R18853 BIT_SEL[34].t1 BIT_SEL[34] 117.727
R18854 BIT_SEL[34].t7 BIT_SEL[34].n6 115.775
R18855 BIT_SEL[34].t5 BIT_SEL[34].n5 115.775
R18856 BIT_SEL[34].t4 BIT_SEL[34].n4 115.775
R18857 BIT_SEL[34].t3 BIT_SEL[34].n3 115.775
R18858 BIT_SEL[34].t6 BIT_SEL[34].n2 115.775
R18859 BIT_SEL[34].n1 BIT_SEL[34].t0 115.775
R18860 BIT_SEL[34].n0 BIT_SEL[34].t2 115.775
R18861 a_14320_12904.t0 a_14320_12904.t1 8.02156
R18862 a_7830_29923.t0 a_7830_29923.t1 5.92569
R18863 a_154_36110.t0 a_154_36110.t1 13.9628
R18864 a_110_36198.t0 a_110_36198.t1 19.5535
R18865 a_110_26833.t0 a_110_26833.n4 4.88081
R18866 a_110_26833.n4 a_110_26833.n5 2.6905
R18867 a_110_26833.n5 a_110_26833.t1 2.06607
R18868 a_110_26833.n5 a_110_26833.t2 2.2382
R18869 a_110_26833.n4 a_110_26833.n0 0.766047
R18870 a_110_26833.n0 a_110_26833.t4 8.68401
R18871 a_110_26833.n2 a_110_26833.n3 5.21793
R18872 a_110_26833.n0 a_110_26833.n2 4.76793
R18873 a_110_26833.n3 a_110_26833.t3 8.51897
R18874 a_110_26833.n3 a_110_26833.t5 4.4523
R18875 a_110_26833.n2 a_110_26833.n1 8.53373
R18876 a_110_26833.n1 a_110_26833.t7 12.3497
R18877 a_110_26833.n1 a_110_26833.t6 17.192
R18878 a_110_25937.t0 a_110_25937.n3 4.44412
R18879 a_110_25937.n3 a_110_25937.n0 0.1805
R18880 a_110_25937.n3 a_110_25937.n2 4.47779
R18881 a_110_25937.n2 a_110_25937.t3 12.3497
R18882 a_110_25937.n2 a_110_25937.t4 17.192
R18883 a_110_25937.n0 a_110_25937.n1 14.1624
R18884 a_110_25937.n1 a_110_25937.t5 12.3497
R18885 a_110_25937.n1 a_110_25937.t2 17.192
R18886 a_110_25937.n0 a_110_25937.t1 8.34715
R18887 a_110_32390.t0 a_110_32390.t1 19.5535
R18888 a_154_32302.t0 a_154_32302.t1 13.9628
R18889 a_638_19518.t0 a_638_19518.n0 7.71211
R18890 a_638_19518.n1 a_638_19518.t66 7.71211
R18891 a_638_19518.n2 a_638_19518.t34 7.71211
R18892 a_638_19518.n3 a_638_19518.t47 7.71211
R18893 a_638_19518.n4 a_638_19518.t60 7.71211
R18894 a_638_19518.n5 a_638_19518.t15 7.71211
R18895 a_638_19518.n6 a_638_19518.t61 7.71211
R18896 a_638_19518.n7 a_638_19518.t40 7.71211
R18897 a_638_19518.n8 a_638_19518.t51 7.71211
R18898 a_638_19518.n9 a_638_19518.t26 7.71211
R18899 a_638_19518.n10 a_638_19518.t6 7.71211
R18900 a_638_19518.n11 a_638_19518.t29 7.71211
R18901 a_638_19518.n12 a_638_19518.t1 7.71211
R18902 a_638_19518.n13 a_638_19518.t45 7.71211
R18903 a_638_19518.n14 a_638_19518.t16 7.71211
R18904 a_638_19518.n15 a_638_19518.t17 7.71211
R18905 a_638_19518.n16 a_638_19518.t35 7.71211
R18906 a_638_19518.n17 a_638_19518.t21 7.71211
R18907 a_638_19518.n18 a_638_19518.t63 7.71211
R18908 a_638_19518.n19 a_638_19518.t39 7.71211
R18909 a_638_19518.n20 a_638_19518.t54 7.71211
R18910 a_638_19518.n21 a_638_19518.t56 7.71211
R18911 a_638_19518.n22 a_638_19518.t68 7.71211
R18912 a_638_19518.n23 a_638_19518.t9 7.71211
R18913 a_638_19518.n24 a_638_19518.t41 7.71211
R18914 a_638_19518.n25 a_638_19518.t19 7.71211
R18915 a_638_19518.n26 a_638_19518.t65 7.71211
R18916 a_638_19518.n27 a_638_19518.t25 7.71211
R18917 a_638_19518.n28 a_638_19518.t38 7.71211
R18918 a_638_19518.n29 a_638_19518.t36 7.71211
R18919 a_638_19518.n30 a_638_19518.t12 7.71211
R18920 a_638_19518.n31 a_638_19518.t43 7.71211
R18921 a_638_19518.n2 a_638_19518.n1 0.427167
R18922 a_638_19518.n3 a_638_19518.n2 0.427167
R18923 a_638_19518.n4 a_638_19518.n3 0.427167
R18924 a_638_19518.n5 a_638_19518.n4 0.427167
R18925 a_638_19518.n6 a_638_19518.n5 0.427167
R18926 a_638_19518.n7 a_638_19518.n6 0.427167
R18927 a_638_19518.n8 a_638_19518.n7 0.427167
R18928 a_638_19518.n9 a_638_19518.n8 0.619389
R18929 a_638_19518.n10 a_638_19518.n9 0.427167
R18930 a_638_19518.n11 a_638_19518.n10 0.427167
R18931 a_638_19518.n12 a_638_19518.n11 0.427167
R18932 a_638_19518.n13 a_638_19518.n12 0.427167
R18933 a_638_19518.n0 a_638_19518.n13 0.427167
R18934 a_638_19518.n0 a_638_19518.n14 0.427167
R18935 a_638_19518.n14 a_638_19518.n15 0.427167
R18936 a_638_19518.n15 a_638_19518.n16 0.619389
R18937 a_638_19518.n16 a_638_19518.n17 0.427167
R18938 a_638_19518.n17 a_638_19518.n18 0.427167
R18939 a_638_19518.n18 a_638_19518.n19 0.427167
R18940 a_638_19518.n19 a_638_19518.n20 0.427167
R18941 a_638_19518.n20 a_638_19518.n21 0.427167
R18942 a_638_19518.n21 a_638_19518.n22 0.427167
R18943 a_638_19518.n22 a_638_19518.n23 0.427167
R18944 a_638_19518.n23 a_638_19518.n24 0.619389
R18945 a_638_19518.n24 a_638_19518.n25 0.427167
R18946 a_638_19518.n25 a_638_19518.n26 0.427167
R18947 a_638_19518.n26 a_638_19518.n27 0.427167
R18948 a_638_19518.n27 a_638_19518.n28 0.427167
R18949 a_638_19518.n28 a_638_19518.n29 0.427167
R18950 a_638_19518.n29 a_638_19518.n30 0.427167
R18951 a_638_19518.n30 a_638_19518.n31 0.427167
R18952 a_638_19518.n31 a_638_19518.n34 0.548278
R18953 a_638_19518.n34 a_638_19518.n70 0.227167
R18954 a_638_19518.n1 a_638_19518.n32 0.466493
R18955 a_638_19518.n36 a_638_19518.t23 7.71211
R18956 a_638_19518.n37 a_638_19518.t44 7.71211
R18957 a_638_19518.n38 a_638_19518.t18 7.71211
R18958 a_638_19518.n39 a_638_19518.t8 7.71211
R18959 a_638_19518.n40 a_638_19518.t33 7.71211
R18960 a_638_19518.n41 a_638_19518.t64 7.71211
R18961 a_638_19518.n42 a_638_19518.t37 7.71211
R18962 a_638_19518.n43 a_638_19518.t48 7.71211
R18963 a_638_19518.n44 a_638_19518.t50 7.71211
R18964 a_638_19518.n45 a_638_19518.t55 7.71211
R18965 a_638_19518.n46 a_638_19518.t28 7.71211
R18966 a_638_19518.n47 a_638_19518.t5 7.71211
R18967 a_638_19518.n48 a_638_19518.t13 7.71211
R18968 a_638_19518.n49 a_638_19518.t20 7.71211
R18969 a_638_19518.n50 a_638_19518.t42 7.71211
R18970 a_638_19518.n51 a_638_19518.t10 7.71211
R18971 a_638_19518.n52 a_638_19518.t67 7.71211
R18972 a_638_19518.n53 a_638_19518.t31 7.71211
R18973 a_638_19518.n54 a_638_19518.t4 7.71211
R18974 a_638_19518.n55 a_638_19518.t22 7.71211
R18975 a_638_19518.n56 a_638_19518.t32 7.71211
R18976 a_638_19518.n57 a_638_19518.t46 7.71211
R18977 a_638_19518.n58 a_638_19518.t7 7.71211
R18978 a_638_19518.n59 a_638_19518.t30 7.71211
R18979 a_638_19518.n60 a_638_19518.t3 7.71211
R18980 a_638_19518.n61 a_638_19518.t27 7.71211
R18981 a_638_19518.n62 a_638_19518.t2 7.71211
R18982 a_638_19518.n63 a_638_19518.t53 7.71211
R18983 a_638_19518.n64 a_638_19518.t62 7.71211
R18984 a_638_19518.n65 a_638_19518.t14 7.71211
R18985 a_638_19518.n66 a_638_19518.t49 7.71211
R18986 a_638_19518.n67 a_638_19518.t11 7.71211
R18987 a_638_19518.n32 a_638_19518.n36 0.69448
R18988 a_638_19518.n36 a_638_19518.n37 0.427167
R18989 a_638_19518.n37 a_638_19518.n38 0.427167
R18990 a_638_19518.n38 a_638_19518.n39 0.427167
R18991 a_638_19518.n39 a_638_19518.n40 0.427167
R18992 a_638_19518.n40 a_638_19518.n41 0.427167
R18993 a_638_19518.n41 a_638_19518.n42 0.427167
R18994 a_638_19518.n42 a_638_19518.n43 0.427167
R18995 a_638_19518.n43 a_638_19518.n44 0.619389
R18996 a_638_19518.n44 a_638_19518.n45 0.427167
R18997 a_638_19518.n45 a_638_19518.n46 0.427167
R18998 a_638_19518.n46 a_638_19518.n47 0.427167
R18999 a_638_19518.n47 a_638_19518.n48 0.427167
R19000 a_638_19518.n48 a_638_19518.n49 0.427167
R19001 a_638_19518.n49 a_638_19518.n50 0.427167
R19002 a_638_19518.n50 a_638_19518.n51 0.427167
R19003 a_638_19518.n51 a_638_19518.n52 0.619389
R19004 a_638_19518.n52 a_638_19518.n53 0.427167
R19005 a_638_19518.n53 a_638_19518.n54 0.427167
R19006 a_638_19518.n54 a_638_19518.n55 0.427167
R19007 a_638_19518.n55 a_638_19518.n56 0.427167
R19008 a_638_19518.n56 a_638_19518.n57 0.427167
R19009 a_638_19518.n57 a_638_19518.n58 0.427167
R19010 a_638_19518.n58 a_638_19518.n59 0.427167
R19011 a_638_19518.n59 a_638_19518.n60 0.619389
R19012 a_638_19518.n60 a_638_19518.n61 0.427167
R19013 a_638_19518.n61 a_638_19518.n62 0.427167
R19014 a_638_19518.n62 a_638_19518.n63 0.427167
R19015 a_638_19518.n63 a_638_19518.n64 0.427167
R19016 a_638_19518.n64 a_638_19518.n65 0.427167
R19017 a_638_19518.n66 a_638_19518.n65 0.427167
R19018 a_638_19518.n67 a_638_19518.n66 0.427167
R19019 a_638_19518.n35 a_638_19518.n67 0.334944
R19020 a_638_19518.n35 a_638_19518.n71 0.227167
R19021 a_638_19518.n70 a_638_19518.n72 4.96756
R19022 a_638_19518.n72 a_638_19518.n71 4.83019
R19023 a_638_19518.n72 a_638_19518.t58 0.113082
R19024 a_638_19518.n69 a_638_19518.n68 0.0655
R19025 a_638_19518.n69 a_638_19518.n71 4.60509
R19026 a_638_19518.n70 a_638_19518.n69 4.74618
R19027 a_638_19518.n68 a_638_19518.t59 0.0480817
R19028 a_638_19518.n68 a_638_19518.t57 0.0480817
R19029 a_638_19518.n33 a_638_19518.n35 4.60509
R19030 a_638_19518.n34 a_638_19518.n33 4.74618
R19031 a_638_19518.n33 a_638_19518.t52 0.113082
R19032 a_638_19518.n32 a_638_19518.t24 9.85476
R19033 a_7830_16010.t0 a_7830_16010.t1 9.52407
R19034 a_7830_45677.t0 a_7830_45677.t1 5.92569
R19035 BIT_SEL[17].t7 BIT_SEL[17] 116.918
R19036 BIT_SEL[17] BIT_SEL[17].n0 11.2682
R19037 BIT_SEL[17] BIT_SEL[17].n0 1.36014
R19038 BIT_SEL[17] BIT_SEL[17].n1 11.2682
R19039 BIT_SEL[17].n1 BIT_SEL[17] 1.36014
R19040 BIT_SEL[17] BIT_SEL[17].n2 11.2682
R19041 BIT_SEL[17].n2 BIT_SEL[17] 1.36014
R19042 BIT_SEL[17] BIT_SEL[17].n3 11.2682
R19043 BIT_SEL[17].n3 BIT_SEL[17] 1.36014
R19044 BIT_SEL[17] BIT_SEL[17].n4 11.2682
R19045 BIT_SEL[17].n4 BIT_SEL[17] 1.36014
R19046 BIT_SEL[17] BIT_SEL[17].n5 11.2682
R19047 BIT_SEL[17].n5 BIT_SEL[17] 1.36014
R19048 BIT_SEL[17] BIT_SEL[17].n6 11.2682
R19049 BIT_SEL[17].n6 BIT_SEL[17] 1.36014
R19050 BIT_SEL[17].t3 BIT_SEL[17].n6 115.558
R19051 BIT_SEL[17].t6 BIT_SEL[17].n5 115.558
R19052 BIT_SEL[17].t2 BIT_SEL[17].n4 115.558
R19053 BIT_SEL[17].t4 BIT_SEL[17].n3 115.558
R19054 BIT_SEL[17].t1 BIT_SEL[17].n2 115.558
R19055 BIT_SEL[17].n1 BIT_SEL[17].t0 115.558
R19056 BIT_SEL[17].n0 BIT_SEL[17].t5 115.558
R19057 a_7830_18908.t0 a_7830_18908.t1 6.02155
R19058 BIT_SEL[56].n6 BIT_SEL[56] 8.64211
R19059 BIT_SEL[56] BIT_SEL[56].n6 3.98621
R19060 BIT_SEL[56].n6 BIT_SEL[56].t0 117.008
R19061 BIT_SEL[56] BIT_SEL[56].n0 3.98621
R19062 BIT_SEL[56].n0 BIT_SEL[56] 8.64211
R19063 BIT_SEL[56] BIT_SEL[56].n1 3.98621
R19064 BIT_SEL[56].n1 BIT_SEL[56] 8.64211
R19065 BIT_SEL[56] BIT_SEL[56].n2 3.98621
R19066 BIT_SEL[56].n2 BIT_SEL[56] 8.64211
R19067 BIT_SEL[56] BIT_SEL[56].n3 3.98621
R19068 BIT_SEL[56].n3 BIT_SEL[56] 8.64211
R19069 BIT_SEL[56] BIT_SEL[56].n4 3.98621
R19070 BIT_SEL[56].n4 BIT_SEL[56] 8.64211
R19071 BIT_SEL[56] BIT_SEL[56].n5 3.98621
R19072 BIT_SEL[56].n5 BIT_SEL[56] 8.64211
R19073 BIT_SEL[56].t2 BIT_SEL[56] 120.995
R19074 BIT_SEL[56].t4 BIT_SEL[56].n5 117.008
R19075 BIT_SEL[56].t1 BIT_SEL[56].n4 117.008
R19076 BIT_SEL[56].t7 BIT_SEL[56].n3 117.008
R19077 BIT_SEL[56].t6 BIT_SEL[56].n2 117.008
R19078 BIT_SEL[56].t5 BIT_SEL[56].n1 117.008
R19079 BIT_SEL[56].t3 BIT_SEL[56].n0 117.008
R19080 a_20810_6292.t0 a_20810_6292.t1 5.92569
R19081 a_154_8671.t0 a_154_8671.t1 13.9628
R19082 a_110_8759.t0 a_110_8759.t1 19.5535
R19083 a_14320_14169.t0 a_14320_14169.t1 5.92611
R19084 BIT_SEL[13].n6 BIT_SEL[13] 5.42621
R19085 BIT_SEL[13] BIT_SEL[13].n6 7.20211
R19086 BIT_SEL[13] BIT_SEL[13].t3 123.463
R19087 BIT_SEL[13].n6 BIT_SEL[13].t4 118.037
R19088 BIT_SEL[13] BIT_SEL[13].n0 7.20211
R19089 BIT_SEL[13].n0 BIT_SEL[13] 5.42621
R19090 BIT_SEL[13] BIT_SEL[13].n1 7.20211
R19091 BIT_SEL[13].n1 BIT_SEL[13] 5.42621
R19092 BIT_SEL[13] BIT_SEL[13].n2 7.20211
R19093 BIT_SEL[13].n2 BIT_SEL[13] 5.42621
R19094 BIT_SEL[13] BIT_SEL[13].n3 7.20211
R19095 BIT_SEL[13].n3 BIT_SEL[13] 5.42621
R19096 BIT_SEL[13] BIT_SEL[13].n4 7.20211
R19097 BIT_SEL[13].n4 BIT_SEL[13] 5.42621
R19098 BIT_SEL[13] BIT_SEL[13].n5 7.20211
R19099 BIT_SEL[13].n5 BIT_SEL[13] 5.42621
R19100 BIT_SEL[13].t0 BIT_SEL[13].n5 118.037
R19101 BIT_SEL[13].t6 BIT_SEL[13].n4 118.037
R19102 BIT_SEL[13].t5 BIT_SEL[13].n3 118.037
R19103 BIT_SEL[13].t2 BIT_SEL[13].n2 118.037
R19104 BIT_SEL[13].t1 BIT_SEL[13].n1 118.037
R19105 BIT_SEL[13].t7 BIT_SEL[13].n0 118.037
R19106 a_1340_55763.t0 a_1340_55763.t1 8.49425
R19107 BIT_SEL[16].n6 BIT_SEL[16] 11.2666
R19108 BIT_SEL[16] BIT_SEL[16].n6 1.36175
R19109 BIT_SEL[16].n6 BIT_SEL[16].t3 115.474
R19110 BIT_SEL[16] BIT_SEL[16].n0 1.36175
R19111 BIT_SEL[16].n0 BIT_SEL[16] 11.2666
R19112 BIT_SEL[16] BIT_SEL[16].n1 1.36175
R19113 BIT_SEL[16].n1 BIT_SEL[16] 11.2666
R19114 BIT_SEL[16] BIT_SEL[16].n2 1.36175
R19115 BIT_SEL[16].n2 BIT_SEL[16] 11.2666
R19116 BIT_SEL[16] BIT_SEL[16].n3 1.36175
R19117 BIT_SEL[16].n3 BIT_SEL[16] 11.2666
R19118 BIT_SEL[16] BIT_SEL[16].n4 1.36175
R19119 BIT_SEL[16].n4 BIT_SEL[16] 11.2666
R19120 BIT_SEL[16] BIT_SEL[16].n5 1.36175
R19121 BIT_SEL[16].n5 BIT_SEL[16] 11.2666
R19122 BIT_SEL[16].t4 BIT_SEL[16] 116.835
R19123 BIT_SEL[16].t7 BIT_SEL[16].n5 115.474
R19124 BIT_SEL[16].t1 BIT_SEL[16].n4 115.474
R19125 BIT_SEL[16].t6 BIT_SEL[16].n3 115.474
R19126 BIT_SEL[16].t5 BIT_SEL[16].n2 115.474
R19127 BIT_SEL[16].t2 BIT_SEL[16].n1 115.474
R19128 BIT_SEL[16].t0 BIT_SEL[16].n0 115.474
R19129 a_7738_11958.t0 a_7738_11958.t1 6.66648
R19130 a_7830_31764.t0 a_7830_31764.t1 9.52407
R19131 a_154_31145.t0 a_154_31145.t1 13.9628
R19132 a_110_31233.t0 a_110_31233.t1 19.5535
R19133 a_14320_20781.t0 a_14320_20781.t1 8.02156
R19134 BIT_SEL[5].t6 BIT_SEL[5] 118.936
R19135 BIT_SEL[5] BIT_SEL[5].n0 10.0837
R19136 BIT_SEL[5] BIT_SEL[5].n0 2.54461
R19137 BIT_SEL[5] BIT_SEL[5].n1 10.0837
R19138 BIT_SEL[5].n1 BIT_SEL[5] 2.54461
R19139 BIT_SEL[5] BIT_SEL[5].n2 10.0837
R19140 BIT_SEL[5].n2 BIT_SEL[5] 2.54461
R19141 BIT_SEL[5] BIT_SEL[5].n3 10.0837
R19142 BIT_SEL[5].n3 BIT_SEL[5] 2.54461
R19143 BIT_SEL[5] BIT_SEL[5].n4 10.0837
R19144 BIT_SEL[5].n4 BIT_SEL[5] 2.54461
R19145 BIT_SEL[5] BIT_SEL[5].n5 10.0837
R19146 BIT_SEL[5].n5 BIT_SEL[5] 2.54461
R19147 BIT_SEL[5] BIT_SEL[5].n6 10.0837
R19148 BIT_SEL[5].n6 BIT_SEL[5] 2.54461
R19149 BIT_SEL[5].t7 BIT_SEL[5].n6 116.391
R19150 BIT_SEL[5].t4 BIT_SEL[5].n5 116.391
R19151 BIT_SEL[5].t2 BIT_SEL[5].n4 116.391
R19152 BIT_SEL[5].t0 BIT_SEL[5].n3 116.391
R19153 BIT_SEL[5].t5 BIT_SEL[5].n2 116.391
R19154 BIT_SEL[5].n1 BIT_SEL[5].t1 116.391
R19155 BIT_SEL[5].n0 BIT_SEL[5].t3 116.391
R19156 a_1340_33925.t0 a_1340_33925.t1 6.71904
R19157 a_110_32838.t0 a_110_32838.t1 19.5535
R19158 a_154_32750.t0 a_154_32750.t1 13.9628
R19159 BIT_SEL[42].n6 BIT_SEL[42] 8.05068
R19160 BIT_SEL[42] BIT_SEL[42].n6 4.57764
R19161 BIT_SEL[42].n6 BIT_SEL[42].t6 117.419
R19162 BIT_SEL[42] BIT_SEL[42].n0 4.57764
R19163 BIT_SEL[42].n0 BIT_SEL[42] 8.05068
R19164 BIT_SEL[42] BIT_SEL[42].n1 4.57764
R19165 BIT_SEL[42].n1 BIT_SEL[42] 8.05068
R19166 BIT_SEL[42] BIT_SEL[42].n2 4.57764
R19167 BIT_SEL[42].n2 BIT_SEL[42] 8.05068
R19168 BIT_SEL[42] BIT_SEL[42].n3 4.57764
R19169 BIT_SEL[42].n3 BIT_SEL[42] 8.05068
R19170 BIT_SEL[42] BIT_SEL[42].n4 4.57764
R19171 BIT_SEL[42].n4 BIT_SEL[42] 8.05068
R19172 BIT_SEL[42] BIT_SEL[42].n5 4.57764
R19173 BIT_SEL[42].n5 BIT_SEL[42] 8.05068
R19174 BIT_SEL[42].t4 BIT_SEL[42] 121.998
R19175 BIT_SEL[42].t3 BIT_SEL[42].n5 117.419
R19176 BIT_SEL[42].t1 BIT_SEL[42].n4 117.419
R19177 BIT_SEL[42].t7 BIT_SEL[42].n3 117.419
R19178 BIT_SEL[42].t5 BIT_SEL[42].n2 117.419
R19179 BIT_SEL[42].t2 BIT_SEL[42].n1 117.419
R19180 BIT_SEL[42].t0 BIT_SEL[42].n0 117.419
R19181 a_14320_14537.t0 a_14320_14537.t1 6.9546
R19182 a_110_58341.t0 a_110_58341.n4 4.88081
R19183 a_110_58341.n4 a_110_58341.n5 2.6905
R19184 a_110_58341.n5 a_110_58341.t1 2.06607
R19185 a_110_58341.n5 a_110_58341.t2 2.2382
R19186 a_110_58341.n4 a_110_58341.n0 0.766047
R19187 a_110_58341.n0 a_110_58341.t3 8.68401
R19188 a_110_58341.n2 a_110_58341.n3 5.21793
R19189 a_110_58341.n0 a_110_58341.n2 4.76793
R19190 a_110_58341.n3 a_110_58341.t4 8.51897
R19191 a_110_58341.n3 a_110_58341.t5 4.4523
R19192 a_110_58341.n2 a_110_58341.n1 8.53373
R19193 a_110_58341.n1 a_110_58341.t7 12.3497
R19194 a_110_58341.n1 a_110_58341.t6 17.192
R19195 a_110_57445.t0 a_110_57445.n3 4.44412
R19196 a_110_57445.n3 a_110_57445.n0 0.1805
R19197 a_110_57445.n3 a_110_57445.n2 4.47779
R19198 a_110_57445.n2 a_110_57445.t3 12.3497
R19199 a_110_57445.n2 a_110_57445.t4 17.192
R19200 a_110_57445.n0 a_110_57445.n1 14.1624
R19201 a_110_57445.n1 a_110_57445.t5 12.3497
R19202 a_110_57445.n1 a_110_57445.t2 17.192
R19203 a_110_57445.n0 a_110_57445.t1 8.34715
R19204 BIT_SEL[9].t0 BIT_SEL[9] 121.198
R19205 BIT_SEL[9] BIT_SEL[9].n0 8.64371
R19206 BIT_SEL[9] BIT_SEL[9].n0 3.98461
R19207 BIT_SEL[9] BIT_SEL[9].n1 8.64371
R19208 BIT_SEL[9].n1 BIT_SEL[9] 3.98461
R19209 BIT_SEL[9] BIT_SEL[9].n2 8.64371
R19210 BIT_SEL[9].n2 BIT_SEL[9] 3.98461
R19211 BIT_SEL[9] BIT_SEL[9].n3 8.64371
R19212 BIT_SEL[9].n3 BIT_SEL[9] 3.98461
R19213 BIT_SEL[9] BIT_SEL[9].n4 8.64371
R19214 BIT_SEL[9].n4 BIT_SEL[9] 3.98461
R19215 BIT_SEL[9] BIT_SEL[9].n5 8.64371
R19216 BIT_SEL[9].n5 BIT_SEL[9] 3.98461
R19217 BIT_SEL[9] BIT_SEL[9].n6 8.64371
R19218 BIT_SEL[9].n6 BIT_SEL[9] 3.98461
R19219 BIT_SEL[9].t4 BIT_SEL[9].n6 117.215
R19220 BIT_SEL[9].t2 BIT_SEL[9].n5 117.215
R19221 BIT_SEL[9].t6 BIT_SEL[9].n4 117.215
R19222 BIT_SEL[9].t1 BIT_SEL[9].n3 117.215
R19223 BIT_SEL[9].t5 BIT_SEL[9].n2 117.215
R19224 BIT_SEL[9].n1 BIT_SEL[9].t3 117.215
R19225 BIT_SEL[9].n0 BIT_SEL[9].t7 117.215
R19226 a_1340_1521.t0 a_1340_1521.t1 6.39548
R19227 a_14320_36535.t0 a_14320_36535.t1 8.02156
R19228 BIT_SEL[55].n6 BIT_SEL[55] 3.39318
R19229 BIT_SEL[55] BIT_SEL[55].n6 9.23514
R19230 BIT_SEL[55] BIT_SEL[55].t3 120.195
R19231 BIT_SEL[55].n6 BIT_SEL[55].t1 116.802
R19232 BIT_SEL[55] BIT_SEL[55].n0 9.23514
R19233 BIT_SEL[55].n0 BIT_SEL[55] 3.39318
R19234 BIT_SEL[55] BIT_SEL[55].n1 9.23514
R19235 BIT_SEL[55].n1 BIT_SEL[55] 3.39318
R19236 BIT_SEL[55] BIT_SEL[55].n2 9.23514
R19237 BIT_SEL[55].n2 BIT_SEL[55] 3.39318
R19238 BIT_SEL[55] BIT_SEL[55].n3 9.23514
R19239 BIT_SEL[55].n3 BIT_SEL[55] 3.39318
R19240 BIT_SEL[55] BIT_SEL[55].n4 9.23514
R19241 BIT_SEL[55].n4 BIT_SEL[55] 3.39318
R19242 BIT_SEL[55] BIT_SEL[55].n5 9.23514
R19243 BIT_SEL[55].n5 BIT_SEL[55] 3.39318
R19244 BIT_SEL[55].t2 BIT_SEL[55].n5 116.802
R19245 BIT_SEL[55].t5 BIT_SEL[55].n4 116.802
R19246 BIT_SEL[55].t0 BIT_SEL[55].n3 116.802
R19247 BIT_SEL[55].t7 BIT_SEL[55].n2 116.802
R19248 BIT_SEL[55].t6 BIT_SEL[55].n1 116.802
R19249 BIT_SEL[55].t4 BIT_SEL[55].n0 116.802
R19250 a_20810_41274.t0 a_20810_41274.t1 5.92075
R19251 BIT_SEL[32] BIT_SEL[32].n0 1.36175
R19252 BIT_SEL[32] BIT_SEL[32].n0 11.2666
R19253 BIT_SEL[32] BIT_SEL[32].n1 1.36175
R19254 BIT_SEL[32].n1 BIT_SEL[32] 11.2666
R19255 BIT_SEL[32] BIT_SEL[32].n2 1.36175
R19256 BIT_SEL[32].n2 BIT_SEL[32] 11.2666
R19257 BIT_SEL[32] BIT_SEL[32].n3 1.36175
R19258 BIT_SEL[32].n3 BIT_SEL[32] 11.2666
R19259 BIT_SEL[32] BIT_SEL[32].n4 1.36175
R19260 BIT_SEL[32].n4 BIT_SEL[32] 11.2666
R19261 BIT_SEL[32] BIT_SEL[32].n5 1.36175
R19262 BIT_SEL[32].n5 BIT_SEL[32] 11.2666
R19263 BIT_SEL[32] BIT_SEL[32].n6 1.36175
R19264 BIT_SEL[32].n6 BIT_SEL[32] 11.2666
R19265 BIT_SEL[32].t1 BIT_SEL[32] 116.835
R19266 BIT_SEL[32].t4 BIT_SEL[32].n6 115.474
R19267 BIT_SEL[32].t6 BIT_SEL[32].n5 115.474
R19268 BIT_SEL[32].t3 BIT_SEL[32].n4 115.474
R19269 BIT_SEL[32].t2 BIT_SEL[32].n3 115.474
R19270 BIT_SEL[32].t7 BIT_SEL[32].n2 115.474
R19271 BIT_SEL[32].n1 BIT_SEL[32].t5 115.474
R19272 BIT_SEL[32].n0 BIT_SEL[32].t0 115.474
R19273 a_1340_13272.t0 a_1340_13272.t1 7.18327
R19274 a_14320_60166.t0 a_14320_60166.t1 8.02156
R19275 a_110_54864.t0 a_110_54864.t1 19.5535
R19276 a_154_54776.t0 a_154_54776.t1 13.9628
R19277 a_14320_58293.t0 a_14320_58293.t1 6.02155
R19278 PRESET_N.n2 PRESET_N 0.008
R19279 PRESET_N PRESET_N.n20 0.008
R19280 PRESET_N PRESET_N.n2 12.6253
R19281 PRESET_N PRESET_N.n20 12.6253
R19282 PRESET_N.n22 PRESET_N.n21 0.2555
R19283 PRESET_N.n21 PRESET_N 5.13582
R19284 PRESET_N.t21 PRESET_N.n22 21.3045
R19285 PRESET_N.t16 PRESET_N.n22 20.9945
R19286 PRESET_N.t12 PRESET_N.n21 20.9945
R19287 PRESET_N.n18 PRESET_N.n19 0.2555
R19288 PRESET_N.n20 PRESET_N.n18 5.12832
R19289 PRESET_N.n19 PRESET_N.t14 21.3045
R19290 PRESET_N.n19 PRESET_N.t11 20.9945
R19291 PRESET_N.n18 PRESET_N.t3 20.9945
R19292 PRESET_N PRESET_N.n5 12.6253
R19293 PRESET_N.n5 PRESET_N 0.008
R19294 PRESET_N PRESET_N.n8 12.6253
R19295 PRESET_N.n8 PRESET_N 0.008
R19296 PRESET_N PRESET_N.n11 12.6253
R19297 PRESET_N.n11 PRESET_N 0.008
R19298 PRESET_N PRESET_N.n14 12.6253
R19299 PRESET_N.n14 PRESET_N 0.008
R19300 PRESET_N PRESET_N.n17 12.6253
R19301 PRESET_N.n17 PRESET_N 0.008
R19302 PRESET_N.n16 PRESET_N.n15 0.2555
R19303 PRESET_N.n15 PRESET_N.n17 5.12832
R19304 PRESET_N.t5 PRESET_N.n16 21.3045
R19305 PRESET_N.t23 PRESET_N.n16 20.9945
R19306 PRESET_N.t17 PRESET_N.n15 20.9945
R19307 PRESET_N.n13 PRESET_N.n12 0.2555
R19308 PRESET_N.n12 PRESET_N.n14 5.12832
R19309 PRESET_N.t10 PRESET_N.n13 21.3045
R19310 PRESET_N.t8 PRESET_N.n13 20.9945
R19311 PRESET_N.t9 PRESET_N.n12 20.9945
R19312 PRESET_N.n10 PRESET_N.n9 0.2555
R19313 PRESET_N.n9 PRESET_N.n11 5.12832
R19314 PRESET_N.t7 PRESET_N.n10 21.3045
R19315 PRESET_N.t2 PRESET_N.n10 20.9945
R19316 PRESET_N.t4 PRESET_N.n9 20.9945
R19317 PRESET_N.n7 PRESET_N.n6 0.2555
R19318 PRESET_N.n6 PRESET_N.n8 5.12832
R19319 PRESET_N.t13 PRESET_N.n7 21.3045
R19320 PRESET_N.t0 PRESET_N.n7 20.9945
R19321 PRESET_N.t20 PRESET_N.n6 20.9945
R19322 PRESET_N.n4 PRESET_N.n3 0.2555
R19323 PRESET_N.n3 PRESET_N.n5 5.12832
R19324 PRESET_N.t6 PRESET_N.n4 21.3045
R19325 PRESET_N.t22 PRESET_N.n4 20.9945
R19326 PRESET_N.t15 PRESET_N.n3 20.9945
R19327 PRESET_N.n0 PRESET_N.n1 0.2555
R19328 PRESET_N.n2 PRESET_N.n0 5.12832
R19329 PRESET_N.n1 PRESET_N.t1 21.3045
R19330 PRESET_N.n1 PRESET_N.t18 20.9945
R19331 PRESET_N.n0 PRESET_N.t19 20.9945
R19332 BIT_SEL[12].n6 BIT_SEL[12] 7.2005
R19333 BIT_SEL[12] BIT_SEL[12].n6 5.42782
R19334 BIT_SEL[12].n6 BIT_SEL[12].t1 117.832
R19335 BIT_SEL[12] BIT_SEL[12].n0 5.42782
R19336 BIT_SEL[12].n0 BIT_SEL[12] 7.2005
R19337 BIT_SEL[12] BIT_SEL[12].n1 5.42782
R19338 BIT_SEL[12].n1 BIT_SEL[12] 7.2005
R19339 BIT_SEL[12] BIT_SEL[12].n2 5.42782
R19340 BIT_SEL[12].n2 BIT_SEL[12] 7.2005
R19341 BIT_SEL[12] BIT_SEL[12].n3 5.42782
R19342 BIT_SEL[12].n3 BIT_SEL[12] 7.2005
R19343 BIT_SEL[12] BIT_SEL[12].n4 5.42782
R19344 BIT_SEL[12].n4 BIT_SEL[12] 7.2005
R19345 BIT_SEL[12] BIT_SEL[12].n5 5.42782
R19346 BIT_SEL[12].n5 BIT_SEL[12] 7.2005
R19347 BIT_SEL[12].t6 BIT_SEL[12] 123.258
R19348 BIT_SEL[12].t3 BIT_SEL[12].n5 117.832
R19349 BIT_SEL[12].t5 BIT_SEL[12].n4 117.832
R19350 BIT_SEL[12].t2 BIT_SEL[12].n3 117.832
R19351 BIT_SEL[12].t4 BIT_SEL[12].n2 117.832
R19352 BIT_SEL[12].t0 BIT_SEL[12].n1 117.832
R19353 BIT_SEL[12].t7 BIT_SEL[12].n0 117.832
R19354 a_1340_22943.t0 a_1340_22943.t1 8.02468
R19355 a_110_48592.t0 a_110_48592.t1 19.5535
R19356 a_154_48504.t0 a_154_48504.t1 13.9628
R19357 BIT_SEL[63].t5 BIT_SEL[63] 124.466
R19358 BIT_SEL[63] BIT_SEL[63].n0 6.61068
R19359 BIT_SEL[63] BIT_SEL[63].n0 6.01764
R19360 BIT_SEL[63] BIT_SEL[63].n1 6.61068
R19361 BIT_SEL[63].n1 BIT_SEL[63] 6.01764
R19362 BIT_SEL[63] BIT_SEL[63].n2 6.61068
R19363 BIT_SEL[63].n2 BIT_SEL[63] 6.01764
R19364 BIT_SEL[63] BIT_SEL[63].n3 6.61068
R19365 BIT_SEL[63].n3 BIT_SEL[63] 6.01764
R19366 BIT_SEL[63] BIT_SEL[63].n4 6.61068
R19367 BIT_SEL[63].n4 BIT_SEL[63] 6.01764
R19368 BIT_SEL[63] BIT_SEL[63].n5 6.61068
R19369 BIT_SEL[63].n5 BIT_SEL[63] 6.01764
R19370 BIT_SEL[63] BIT_SEL[63].n6 6.61068
R19371 BIT_SEL[63].n6 BIT_SEL[63] 6.01764
R19372 BIT_SEL[63].t4 BIT_SEL[63].n6 118.448
R19373 BIT_SEL[63].t2 BIT_SEL[63].n5 118.448
R19374 BIT_SEL[63].t1 BIT_SEL[63].n4 118.448
R19375 BIT_SEL[63].t7 BIT_SEL[63].n3 118.448
R19376 BIT_SEL[63].t3 BIT_SEL[63].n2 118.448
R19377 BIT_SEL[63].n1 BIT_SEL[63].t6 118.448
R19378 BIT_SEL[63].n0 BIT_SEL[63].t0 118.448
R19379 a_20810_8133.t0 a_20810_8133.t1 9.52293
R19380 a_7830_17643.t0 a_7830_17643.t1 5.92117
R19381 BIT_SEL[36] BIT_SEL[36].n0 2.54461
R19382 BIT_SEL[36] BIT_SEL[36].n0 10.0837
R19383 BIT_SEL[36] BIT_SEL[36].n1 2.54461
R19384 BIT_SEL[36].n1 BIT_SEL[36] 10.0837
R19385 BIT_SEL[36] BIT_SEL[36].n2 2.54461
R19386 BIT_SEL[36].n2 BIT_SEL[36] 10.0837
R19387 BIT_SEL[36] BIT_SEL[36].n3 2.54461
R19388 BIT_SEL[36].n3 BIT_SEL[36] 10.0837
R19389 BIT_SEL[36] BIT_SEL[36].n4 2.54461
R19390 BIT_SEL[36].n4 BIT_SEL[36] 10.0837
R19391 BIT_SEL[36] BIT_SEL[36].n5 2.54461
R19392 BIT_SEL[36].n5 BIT_SEL[36] 10.0837
R19393 BIT_SEL[36] BIT_SEL[36].n6 2.54461
R19394 BIT_SEL[36].n6 BIT_SEL[36] 10.0837
R19395 BIT_SEL[36].t0 BIT_SEL[36] 118.73
R19396 BIT_SEL[36].t6 BIT_SEL[36].n6 116.186
R19397 BIT_SEL[36].t4 BIT_SEL[36].n5 116.186
R19398 BIT_SEL[36].t5 BIT_SEL[36].n4 116.186
R19399 BIT_SEL[36].t3 BIT_SEL[36].n3 116.186
R19400 BIT_SEL[36].t7 BIT_SEL[36].n2 116.186
R19401 BIT_SEL[36].n1 BIT_SEL[36].t1 116.186
R19402 BIT_SEL[36].n0 BIT_SEL[36].t2 116.186
R19403 a_14320_60534.t0 a_14320_60534.t1 7.18327
R19404 a_20810_13801.t0 a_20810_13801.t1 6.38524
R19405 a_14320_46045.t0 a_14320_46045.t1 6.9546
R19406 a_1340_29026.t0 a_1340_29026.t1 7.18213
R19407 a_110_9207.t0 a_110_9207.t1 19.5535
R19408 a_154_9119.t0 a_154_9119.t1 13.9628
R19409 BIT_SEL[18] BIT_SEL[18].n0 1.95318
R19410 BIT_SEL[18] BIT_SEL[18].n0 10.6751
R19411 BIT_SEL[18] BIT_SEL[18].n1 1.95318
R19412 BIT_SEL[18].n1 BIT_SEL[18] 10.6751
R19413 BIT_SEL[18] BIT_SEL[18].n2 1.95318
R19414 BIT_SEL[18].n2 BIT_SEL[18] 10.6751
R19415 BIT_SEL[18] BIT_SEL[18].n3 1.95318
R19416 BIT_SEL[18].n3 BIT_SEL[18] 10.6751
R19417 BIT_SEL[18] BIT_SEL[18].n4 1.95318
R19418 BIT_SEL[18].n4 BIT_SEL[18] 10.6751
R19419 BIT_SEL[18] BIT_SEL[18].n5 1.95318
R19420 BIT_SEL[18].n5 BIT_SEL[18] 10.6751
R19421 BIT_SEL[18] BIT_SEL[18].n6 1.95318
R19422 BIT_SEL[18].n6 BIT_SEL[18] 10.6751
R19423 BIT_SEL[18].t4 BIT_SEL[18] 117.727
R19424 BIT_SEL[18].t2 BIT_SEL[18].n6 115.775
R19425 BIT_SEL[18].t0 BIT_SEL[18].n5 115.775
R19426 BIT_SEL[18].t7 BIT_SEL[18].n4 115.775
R19427 BIT_SEL[18].t6 BIT_SEL[18].n3 115.775
R19428 BIT_SEL[18].t1 BIT_SEL[18].n2 115.775
R19429 BIT_SEL[18].n1 BIT_SEL[18].t3 115.775
R19430 BIT_SEL[18].n0 BIT_SEL[18].t5 115.775
R19431 a_7830_44412.t0 a_7830_44412.t1 8.02269
R19432 a_20810_62328.t0 a_20810_62328.t1 8.02468
R19433 a_7830_33397.t0 a_7830_33397.t1 5.92117
R19434 a_1340_24255.t0 a_1340_24255.t1 8.49425
R19435 BIT_SEL[0].n6 BIT_SEL[0] 11.2666
R19436 BIT_SEL[0] BIT_SEL[0].n6 1.36175
R19437 BIT_SEL[0].n6 BIT_SEL[0].t7 115.474
R19438 BIT_SEL[0] BIT_SEL[0].n0 1.36175
R19439 BIT_SEL[0].n0 BIT_SEL[0] 11.2666
R19440 BIT_SEL[0] BIT_SEL[0].n1 1.36175
R19441 BIT_SEL[0].n1 BIT_SEL[0] 11.2666
R19442 BIT_SEL[0] BIT_SEL[0].n2 1.36175
R19443 BIT_SEL[0].n2 BIT_SEL[0] 11.2666
R19444 BIT_SEL[0] BIT_SEL[0].n3 1.36175
R19445 BIT_SEL[0].n3 BIT_SEL[0] 11.2666
R19446 BIT_SEL[0] BIT_SEL[0].n4 1.36175
R19447 BIT_SEL[0].n4 BIT_SEL[0] 11.2666
R19448 BIT_SEL[0] BIT_SEL[0].n5 1.36175
R19449 BIT_SEL[0].n5 BIT_SEL[0] 11.2666
R19450 BIT_SEL[0].t0 BIT_SEL[0] 116.835
R19451 BIT_SEL[0].t3 BIT_SEL[0].n5 115.474
R19452 BIT_SEL[0].t5 BIT_SEL[0].n4 115.474
R19453 BIT_SEL[0].t2 BIT_SEL[0].n3 115.474
R19454 BIT_SEL[0].t1 BIT_SEL[0].n2 115.474
R19455 BIT_SEL[0].t6 BIT_SEL[0].n1 115.474
R19456 BIT_SEL[0].t4 BIT_SEL[0].n0 115.474
R19457 BIT_SEL[35].t3 BIT_SEL[35] 117.93
R19458 BIT_SEL[35] BIT_SEL[35].n0 10.6768
R19459 BIT_SEL[35] BIT_SEL[35].n0 1.95157
R19460 BIT_SEL[35] BIT_SEL[35].n1 10.6768
R19461 BIT_SEL[35].n1 BIT_SEL[35] 1.95157
R19462 BIT_SEL[35] BIT_SEL[35].n2 10.6768
R19463 BIT_SEL[35].n2 BIT_SEL[35] 1.95157
R19464 BIT_SEL[35] BIT_SEL[35].n3 10.6768
R19465 BIT_SEL[35].n3 BIT_SEL[35] 1.95157
R19466 BIT_SEL[35] BIT_SEL[35].n4 10.6768
R19467 BIT_SEL[35].n4 BIT_SEL[35] 1.95157
R19468 BIT_SEL[35] BIT_SEL[35].n5 10.6768
R19469 BIT_SEL[35].n5 BIT_SEL[35] 1.95157
R19470 BIT_SEL[35] BIT_SEL[35].n6 10.6768
R19471 BIT_SEL[35].n6 BIT_SEL[35] 1.95157
R19472 BIT_SEL[35].t5 BIT_SEL[35].n6 115.98
R19473 BIT_SEL[35].t4 BIT_SEL[35].n5 115.98
R19474 BIT_SEL[35].t2 BIT_SEL[35].n4 115.98
R19475 BIT_SEL[35].t0 BIT_SEL[35].n3 115.98
R19476 BIT_SEL[35].t7 BIT_SEL[35].n2 115.98
R19477 BIT_SEL[35].n1 BIT_SEL[35].t6 115.98
R19478 BIT_SEL[35].n0 BIT_SEL[35].t1 115.98
R19479 a_14320_34294.t0 a_14320_34294.t1 7.55862
R19480 a_7830_6660.t0 a_7830_6660.t1 6.95418
R19481 SENSE.n5 SENSE 0.0620789
R19482 SENSE.n5 SENSE.n0 12.5378
R19483 SENSE.n4 SENSE.n5 12.5378
R19484 SENSE SENSE.n4 0.0620789
R19485 SENSE SENSE.t1 21.0993
R19486 SENSE.n4 SENSE.n3 12.5378
R19487 SENSE.n3 SENSE 0.0620789
R19488 SENSE SENSE.t5 21.0993
R19489 SENSE.n3 SENSE.n2 12.5378
R19490 SENSE.n2 SENSE 0.0620789
R19491 SENSE SENSE.t2 21.0993
R19492 SENSE.n2 SENSE.n1 12.5378
R19493 SENSE.n1 SENSE 0.0620789
R19494 SENSE SENSE.t4 21.0993
R19495 SENSE.n1 SENSE 12.5994
R19496 SENSE SENSE.t0 21.0993
R19497 SENSE.n0 SENSE 0.0620789
R19498 SENSE SENSE.t6 21.0993
R19499 SENSE.n0 SENSE 12.5994
R19500 SENSE SENSE.t3 21.0993
R19501 SENSE SENSE.t7 21.0993
R19502 a_1340_44780.t0 a_1340_44780.t1 7.18213
R19503 OUT[4] OUT[4].n0 9.0005
R19504 OUT[4].n0 OUT[4].t1 8.56064
R19505 OUT[4].n0 OUT[4].t0 4.38216
R19506 a_154_1242.t0 a_154_1242.t1 13.9628
R19507 a_110_1330.t0 a_110_1330.t1 19.5535
R19508 BIT_SEL[33].t3 BIT_SEL[33] 116.918
R19509 BIT_SEL[33] BIT_SEL[33].n0 11.2682
R19510 BIT_SEL[33] BIT_SEL[33].n0 1.36014
R19511 BIT_SEL[33] BIT_SEL[33].n1 11.2682
R19512 BIT_SEL[33].n1 BIT_SEL[33] 1.36014
R19513 BIT_SEL[33] BIT_SEL[33].n2 11.2682
R19514 BIT_SEL[33].n2 BIT_SEL[33] 1.36014
R19515 BIT_SEL[33] BIT_SEL[33].n3 11.2682
R19516 BIT_SEL[33].n3 BIT_SEL[33] 1.36014
R19517 BIT_SEL[33] BIT_SEL[33].n4 11.2682
R19518 BIT_SEL[33].n4 BIT_SEL[33] 1.36014
R19519 BIT_SEL[33] BIT_SEL[33].n5 11.2682
R19520 BIT_SEL[33].n5 BIT_SEL[33] 1.36014
R19521 BIT_SEL[33] BIT_SEL[33].n6 11.2682
R19522 BIT_SEL[33].n6 BIT_SEL[33] 1.36014
R19523 BIT_SEL[33].t7 BIT_SEL[33].n6 115.558
R19524 BIT_SEL[33].t2 BIT_SEL[33].n5 115.558
R19525 BIT_SEL[33].t6 BIT_SEL[33].n4 115.558
R19526 BIT_SEL[33].t0 BIT_SEL[33].n3 115.558
R19527 BIT_SEL[33].t5 BIT_SEL[33].n2 115.558
R19528 BIT_SEL[33].n1 BIT_SEL[33].t4 115.558
R19529 BIT_SEL[33].n0 BIT_SEL[33].t1 115.558
R19530 a_14320_34662.t0 a_14320_34662.t1 6.02155
R19531 a_14320_53554.t0 a_14320_53554.t1 5.92569
R19532 a_110_23356.t0 a_110_23356.t1 19.5535
R19533 a_154_23268.t0 a_154_23268.t1 13.9628
R19534 a_14320_13272.t0 a_14320_13272.t1 7.18327
R19535 a_20810_45309.t0 a_20810_45309.t1 6.38411
R19536 a_110_42587.n0 a_110_42587.t0 2.06607
R19537 a_110_42587.t2 a_110_42587.n0 2.2382
R19538 a_110_42587.n0 a_110_42587.n5 2.6905
R19539 a_110_42587.n5 a_110_42587.t1 4.88081
R19540 a_110_42587.n5 a_110_42587.n1 0.766047
R19541 a_110_42587.n1 a_110_42587.t5 8.68401
R19542 a_110_42587.n3 a_110_42587.n4 5.21793
R19543 a_110_42587.n1 a_110_42587.n3 4.76793
R19544 a_110_42587.n4 a_110_42587.t4 8.51897
R19545 a_110_42587.n4 a_110_42587.t3 4.4523
R19546 a_110_42587.n3 a_110_42587.n2 8.53373
R19547 a_110_42587.n2 a_110_42587.t6 12.3497
R19548 a_110_42587.n2 a_110_42587.t7 17.192
R19549 a_110_41691.t0 a_110_41691.n3 4.44412
R19550 a_110_41691.n3 a_110_41691.n0 0.1805
R19551 a_110_41691.n3 a_110_41691.n2 4.47779
R19552 a_110_41691.n2 a_110_41691.t3 12.3497
R19553 a_110_41691.n2 a_110_41691.t5 17.192
R19554 a_110_41691.n0 a_110_41691.n1 14.1624
R19555 a_110_41691.n1 a_110_41691.t2 12.3497
R19556 a_110_41691.n1 a_110_41691.t4 17.192
R19557 a_110_41691.n0 a_110_41691.t1 8.34715
R19558 a_1340_18171.t0 a_1340_18171.t1 6.71904
R19559 BIT_SEL[19].t6 BIT_SEL[19] 117.93
R19560 BIT_SEL[19] BIT_SEL[19].n0 10.6768
R19561 BIT_SEL[19] BIT_SEL[19].n0 1.95157
R19562 BIT_SEL[19] BIT_SEL[19].n1 10.6768
R19563 BIT_SEL[19].n1 BIT_SEL[19] 1.95157
R19564 BIT_SEL[19] BIT_SEL[19].n2 10.6768
R19565 BIT_SEL[19].n2 BIT_SEL[19] 1.95157
R19566 BIT_SEL[19] BIT_SEL[19].n3 10.6768
R19567 BIT_SEL[19].n3 BIT_SEL[19] 1.95157
R19568 BIT_SEL[19] BIT_SEL[19].n4 10.6768
R19569 BIT_SEL[19].n4 BIT_SEL[19] 1.95157
R19570 BIT_SEL[19] BIT_SEL[19].n5 10.6768
R19571 BIT_SEL[19].n5 BIT_SEL[19] 1.95157
R19572 BIT_SEL[19] BIT_SEL[19].n6 10.6768
R19573 BIT_SEL[19].n6 BIT_SEL[19] 1.95157
R19574 BIT_SEL[19].t7 BIT_SEL[19].n6 115.98
R19575 BIT_SEL[19].t5 BIT_SEL[19].n5 115.98
R19576 BIT_SEL[19].t4 BIT_SEL[19].n4 115.98
R19577 BIT_SEL[19].t2 BIT_SEL[19].n3 115.98
R19578 BIT_SEL[19].t1 BIT_SEL[19].n2 115.98
R19579 BIT_SEL[19].n1 BIT_SEL[19].t0 115.98
R19580 BIT_SEL[19].n0 BIT_SEL[19].t3 115.98
R19581 a_7830_18540.t0 a_7830_18540.t1 7.5582
R19582 a_14320_16378.t0 a_14320_16378.t1 8.49538
R19583 a_110_17084.t0 a_110_17084.t1 19.5535
R19584 a_154_16996.t0 a_154_16996.t1 13.9628
R19585 a_20810_45677.t0 a_20810_45677.t1 5.92569
R19586 BIT_SEL[21].t3 BIT_SEL[21] 118.936
R19587 BIT_SEL[21] BIT_SEL[21].n0 10.0837
R19588 BIT_SEL[21] BIT_SEL[21].n0 2.54461
R19589 BIT_SEL[21] BIT_SEL[21].n1 10.0837
R19590 BIT_SEL[21].n1 BIT_SEL[21] 2.54461
R19591 BIT_SEL[21] BIT_SEL[21].n2 10.0837
R19592 BIT_SEL[21].n2 BIT_SEL[21] 2.54461
R19593 BIT_SEL[21] BIT_SEL[21].n3 10.0837
R19594 BIT_SEL[21].n3 BIT_SEL[21] 2.54461
R19595 BIT_SEL[21] BIT_SEL[21].n4 10.0837
R19596 BIT_SEL[21].n4 BIT_SEL[21] 2.54461
R19597 BIT_SEL[21] BIT_SEL[21].n5 10.0837
R19598 BIT_SEL[21].n5 BIT_SEL[21] 2.54461
R19599 BIT_SEL[21] BIT_SEL[21].n6 10.0837
R19600 BIT_SEL[21].n6 BIT_SEL[21] 2.54461
R19601 BIT_SEL[21].t5 BIT_SEL[21].n6 116.391
R19602 BIT_SEL[21].t2 BIT_SEL[21].n5 116.391
R19603 BIT_SEL[21].t0 BIT_SEL[21].n4 116.391
R19604 BIT_SEL[21].t6 BIT_SEL[21].n3 116.391
R19605 BIT_SEL[21].t4 BIT_SEL[21].n2 116.391
R19606 BIT_SEL[21].n1 BIT_SEL[21].t7 116.391
R19607 BIT_SEL[21].n0 BIT_SEL[21].t1 116.391
R19608 a_7830_41802.t0 a_7830_41802.t1 6.71904
R19609 a_20810_61431.t0 a_20810_61431.t1 5.92569
R19610 a_14320_32132.t0 a_14320_32132.t1 8.49425
R19611 BIT_SEL[10] BIT_SEL[10].n0 4.57764
R19612 BIT_SEL[10] BIT_SEL[10].n0 8.05068
R19613 BIT_SEL[10] BIT_SEL[10].n1 4.57764
R19614 BIT_SEL[10].n1 BIT_SEL[10] 8.05068
R19615 BIT_SEL[10] BIT_SEL[10].n2 4.57764
R19616 BIT_SEL[10].n2 BIT_SEL[10] 8.05068
R19617 BIT_SEL[10] BIT_SEL[10].n3 4.57764
R19618 BIT_SEL[10].n3 BIT_SEL[10] 8.05068
R19619 BIT_SEL[10] BIT_SEL[10].n4 4.57764
R19620 BIT_SEL[10].n4 BIT_SEL[10] 8.05068
R19621 BIT_SEL[10] BIT_SEL[10].n5 4.57764
R19622 BIT_SEL[10].n5 BIT_SEL[10] 8.05068
R19623 BIT_SEL[10] BIT_SEL[10].n6 4.57764
R19624 BIT_SEL[10].n6 BIT_SEL[10] 8.05068
R19625 BIT_SEL[10].t6 BIT_SEL[10] 121.998
R19626 BIT_SEL[10].t5 BIT_SEL[10].n6 117.419
R19627 BIT_SEL[10].t3 BIT_SEL[10].n5 117.419
R19628 BIT_SEL[10].t1 BIT_SEL[10].n4 117.419
R19629 BIT_SEL[10].t7 BIT_SEL[10].n3 117.419
R19630 BIT_SEL[10].t4 BIT_SEL[10].n2 117.419
R19631 BIT_SEL[10].n1 BIT_SEL[10].t2 117.419
R19632 BIT_SEL[10].n0 BIT_SEL[10].t0 117.419
R19633 a_1340_6660.t0 a_1340_6660.t1 6.9546
R19634 a_20810_60534.t0 a_20810_60534.t1 7.18213
R19635 a_154_61757.t0 a_154_61757.t1 13.9628
R19636 a_110_61845.t0 a_110_61845.t1 19.5535
R19637 a_7830_47886.t0 a_7830_47886.t1 8.49425
R19638 a_1248_27712.t0 a_1248_27712.t1 6.66648
R19639 a_154_55485.t0 a_154_55485.t1 13.9628
R19640 a_110_55573.t0 a_110_55573.t1 19.5535
R19641 a_7830_48783.t0 a_7830_48783.t1 6.39662
R19642 BIT_SEL[3].t1 BIT_SEL[3] 117.93
R19643 BIT_SEL[3] BIT_SEL[3].n0 10.6768
R19644 BIT_SEL[3] BIT_SEL[3].n0 1.95157
R19645 BIT_SEL[3] BIT_SEL[3].n1 10.6768
R19646 BIT_SEL[3].n1 BIT_SEL[3] 1.95157
R19647 BIT_SEL[3] BIT_SEL[3].n2 10.6768
R19648 BIT_SEL[3].n2 BIT_SEL[3] 1.95157
R19649 BIT_SEL[3] BIT_SEL[3].n3 10.6768
R19650 BIT_SEL[3].n3 BIT_SEL[3] 1.95157
R19651 BIT_SEL[3] BIT_SEL[3].n4 10.6768
R19652 BIT_SEL[3].n4 BIT_SEL[3] 1.95157
R19653 BIT_SEL[3] BIT_SEL[3].n5 10.6768
R19654 BIT_SEL[3].n5 BIT_SEL[3] 1.95157
R19655 BIT_SEL[3] BIT_SEL[3].n6 10.6768
R19656 BIT_SEL[3].n6 BIT_SEL[3] 1.95157
R19657 BIT_SEL[3].t2 BIT_SEL[3].n6 115.98
R19658 BIT_SEL[3].t0 BIT_SEL[3].n5 115.98
R19659 BIT_SEL[3].t7 BIT_SEL[3].n4 115.98
R19660 BIT_SEL[3].t5 BIT_SEL[3].n3 115.98
R19661 BIT_SEL[3].t4 BIT_SEL[3].n2 115.98
R19662 BIT_SEL[3].n1 BIT_SEL[3].t3 115.98
R19663 BIT_SEL[3].n0 BIT_SEL[3].t6 115.98
R19664 a_1340_50048.t0 a_1340_50048.t1 7.55862
R19665 COL_PROG_N[4] COL_PROG_N[4].n0 0.0965
R19666 COL_PROG_N[4].n0 COL_PROG_N[4].n1 0.3065
R19667 COL_PROG_N[4].n1 COL_PROG_N[4].n2 0.3065
R19668 COL_PROG_N[4].n2 COL_PROG_N[4].t0 292.788
R19669 COL_PROG_N[4].n2 COL_PROG_N[4].t2 292.481
R19670 COL_PROG_N[4].n1 COL_PROG_N[4].t1 292.481
R19671 COL_PROG_N[4].n0 COL_PROG_N[4].t3 292.481
R19672 a_20810_12904.t0 a_20810_12904.t1 8.02269
R19673 BIT_SEL[2] BIT_SEL[2].n0 1.95318
R19674 BIT_SEL[2] BIT_SEL[2].n0 10.6751
R19675 BIT_SEL[2] BIT_SEL[2].n1 1.95318
R19676 BIT_SEL[2].n1 BIT_SEL[2] 10.6751
R19677 BIT_SEL[2] BIT_SEL[2].n2 1.95318
R19678 BIT_SEL[2].n2 BIT_SEL[2] 10.6751
R19679 BIT_SEL[2] BIT_SEL[2].n3 1.95318
R19680 BIT_SEL[2].n3 BIT_SEL[2] 10.6751
R19681 BIT_SEL[2] BIT_SEL[2].n4 1.95318
R19682 BIT_SEL[2].n4 BIT_SEL[2] 10.6751
R19683 BIT_SEL[2] BIT_SEL[2].n5 1.95318
R19684 BIT_SEL[2].n5 BIT_SEL[2] 10.6751
R19685 BIT_SEL[2] BIT_SEL[2].n6 1.95318
R19686 BIT_SEL[2].n6 BIT_SEL[2] 10.6751
R19687 BIT_SEL[2].t6 BIT_SEL[2] 117.727
R19688 BIT_SEL[2].t4 BIT_SEL[2].n6 115.775
R19689 BIT_SEL[2].t2 BIT_SEL[2].n5 115.775
R19690 BIT_SEL[2].t1 BIT_SEL[2].n4 115.775
R19691 BIT_SEL[2].t0 BIT_SEL[2].n3 115.775
R19692 BIT_SEL[2].t3 BIT_SEL[2].n2 115.775
R19693 BIT_SEL[2].n1 BIT_SEL[2].t5 115.775
R19694 BIT_SEL[2].n0 BIT_SEL[2].t7 115.775
R19695 a_1340_28658.t0 a_1340_28658.t1 8.02269
R19696 a_7830_23311.t0 a_7830_23311.t1 9.05337
R19697 a_1340_61799.t0 a_1340_61799.t1 6.9546
R19698 a_14228_51343.t0 a_14228_51343.t1 6.66648
R19699 BIT_SEL[44].n6 BIT_SEL[44] 7.2005
R19700 BIT_SEL[44] BIT_SEL[44].n6 5.42782
R19701 BIT_SEL[44].n6 BIT_SEL[44].t7 117.832
R19702 BIT_SEL[44] BIT_SEL[44].n0 5.42782
R19703 BIT_SEL[44].n0 BIT_SEL[44] 7.2005
R19704 BIT_SEL[44] BIT_SEL[44].n1 5.42782
R19705 BIT_SEL[44].n1 BIT_SEL[44] 7.2005
R19706 BIT_SEL[44] BIT_SEL[44].n2 5.42782
R19707 BIT_SEL[44].n2 BIT_SEL[44] 7.2005
R19708 BIT_SEL[44] BIT_SEL[44].n3 5.42782
R19709 BIT_SEL[44].n3 BIT_SEL[44] 7.2005
R19710 BIT_SEL[44] BIT_SEL[44].n4 5.42782
R19711 BIT_SEL[44].n4 BIT_SEL[44] 7.2005
R19712 BIT_SEL[44] BIT_SEL[44].n5 5.42782
R19713 BIT_SEL[44].n5 BIT_SEL[44] 7.2005
R19714 BIT_SEL[44].t4 BIT_SEL[44] 123.258
R19715 BIT_SEL[44].t1 BIT_SEL[44].n5 117.832
R19716 BIT_SEL[44].t3 BIT_SEL[44].n4 117.832
R19717 BIT_SEL[44].t0 BIT_SEL[44].n3 117.832
R19718 BIT_SEL[44].t2 BIT_SEL[44].n2 117.832
R19719 BIT_SEL[44].t6 BIT_SEL[44].n1 117.832
R19720 BIT_SEL[44].t5 BIT_SEL[44].n0 117.832
R19721 a_14320_38697.t0 a_14320_38697.t1 8.02468
R19722 a_14320_5027.t0 a_14320_5027.t1 8.02156
R19723 a_1340_24783.t0 a_1340_24783.t1 7.42442
R19724 OUT[3] OUT[3].n0 9.0005
R19725 OUT[3].n0 OUT[3].t1 8.56064
R19726 OUT[3].n0 OUT[3].t0 4.38216
R19727 a_20810_5924.t0 a_20810_5924.t1 6.38411
R19728 a_14320_18171.t0 a_14320_18171.t1 6.71945
R19729 a_110_18060.t0 a_110_18060.n0 8.34715
R19730 a_110_18060.n0 a_110_18060.n3 0.1805
R19731 a_110_18060.n3 a_110_18060.n2 4.47779
R19732 a_110_18060.n2 a_110_18060.t3 12.3497
R19733 a_110_18060.n2 a_110_18060.t5 17.192
R19734 a_110_18060.n0 a_110_18060.n1 14.1624
R19735 a_110_18060.n1 a_110_18060.t2 12.3497
R19736 a_110_18060.n1 a_110_18060.t4 17.192
R19737 a_110_18060.n3 a_110_18060.t1 4.44412
R19738 OUT[2] OUT[2].n0 9.0005
R19739 OUT[2].n0 OUT[2].t1 8.56064
R19740 OUT[2].n0 OUT[2].t0 4.38216
R19741 a_7830_39065.t0 a_7830_39065.t1 9.05295
R19742 a_14320_54451.t0 a_14320_54451.t1 8.02468
R19743 BIT_SEL[24].n6 BIT_SEL[24] 8.64211
R19744 BIT_SEL[24] BIT_SEL[24].n6 3.98621
R19745 BIT_SEL[24].n6 BIT_SEL[24].t7 117.008
R19746 BIT_SEL[24] BIT_SEL[24].n0 3.98621
R19747 BIT_SEL[24].n0 BIT_SEL[24] 8.64211
R19748 BIT_SEL[24] BIT_SEL[24].n1 3.98621
R19749 BIT_SEL[24].n1 BIT_SEL[24] 8.64211
R19750 BIT_SEL[24] BIT_SEL[24].n2 3.98621
R19751 BIT_SEL[24].n2 BIT_SEL[24] 8.64211
R19752 BIT_SEL[24] BIT_SEL[24].n3 3.98621
R19753 BIT_SEL[24].n3 BIT_SEL[24] 8.64211
R19754 BIT_SEL[24] BIT_SEL[24].n4 3.98621
R19755 BIT_SEL[24].n4 BIT_SEL[24] 8.64211
R19756 BIT_SEL[24] BIT_SEL[24].n5 3.98621
R19757 BIT_SEL[24].n5 BIT_SEL[24] 8.64211
R19758 BIT_SEL[24].t2 BIT_SEL[24] 120.995
R19759 BIT_SEL[24].t4 BIT_SEL[24].n5 117.008
R19760 BIT_SEL[24].t1 BIT_SEL[24].n4 117.008
R19761 BIT_SEL[24].t0 BIT_SEL[24].n3 117.008
R19762 BIT_SEL[24].t6 BIT_SEL[24].n2 117.008
R19763 BIT_SEL[24].t5 BIT_SEL[24].n1 117.008
R19764 BIT_SEL[24].t3 BIT_SEL[24].n0 117.008
R19765 a_7830_37800.t0 a_7830_37800.t1 5.92569
R19766 a_154_14495.t0 a_154_14495.t1 13.9628
R19767 a_110_14583.t0 a_110_14583.t1 19.5535
R19768 a_1340_40537.t0 a_1340_40537.t1 7.42442
R19769 a_1340_5924.t0 a_1340_5924.t1 6.38411
R19770 a_7830_10294.t0 a_7830_10294.t1 6.71904
R19771 a_20810_14169.t0 a_20810_14169.t1 5.92569
R19772 a_110_60501.t0 a_110_60501.t1 19.5535
R19773 a_154_60413.t0 a_154_60413.t1 13.9628
R19774 BIT_SEL[45].n6 BIT_SEL[45] 5.42621
R19775 BIT_SEL[45] BIT_SEL[45].n6 7.20211
R19776 BIT_SEL[45] BIT_SEL[45].t7 123.463
R19777 BIT_SEL[45].n6 BIT_SEL[45].t6 118.037
R19778 BIT_SEL[45] BIT_SEL[45].n0 7.20211
R19779 BIT_SEL[45].n0 BIT_SEL[45] 5.42621
R19780 BIT_SEL[45] BIT_SEL[45].n1 7.20211
R19781 BIT_SEL[45].n1 BIT_SEL[45] 5.42621
R19782 BIT_SEL[45] BIT_SEL[45].n2 7.20211
R19783 BIT_SEL[45].n2 BIT_SEL[45] 5.42621
R19784 BIT_SEL[45] BIT_SEL[45].n3 7.20211
R19785 BIT_SEL[45].n3 BIT_SEL[45] 5.42621
R19786 BIT_SEL[45] BIT_SEL[45].n4 7.20211
R19787 BIT_SEL[45].n4 BIT_SEL[45] 5.42621
R19788 BIT_SEL[45] BIT_SEL[45].n5 7.20211
R19789 BIT_SEL[45].n5 BIT_SEL[45] 5.42621
R19790 BIT_SEL[45].t3 BIT_SEL[45].n5 118.037
R19791 BIT_SEL[45].t1 BIT_SEL[45].n4 118.037
R19792 BIT_SEL[45].t0 BIT_SEL[45].n3 118.037
R19793 BIT_SEL[45].t5 BIT_SEL[45].n2 118.037
R19794 BIT_SEL[45].t4 BIT_SEL[45].n1 118.037
R19795 BIT_SEL[45].t2 BIT_SEL[45].n0 118.037
R19796 a_14320_40009.t0 a_14320_40009.t1 8.49425
R19797 a_14320_33925.t0 a_14320_33925.t1 6.71945
R19798 BIT_SEL[46].n6 BIT_SEL[46] 6.60907
R19799 BIT_SEL[46] BIT_SEL[46].n6 6.01925
R19800 BIT_SEL[46].n6 BIT_SEL[46].t7 118.243
R19801 BIT_SEL[46] BIT_SEL[46].n0 6.01925
R19802 BIT_SEL[46].n0 BIT_SEL[46] 6.60907
R19803 BIT_SEL[46] BIT_SEL[46].n1 6.01925
R19804 BIT_SEL[46].n1 BIT_SEL[46] 6.60907
R19805 BIT_SEL[46] BIT_SEL[46].n2 6.01925
R19806 BIT_SEL[46].n2 BIT_SEL[46] 6.60907
R19807 BIT_SEL[46] BIT_SEL[46].n3 6.01925
R19808 BIT_SEL[46].n3 BIT_SEL[46] 6.60907
R19809 BIT_SEL[46] BIT_SEL[46].n4 6.01925
R19810 BIT_SEL[46].n4 BIT_SEL[46] 6.60907
R19811 BIT_SEL[46] BIT_SEL[46].n5 6.01925
R19812 BIT_SEL[46].n5 BIT_SEL[46] 6.60907
R19813 BIT_SEL[46].t5 BIT_SEL[46] 124.261
R19814 BIT_SEL[46].t0 BIT_SEL[46].n5 118.243
R19815 BIT_SEL[46].t3 BIT_SEL[46].n4 118.243
R19816 BIT_SEL[46].t1 BIT_SEL[46].n3 118.243
R19817 BIT_SEL[46].t6 BIT_SEL[46].n2 118.243
R19818 BIT_SEL[46].t4 BIT_SEL[46].n1 118.243
R19819 BIT_SEL[46].t2 BIT_SEL[46].n0 118.243
R19820 a_14320_54819.t0 a_14320_54819.t1 9.05295
R19821 a_154_30249.t0 a_154_30249.t1 13.9628
R19822 a_110_30337.t0 a_110_30337.t1 19.5535
R19823 a_110_28321.t0 a_110_28321.t1 19.5535
R19824 a_154_28233.t0 a_154_28233.t1 13.9628
R19825 a_20810_14537.t0 a_20810_14537.t1 6.9546
R19826 a_1340_62696.t0 a_1340_62696.t1 9.05337
R19827 a_1340_33029.t0 a_1340_33029.t1 6.39548
R19828 a_1340_624.t0 a_1340_624.t1 8.49538
R19829 a_110_18956.t2 a_110_18956.n0 2.06607
R19830 a_110_18956.n0 a_110_18956.t1 2.2382
R19831 a_110_18956.n0 a_110_18956.n5 2.6905
R19832 a_110_18956.n5 a_110_18956.t0 4.88081
R19833 a_110_18956.n5 a_110_18956.n1 0.766047
R19834 a_110_18956.n1 a_110_18956.t5 8.68401
R19835 a_110_18956.n3 a_110_18956.n4 5.21793
R19836 a_110_18956.n1 a_110_18956.n3 4.76793
R19837 a_110_18956.n4 a_110_18956.t4 8.51897
R19838 a_110_18956.n4 a_110_18956.t3 4.4523
R19839 a_110_18956.n3 a_110_18956.n2 8.53373
R19840 a_110_18956.n2 a_110_18956.t6 12.3497
R19841 a_110_18956.n2 a_110_18956.t7 17.192
R19842 a_7830_60166.t0 a_7830_60166.t1 8.02156
R19843 BIT_SEL[4].n6 BIT_SEL[4] 10.0837
R19844 BIT_SEL[4] BIT_SEL[4].n6 2.54461
R19845 BIT_SEL[4].n6 BIT_SEL[4].t0 116.186
R19846 BIT_SEL[4] BIT_SEL[4].n0 2.54461
R19847 BIT_SEL[4].n0 BIT_SEL[4] 10.0837
R19848 BIT_SEL[4] BIT_SEL[4].n1 2.54461
R19849 BIT_SEL[4].n1 BIT_SEL[4] 10.0837
R19850 BIT_SEL[4] BIT_SEL[4].n2 2.54461
R19851 BIT_SEL[4].n2 BIT_SEL[4] 10.0837
R19852 BIT_SEL[4] BIT_SEL[4].n3 2.54461
R19853 BIT_SEL[4].n3 BIT_SEL[4] 10.0837
R19854 BIT_SEL[4] BIT_SEL[4].n4 2.54461
R19855 BIT_SEL[4].n4 BIT_SEL[4] 10.0837
R19856 BIT_SEL[4] BIT_SEL[4].n5 2.54461
R19857 BIT_SEL[4].n5 BIT_SEL[4] 10.0837
R19858 BIT_SEL[4].t6 BIT_SEL[4] 118.73
R19859 BIT_SEL[4].t4 BIT_SEL[4].n5 116.186
R19860 BIT_SEL[4].t2 BIT_SEL[4].n4 116.186
R19861 BIT_SEL[4].t3 BIT_SEL[4].n3 116.186
R19862 BIT_SEL[4].t1 BIT_SEL[4].n2 116.186
R19863 BIT_SEL[4].t5 BIT_SEL[4].n1 116.186
R19864 BIT_SEL[4].t7 BIT_SEL[4].n0 116.186
R19865 a_1340_5395.t0 a_1340_5395.t1 7.18327
R19866 a_154_23977.t0 a_154_23977.t1 13.9628
R19867 a_110_24065.t0 a_110_24065.t1 19.5535
R19868 a_110_3202.t2 a_110_3202.n4 4.88081
R19869 a_110_3202.n4 a_110_3202.n5 2.6905
R19870 a_110_3202.n5 a_110_3202.t0 2.06607
R19871 a_110_3202.n5 a_110_3202.t1 2.2382
R19872 a_110_3202.n4 a_110_3202.n0 0.766047
R19873 a_110_3202.n0 a_110_3202.t5 8.68401
R19874 a_110_3202.n2 a_110_3202.n3 5.21793
R19875 a_110_3202.n0 a_110_3202.n2 4.76793
R19876 a_110_3202.n3 a_110_3202.t4 8.51897
R19877 a_110_3202.n3 a_110_3202.t3 4.4523
R19878 a_110_3202.n2 a_110_3202.n1 8.53373
R19879 a_110_3202.n1 a_110_3202.t7 12.3497
R19880 a_110_3202.n1 a_110_3202.t6 17.192
R19881 BIT_SEL[37].t0 BIT_SEL[37] 118.936
R19882 BIT_SEL[37] BIT_SEL[37].n0 10.0837
R19883 BIT_SEL[37] BIT_SEL[37].n0 2.54461
R19884 BIT_SEL[37] BIT_SEL[37].n1 10.0837
R19885 BIT_SEL[37].n1 BIT_SEL[37] 2.54461
R19886 BIT_SEL[37] BIT_SEL[37].n2 10.0837
R19887 BIT_SEL[37].n2 BIT_SEL[37] 2.54461
R19888 BIT_SEL[37] BIT_SEL[37].n3 10.0837
R19889 BIT_SEL[37].n3 BIT_SEL[37] 2.54461
R19890 BIT_SEL[37] BIT_SEL[37].n4 10.0837
R19891 BIT_SEL[37].n4 BIT_SEL[37] 2.54461
R19892 BIT_SEL[37] BIT_SEL[37].n5 10.0837
R19893 BIT_SEL[37].n5 BIT_SEL[37] 2.54461
R19894 BIT_SEL[37] BIT_SEL[37].n6 10.0837
R19895 BIT_SEL[37].n6 BIT_SEL[37] 2.54461
R19896 BIT_SEL[37].t3 BIT_SEL[37].n6 116.391
R19897 BIT_SEL[37].t1 BIT_SEL[37].n5 116.391
R19898 BIT_SEL[37].t6 BIT_SEL[37].n4 116.391
R19899 BIT_SEL[37].t4 BIT_SEL[37].n3 116.391
R19900 BIT_SEL[37].t2 BIT_SEL[37].n2 116.391
R19901 BIT_SEL[37].n1 BIT_SEL[37].t5 116.391
R19902 BIT_SEL[37].n0 BIT_SEL[37].t7 116.391
R19903 a_14320_2417.t0 a_14320_2417.t1 6.71904
R19904 OUT[7] OUT[7].n0 9.0005
R19905 OUT[7].n0 OUT[7].t1 8.56064
R19906 OUT[7].n0 OUT[7].t0 4.38216
R19907 a_14320_21678.t0 a_14320_21678.t1 6.38524
R19908 a_7830_22414.t0 a_7830_22414.t1 6.95418
R19909 a_20810_60166.t0 a_20810_60166.t1 8.02269
R19910 a_1340_22046.t0 a_1340_22046.t1 5.92569
R19911 a_7830_21678.t0 a_7830_21678.t1 6.38411
R19912 a_110_53968.t0 a_110_53968.t1 19.5535
R19913 a_154_53880.t0 a_154_53880.t1 13.9628
R19914 BIT_SEL[6] BIT_SEL[6].n0 3.39479
R19915 BIT_SEL[6] BIT_SEL[6].n0 9.23354
R19916 BIT_SEL[6] BIT_SEL[6].n1 3.39479
R19917 BIT_SEL[6].n1 BIT_SEL[6] 9.23354
R19918 BIT_SEL[6] BIT_SEL[6].n2 3.39479
R19919 BIT_SEL[6].n2 BIT_SEL[6] 9.23354
R19920 BIT_SEL[6] BIT_SEL[6].n3 3.39479
R19921 BIT_SEL[6].n3 BIT_SEL[6] 9.23354
R19922 BIT_SEL[6] BIT_SEL[6].n4 3.39479
R19923 BIT_SEL[6].n4 BIT_SEL[6] 9.23354
R19924 BIT_SEL[6] BIT_SEL[6].n5 3.39479
R19925 BIT_SEL[6].n5 BIT_SEL[6] 9.23354
R19926 BIT_SEL[6] BIT_SEL[6].n6 3.39479
R19927 BIT_SEL[6].n6 BIT_SEL[6] 9.23354
R19928 BIT_SEL[6].t7 BIT_SEL[6] 119.992
R19929 BIT_SEL[6].t6 BIT_SEL[6].n6 116.597
R19930 BIT_SEL[6].t4 BIT_SEL[6].n5 116.597
R19931 BIT_SEL[6].t2 BIT_SEL[6].n4 116.597
R19932 BIT_SEL[6].t1 BIT_SEL[6].n3 116.597
R19933 BIT_SEL[6].t5 BIT_SEL[6].n2 116.597
R19934 BIT_SEL[6].n1 BIT_SEL[6].t3 116.597
R19935 BIT_SEL[6].n0 BIT_SEL[6].t0 116.597
R19936 a_154_46003.t0 a_154_46003.t1 13.9628
R19937 a_110_46091.t0 a_110_46091.t1 19.5535
R19938 a_7830_5027.t0 a_7830_5027.t1 8.02156
R19939 a_20810_55395.t0 a_20810_55395.t1 9.52293
R19940 a_1340_48783.t0 a_1340_48783.t1 6.39548
R19941 a_7830_38168.t0 a_7830_38168.t1 6.95418
R19942 a_20810_56291.t0 a_20810_56291.t1 7.42556
R19943 a_110_47696.t0 a_110_47696.t1 19.5535
R19944 a_154_47608.t0 a_154_47608.t1 13.9628
R19945 a_7830_37432.t0 a_7830_37432.t1 6.38411
R19946 a_7830_20781.t0 a_7830_20781.t1 8.02156
R19947 a_1340_37800.t0 a_1340_37800.t1 5.92611
R19948 a_20810_46045.t0 a_20810_46045.t1 6.9546
R19949 a_7830_9398.t0 a_7830_9398.t1 6.39662
R19950 a_14320_49679.t0 a_14320_49679.t1 6.71904
R19951 a_20810_50048.t0 a_20810_50048.t1 7.5582
R19952 a_20810_34294.t0 a_20810_34294.t1 7.5582
R19953 a_154_46451.t0 a_154_46451.t1 13.9628
R19954 a_110_46539.t0 a_110_46539.t1 19.5535
R19955 a_14320_53186.t0 a_14320_53186.t1 6.38411
R19956 a_7830_9766.t0 a_7830_9766.t1 5.92117
R19957 a_14320_49151.t0 a_14320_49151.t1 5.92117
R19958 a_1340_31188.t0 a_1340_31188.t1 9.05337
R19959 a_1340_16010.t0 a_1340_16010.t1 9.52293
R19960 a_20810_34662.t0 a_20810_34662.t1 6.02155
R19961 a_14320_22943.t0 a_14320_22943.t1 8.02468
R19962 a_154_12479.t0 a_154_12479.t1 13.9628
R19963 a_110_12567.t0 a_110_12567.t1 19.5535
R19964 a_7830_52289.t0 a_7830_52289.t1 8.02156
R19965 a_7830_36903.t0 a_7830_36903.t1 7.18327
R19966 a_1248_19835.t0 a_1248_19835.t1 6.66648
R19967 a_20810_13272.t0 a_20810_13272.t1 7.18213
R19968 BIT_SEL[43].n6 BIT_SEL[43] 4.57764
R19969 BIT_SEL[43] BIT_SEL[43].n6 8.05068
R19970 BIT_SEL[43] BIT_SEL[43].t7 122.203
R19971 BIT_SEL[43].n6 BIT_SEL[43].t2 117.626
R19972 BIT_SEL[43] BIT_SEL[43].n0 8.05068
R19973 BIT_SEL[43].n0 BIT_SEL[43] 4.57764
R19974 BIT_SEL[43] BIT_SEL[43].n1 8.05068
R19975 BIT_SEL[43].n1 BIT_SEL[43] 4.57764
R19976 BIT_SEL[43] BIT_SEL[43].n2 8.05068
R19977 BIT_SEL[43].n2 BIT_SEL[43] 4.57764
R19978 BIT_SEL[43] BIT_SEL[43].n3 8.05068
R19979 BIT_SEL[43].n3 BIT_SEL[43] 4.57764
R19980 BIT_SEL[43] BIT_SEL[43].n4 8.05068
R19981 BIT_SEL[43].n4 BIT_SEL[43] 4.57764
R19982 BIT_SEL[43] BIT_SEL[43].n5 8.05068
R19983 BIT_SEL[43].n5 BIT_SEL[43] 4.57764
R19984 BIT_SEL[43].t5 BIT_SEL[43].n5 117.626
R19985 BIT_SEL[43].t1 BIT_SEL[43].n4 117.626
R19986 BIT_SEL[43].t4 BIT_SEL[43].n3 117.626
R19987 BIT_SEL[43].t6 BIT_SEL[43].n2 117.626
R19988 BIT_SEL[43].t3 BIT_SEL[43].n1 117.626
R19989 BIT_SEL[43].t0 BIT_SEL[43].n0 117.626
R19990 a_14320_16906.t0 a_14320_16906.t1 7.42442
R19991 a_1340_31764.t0 a_1340_31764.t1 9.52293
R19992 a_14320_39065.t0 a_14320_39065.t1 9.05295
R19993 a_20810_16378.t0 a_20810_16378.t1 8.49425
R19994 a_1340_17275.t0 a_1340_17275.t1 6.39548
R19995 a_1248_35589.t0 a_1248_35589.t1 6.66648
R19996 a_7830_8133.t0 a_7830_8133.t1 9.52293
R19997 a_14320_56291.t0 a_14320_56291.t1 7.42442
R19998 BIT_SEL[47].n6 BIT_SEL[47] 6.01764
R19999 BIT_SEL[47] BIT_SEL[47].n6 6.61068
R20000 BIT_SEL[47] BIT_SEL[47].t7 124.466
R20001 BIT_SEL[47].n6 BIT_SEL[47].t6 118.448
R20002 BIT_SEL[47] BIT_SEL[47].n0 6.61068
R20003 BIT_SEL[47].n0 BIT_SEL[47] 6.01764
R20004 BIT_SEL[47] BIT_SEL[47].n1 6.61068
R20005 BIT_SEL[47].n1 BIT_SEL[47] 6.01764
R20006 BIT_SEL[47] BIT_SEL[47].n2 6.61068
R20007 BIT_SEL[47].n2 BIT_SEL[47] 6.01764
R20008 BIT_SEL[47] BIT_SEL[47].n3 6.61068
R20009 BIT_SEL[47].n3 BIT_SEL[47] 6.01764
R20010 BIT_SEL[47] BIT_SEL[47].n4 6.61068
R20011 BIT_SEL[47].n4 BIT_SEL[47] 6.01764
R20012 BIT_SEL[47] BIT_SEL[47].n5 6.61068
R20013 BIT_SEL[47].n5 BIT_SEL[47] 6.01764
R20014 BIT_SEL[47].t3 BIT_SEL[47].n5 118.448
R20015 BIT_SEL[47].t1 BIT_SEL[47].n4 118.448
R20016 BIT_SEL[47].t0 BIT_SEL[47].n3 118.448
R20017 BIT_SEL[47].t5 BIT_SEL[47].n2 118.448
R20018 BIT_SEL[47].t2 BIT_SEL[47].n1 118.448
R20019 BIT_SEL[47].t4 BIT_SEL[47].n0 118.448
R20020 a_14320_39641.t0 a_14320_39641.t1 9.52293
R20021 a_7830_54451.t0 a_7830_54451.t1 8.02468
R20022 a_7830_40906.t0 a_7830_40906.t1 6.39662
R20023 BIT_SEL[26].n6 BIT_SEL[26] 8.05068
R20024 BIT_SEL[26] BIT_SEL[26].n6 4.57764
R20025 BIT_SEL[26].n6 BIT_SEL[26].t7 117.419
R20026 BIT_SEL[26] BIT_SEL[26].n0 4.57764
R20027 BIT_SEL[26].n0 BIT_SEL[26] 8.05068
R20028 BIT_SEL[26] BIT_SEL[26].n1 4.57764
R20029 BIT_SEL[26].n1 BIT_SEL[26] 8.05068
R20030 BIT_SEL[26] BIT_SEL[26].n2 4.57764
R20031 BIT_SEL[26].n2 BIT_SEL[26] 8.05068
R20032 BIT_SEL[26] BIT_SEL[26].n3 4.57764
R20033 BIT_SEL[26].n3 BIT_SEL[26] 8.05068
R20034 BIT_SEL[26] BIT_SEL[26].n4 4.57764
R20035 BIT_SEL[26].n4 BIT_SEL[26] 8.05068
R20036 BIT_SEL[26] BIT_SEL[26].n5 4.57764
R20037 BIT_SEL[26].n5 BIT_SEL[26] 8.05068
R20038 BIT_SEL[26].t5 BIT_SEL[26] 121.998
R20039 BIT_SEL[26].t4 BIT_SEL[26].n5 117.419
R20040 BIT_SEL[26].t2 BIT_SEL[26].n4 117.419
R20041 BIT_SEL[26].t0 BIT_SEL[26].n3 117.419
R20042 BIT_SEL[26].t6 BIT_SEL[26].n2 117.419
R20043 BIT_SEL[26].t3 BIT_SEL[26].n1 117.419
R20044 BIT_SEL[26].t1 BIT_SEL[26].n0 117.419
R20045 a_20810_32132.t0 a_20810_32132.t1 8.49538
R20046 a_1340_17643.t0 a_1340_17643.t1 5.92075
R20047 a_7830_26417.t0 a_7830_26417.t1 7.5582
R20048 a_154_60861.t0 a_154_60861.t1 13.9628
R20049 a_110_60949.t0 a_110_60949.t1 19.5535
R20050 a_14320_50048.t0 a_14320_50048.t1 7.55862
R20051 a_154_43987.t0 a_154_43987.t1 13.9628
R20052 a_110_44075.t0 a_110_44075.t1 19.5535
R20053 a_14320_48414.t0 a_14320_48414.t1 7.42442
R20054 a_7830_23887.t0 a_7830_23887.t1 9.52407
R20055 a_7830_26785.t0 a_7830_26785.t1 6.02155
R20056 a_20718_51343.t0 a_20718_51343.t1 6.66648
R20057 a_20810_38697.t0 a_20810_38697.t1 8.02468
R20058 a_14320_22046.t0 a_14320_22046.t1 5.92611
R20059 BIT_SEL[29].n6 BIT_SEL[29] 5.42621
R20060 BIT_SEL[29] BIT_SEL[29].n6 7.20211
R20061 BIT_SEL[29] BIT_SEL[29].t7 123.463
R20062 BIT_SEL[29].n6 BIT_SEL[29].t0 118.037
R20063 BIT_SEL[29] BIT_SEL[29].n0 7.20211
R20064 BIT_SEL[29].n0 BIT_SEL[29] 5.42621
R20065 BIT_SEL[29] BIT_SEL[29].n1 7.20211
R20066 BIT_SEL[29].n1 BIT_SEL[29] 5.42621
R20067 BIT_SEL[29] BIT_SEL[29].n2 7.20211
R20068 BIT_SEL[29].n2 BIT_SEL[29] 5.42621
R20069 BIT_SEL[29] BIT_SEL[29].n3 7.20211
R20070 BIT_SEL[29].n3 BIT_SEL[29] 5.42621
R20071 BIT_SEL[29] BIT_SEL[29].n4 7.20211
R20072 BIT_SEL[29].n4 BIT_SEL[29] 5.42621
R20073 BIT_SEL[29] BIT_SEL[29].n5 7.20211
R20074 BIT_SEL[29].n5 BIT_SEL[29] 5.42621
R20075 BIT_SEL[29].t4 BIT_SEL[29].n5 118.037
R20076 BIT_SEL[29].t2 BIT_SEL[29].n4 118.037
R20077 BIT_SEL[29].t1 BIT_SEL[29].n3 118.037
R20078 BIT_SEL[29].t6 BIT_SEL[29].n2 118.037
R20079 BIT_SEL[29].t5 BIT_SEL[29].n1 118.037
R20080 BIT_SEL[29].t3 BIT_SEL[29].n0 118.037
R20081 a_7830_8501.t0 a_7830_8501.t1 8.49425
R20082 a_7738_19835.t0 a_7738_19835.t1 6.66648
R20083 a_7830_39641.t0 a_7830_39641.t1 9.52407
R20084 a_14320_28658.t0 a_14320_28658.t1 8.02156
R20085 a_7830_5395.t0 a_7830_5395.t1 7.18327
R20086 a_7830_42539.t0 a_7830_42539.t1 6.02155
R20087 a_20810_18908.t0 a_20810_18908.t1 6.02155
R20088 a_20810_18171.t0 a_20810_18171.t1 6.71945
R20089 a_1340_49151.t0 a_1340_49151.t1 5.92075
R20090 a_14320_22414.t0 a_14320_22414.t1 6.9546
R20091 a_20810_54451.t0 a_20810_54451.t1 8.02468
R20092 a_7830_21149.t0 a_7830_21149.t1 7.18327
R20093 a_14320_9029.t0 a_14320_9029.t1 7.42442
R20094 a_14320_44412.t0 a_14320_44412.t1 8.02156
R20095 a_7830_57556.t0 a_7830_57556.t1 6.71904
R20096 a_20810_33925.t0 a_20810_33925.t1 6.71945
R20097 a_1340_2786.t0 a_1340_2786.t1 7.55862
R20098 a_154_4602.t0 a_154_4602.t1 13.9628
R20099 a_110_4690.t0 a_110_4690.t1 19.5535
R20100 a_14320_10663.t0 a_14320_10663.t1 7.55862
R20101 a_154_13599.t0 a_154_13599.t1 13.9628
R20102 a_110_13687.t0 a_110_13687.t1 19.5535
R20103 a_7830_58293.t0 a_7830_58293.t1 6.02155
R20104 a_1340_52289.t0 a_1340_52289.t1 8.02156
R20105 BIT_SEL[61].n6 BIT_SEL[61] 5.42621
R20106 BIT_SEL[61] BIT_SEL[61].n6 7.20211
R20107 BIT_SEL[61] BIT_SEL[61].t6 123.463
R20108 BIT_SEL[61].n6 BIT_SEL[61].t1 118.037
R20109 BIT_SEL[61] BIT_SEL[61].n0 7.20211
R20110 BIT_SEL[61].n0 BIT_SEL[61] 5.42621
R20111 BIT_SEL[61] BIT_SEL[61].n1 7.20211
R20112 BIT_SEL[61].n1 BIT_SEL[61] 5.42621
R20113 BIT_SEL[61] BIT_SEL[61].n2 7.20211
R20114 BIT_SEL[61].n2 BIT_SEL[61] 5.42621
R20115 BIT_SEL[61] BIT_SEL[61].n3 7.20211
R20116 BIT_SEL[61].n3 BIT_SEL[61] 5.42621
R20117 BIT_SEL[61] BIT_SEL[61].n4 7.20211
R20118 BIT_SEL[61].n4 BIT_SEL[61] 5.42621
R20119 BIT_SEL[61] BIT_SEL[61].n5 7.20211
R20120 BIT_SEL[61].n5 BIT_SEL[61] 5.42621
R20121 BIT_SEL[61].t4 BIT_SEL[61].n5 118.037
R20122 BIT_SEL[61].t2 BIT_SEL[61].n4 118.037
R20123 BIT_SEL[61].t0 BIT_SEL[61].n3 118.037
R20124 BIT_SEL[61].t7 BIT_SEL[61].n2 118.037
R20125 BIT_SEL[61].t5 BIT_SEL[61].n1 118.037
R20126 BIT_SEL[61].t3 BIT_SEL[61].n0 118.037
R20127 a_20810_40009.t0 a_20810_40009.t1 8.49425
R20128 a_110_7602.t0 a_110_7602.t1 19.5535
R20129 a_154_7514.t0 a_154_7514.t1 13.9628
R20130 a_20810_54819.t0 a_20810_54819.t1 9.05337
R20131 a_14320_11031.t0 a_14320_11031.t1 6.02155
R20132 a_110_50464.n0 a_110_50464.t0 2.06607
R20133 a_110_50464.t2 a_110_50464.n0 2.2382
R20134 a_110_50464.n0 a_110_50464.n5 2.6905
R20135 a_110_50464.n5 a_110_50464.t1 4.88081
R20136 a_110_50464.n5 a_110_50464.n1 0.766047
R20137 a_110_50464.n1 a_110_50464.t5 8.68401
R20138 a_110_50464.n3 a_110_50464.n4 5.21793
R20139 a_110_50464.n1 a_110_50464.n3 4.76793
R20140 a_110_50464.n4 a_110_50464.t4 8.51897
R20141 a_110_50464.n4 a_110_50464.t3 4.4523
R20142 a_110_50464.n3 a_110_50464.n2 8.53373
R20143 a_110_50464.n2 a_110_50464.t6 12.3497
R20144 a_110_50464.n2 a_110_50464.t7 17.192
R20145 a_20810_21678.t0 a_20810_21678.t1 6.38411
R20146 a_7830_1521.t0 a_7830_1521.t1 6.39662
R20147 a_14320_47518.t0 a_14320_47518.t1 9.52407
R20148 a_14320_7557.t0 a_14320_7557.t1 9.05295
R20149 a_14320_53922.t0 a_14320_53922.t1 6.95418
R20150 a_1340_33397.t0 a_1340_33397.t1 5.92075
R20151 a_7830_41274.t0 a_7830_41274.t1 5.92117
R20152 a_1340_32132.t0 a_1340_32132.t1 8.49425
R20153 a_154_45107.t0 a_154_45107.t1 13.9628
R20154 a_110_45195.t0 a_110_45195.t1 19.5535
R20155 a_14320_42171.t0 a_14320_42171.t1 7.5582
R20156 a_1340_61063.t0 a_1340_61063.t1 6.38524
R20157 a_14320_1889.t0 a_14320_1889.t1 5.92075
R20158 a_154_7066.t0 a_154_7066.t1 13.9628
R20159 a_110_7154.t0 a_110_7154.t1 19.5535
R20160 a_14320_8501.t0 a_14320_8501.t1 8.49425
R20161 BIT_SEL[53].t4 BIT_SEL[53] 118.936
R20162 BIT_SEL[53] BIT_SEL[53].n0 10.0837
R20163 BIT_SEL[53] BIT_SEL[53].n0 2.54461
R20164 BIT_SEL[53] BIT_SEL[53].n1 10.0837
R20165 BIT_SEL[53].n1 BIT_SEL[53] 2.54461
R20166 BIT_SEL[53] BIT_SEL[53].n2 10.0837
R20167 BIT_SEL[53].n2 BIT_SEL[53] 2.54461
R20168 BIT_SEL[53] BIT_SEL[53].n3 10.0837
R20169 BIT_SEL[53].n3 BIT_SEL[53] 2.54461
R20170 BIT_SEL[53] BIT_SEL[53].n4 10.0837
R20171 BIT_SEL[53].n4 BIT_SEL[53] 2.54461
R20172 BIT_SEL[53] BIT_SEL[53].n5 10.0837
R20173 BIT_SEL[53].n5 BIT_SEL[53] 2.54461
R20174 BIT_SEL[53] BIT_SEL[53].n6 10.0837
R20175 BIT_SEL[53].n6 BIT_SEL[53] 2.54461
R20176 BIT_SEL[53].t2 BIT_SEL[53].n6 116.391
R20177 BIT_SEL[53].t0 BIT_SEL[53].n5 116.391
R20178 BIT_SEL[53].t6 BIT_SEL[53].n4 116.391
R20179 BIT_SEL[53].t3 BIT_SEL[53].n3 116.391
R20180 BIT_SEL[53].t1 BIT_SEL[53].n2 116.391
R20181 BIT_SEL[53].n1 BIT_SEL[53].t5 116.391
R20182 BIT_SEL[53].n0 BIT_SEL[53].t7 116.391
R20183 a_20810_49679.t0 a_20810_49679.t1 6.71904
R20184 a_154_29801.t0 a_154_29801.t1 13.9628
R20185 a_110_29889.t0 a_110_29889.t1 19.5535
R20186 a_14320_18908.t0 a_14320_18908.t1 6.02155
R20187 a_20810_53186.t0 a_20810_53186.t1 6.38411
R20188 a_154_31854.t0 a_154_31854.t1 13.9628
R20189 a_110_31942.t0 a_110_31942.t1 19.5535
R20190 a_20810_49151.t0 a_20810_49151.t1 5.92075
R20191 a_154_794.t0 a_154_794.t1 13.9628
R20192 a_110_882.t0 a_110_882.t1 19.5535
R20193 a_14320_24255.t0 a_14320_24255.t1 8.49425
R20194 BIT_SEL[27].n6 BIT_SEL[27] 4.57764
R20195 BIT_SEL[27] BIT_SEL[27].n6 8.05068
R20196 BIT_SEL[27] BIT_SEL[27].t0 122.203
R20197 BIT_SEL[27].n6 BIT_SEL[27].t3 117.626
R20198 BIT_SEL[27] BIT_SEL[27].n0 8.05068
R20199 BIT_SEL[27].n0 BIT_SEL[27] 4.57764
R20200 BIT_SEL[27] BIT_SEL[27].n1 8.05068
R20201 BIT_SEL[27].n1 BIT_SEL[27] 4.57764
R20202 BIT_SEL[27] BIT_SEL[27].n2 8.05068
R20203 BIT_SEL[27].n2 BIT_SEL[27] 4.57764
R20204 BIT_SEL[27] BIT_SEL[27].n3 8.05068
R20205 BIT_SEL[27].n3 BIT_SEL[27] 4.57764
R20206 BIT_SEL[27] BIT_SEL[27].n4 8.05068
R20207 BIT_SEL[27].n4 BIT_SEL[27] 4.57764
R20208 BIT_SEL[27] BIT_SEL[27].n5 8.05068
R20209 BIT_SEL[27].n5 BIT_SEL[27] 4.57764
R20210 BIT_SEL[27].t6 BIT_SEL[27].n5 117.626
R20211 BIT_SEL[27].t2 BIT_SEL[27].n4 117.626
R20212 BIT_SEL[27].t5 BIT_SEL[27].n3 117.626
R20213 BIT_SEL[27].t7 BIT_SEL[27].n2 117.626
R20214 BIT_SEL[27].t4 BIT_SEL[27].n1 117.626
R20215 BIT_SEL[27].t1 BIT_SEL[27].n0 117.626
R20216 a_7830_1152.t0 a_7830_1152.t1 7.42442
R20217 a_20810_53554.t0 a_20810_53554.t1 5.92569
R20218 a_7830_13801.t0 a_7830_13801.t1 6.38411
R20219 a_20810_22943.t0 a_20810_22943.t1 8.02468
R20220 BIT_SEL[59].n6 BIT_SEL[59] 4.57764
R20221 BIT_SEL[59] BIT_SEL[59].n6 8.05068
R20222 BIT_SEL[59] BIT_SEL[59].t2 122.203
R20223 BIT_SEL[59].n6 BIT_SEL[59].t7 117.626
R20224 BIT_SEL[59] BIT_SEL[59].n0 8.05068
R20225 BIT_SEL[59].n0 BIT_SEL[59] 4.57764
R20226 BIT_SEL[59] BIT_SEL[59].n1 8.05068
R20227 BIT_SEL[59].n1 BIT_SEL[59] 4.57764
R20228 BIT_SEL[59] BIT_SEL[59].n2 8.05068
R20229 BIT_SEL[59].n2 BIT_SEL[59] 4.57764
R20230 BIT_SEL[59] BIT_SEL[59].n3 8.05068
R20231 BIT_SEL[59].n3 BIT_SEL[59] 4.57764
R20232 BIT_SEL[59] BIT_SEL[59].n4 8.05068
R20233 BIT_SEL[59].n4 BIT_SEL[59] 4.57764
R20234 BIT_SEL[59] BIT_SEL[59].n5 8.05068
R20235 BIT_SEL[59].n5 BIT_SEL[59] 4.57764
R20236 BIT_SEL[59].t5 BIT_SEL[59].n5 117.626
R20237 BIT_SEL[59].t1 BIT_SEL[59].n4 117.626
R20238 BIT_SEL[59].t4 BIT_SEL[59].n3 117.626
R20239 BIT_SEL[59].t6 BIT_SEL[59].n2 117.626
R20240 BIT_SEL[59].t3 BIT_SEL[59].n1 117.626
R20241 BIT_SEL[59].t0 BIT_SEL[59].n0 117.626
R20242 a_20810_16906.t0 a_20810_16906.t1 7.42442
R20243 a_20810_39065.t0 a_20810_39065.t1 9.05337
R20244 a_7830_15434.t0 a_7830_15434.t1 9.05337
R20245 a_1340_47886.t0 a_1340_47886.t1 8.49538
R20246 a_7830_48414.t0 a_7830_48414.t1 7.42442
R20247 a_14320_30820.t0 a_14320_30820.t1 8.02468
R20248 a_20810_39641.t0 a_20810_39641.t1 9.52293
R20249 a_14320_10294.t0 a_14320_10294.t1 6.71945
R20250 a_1340_57925.t0 a_1340_57925.t1 7.55862
R20251 a_1340_2417.t0 a_1340_2417.t1 6.71904
R20252 a_1340_36535.t0 a_1340_36535.t1 8.02269
R20253 a_7830_31188.t0 a_7830_31188.t1 9.05337
R20254 a_1248_51343.t0 a_1248_51343.t1 6.66648
R20255 a_14320_46574.t0 a_14320_46574.t1 8.02427
R20256 a_14320_61799.t0 a_14320_61799.t1 6.95418
R20257 a_7830_45309.t0 a_7830_45309.t1 6.38524
R20258 a_20810_48414.t0 a_20810_48414.t1 7.42442
R20259 a_7830_46942.t0 a_7830_46942.t1 9.05337
R20260 a_14320_26048.t0 a_14320_26048.t1 6.71945
R20261 a_20810_9766.t0 a_20810_9766.t1 5.92075
R20262 a_20810_22046.t0 a_20810_22046.t1 5.92569
R20263 a_154_22372.t0 a_154_22372.t1 13.9628
R20264 a_110_22460.t0 a_110_22460.t1 19.5535
R20265 BIT_SEL[41].n6 BIT_SEL[41] 3.98461
R20266 BIT_SEL[41] BIT_SEL[41].n6 8.64371
R20267 BIT_SEL[41] BIT_SEL[41].t0 121.198
R20268 BIT_SEL[41].n6 BIT_SEL[41].t6 117.215
R20269 BIT_SEL[41] BIT_SEL[41].n0 8.64371
R20270 BIT_SEL[41].n0 BIT_SEL[41] 3.98461
R20271 BIT_SEL[41] BIT_SEL[41].n1 8.64371
R20272 BIT_SEL[41].n1 BIT_SEL[41] 3.98461
R20273 BIT_SEL[41] BIT_SEL[41].n2 8.64371
R20274 BIT_SEL[41].n2 BIT_SEL[41] 3.98461
R20275 BIT_SEL[41] BIT_SEL[41].n3 8.64371
R20276 BIT_SEL[41].n3 BIT_SEL[41] 3.98461
R20277 BIT_SEL[41] BIT_SEL[41].n4 8.64371
R20278 BIT_SEL[41].n4 BIT_SEL[41] 3.98461
R20279 BIT_SEL[41] BIT_SEL[41].n5 8.64371
R20280 BIT_SEL[41].n5 BIT_SEL[41] 3.98461
R20281 BIT_SEL[41].t4 BIT_SEL[41].n5 117.215
R20282 BIT_SEL[41].t2 BIT_SEL[41].n4 117.215
R20283 BIT_SEL[41].t7 BIT_SEL[41].n3 117.215
R20284 BIT_SEL[41].t1 BIT_SEL[41].n2 117.215
R20285 BIT_SEL[41].t5 BIT_SEL[41].n1 117.215
R20286 BIT_SEL[41].t3 BIT_SEL[41].n0 117.215
R20287 a_7830_14537.t0 a_7830_14537.t1 6.95418
R20288 a_14320_47886.t0 a_14320_47886.t1 8.49425
R20289 a_14320_41802.t0 a_14320_41802.t1 6.71945
R20290 a_1340_14169.t0 a_1340_14169.t1 5.92611
R20291 a_7830_60534.t0 a_7830_60534.t1 7.18327
R20292 a_1340_49679.t0 a_1340_49679.t1 6.71945
R20293 a_20810_37800.t0 a_20810_37800.t1 5.92569
R20294 a_7830_61431.t0 a_7830_61431.t1 5.92611
R20295 a_20810_22414.t0 a_20810_22414.t1 6.9546
R20296 a_7830_256.t0 a_7830_256.t1 9.52407
R20297 a_1340_22414.t0 a_1340_22414.t1 6.9546
R20298 a_20810_10663.t0 a_20810_10663.t1 7.55862
R20299 a_154_51864.t0 a_154_51864.t1 13.9628
R20300 a_110_51952.t0 a_110_51952.t1 19.5535
R20301 a_7830_30291.t0 a_7830_30291.t1 6.95418
R20302 a_154_22820.t0 a_154_22820.t1 13.9628
R20303 a_110_22908.t0 a_110_22908.t1 19.5535
R20304 a_7830_12904.t0 a_7830_12904.t1 8.02156
R20305 a_1340_29923.t0 a_1340_29923.t1 5.92611
R20306 a_110_6706.t0 a_110_6706.t1 19.5535
R20307 a_154_6618.t0 a_154_6618.t1 13.9628
R20308 a_1340_38168.t0 a_1340_38168.t1 6.9546
R20309 a_20810_11031.t0 a_20810_11031.t1 6.02155
R20310 a_14320_15066.t0 a_14320_15066.t1 8.02427
R20311 a_154_16548.t0 a_154_16548.t1 13.9628
R20312 a_110_16636.t0 a_110_16636.t1 19.5535
R20313 a_1340_56660.t0 a_1340_56660.t1 6.39548
R20314 a_14320_30291.t0 a_14320_30291.t1 6.9546
R20315 a_7830_46045.t0 a_7830_46045.t1 6.9546
R20316 a_1340_45677.t0 a_1340_45677.t1 5.92569
R20317 a_154_38574.t0 a_154_38574.t1 13.9628
R20318 a_110_38662.t0 a_110_38662.t1 19.5535
R20319 a_14320_256.t0 a_14320_256.t1 9.52407
R20320 a_20810_53922.t0 a_20810_53922.t1 6.9546
R20321 a_14320_15434.t0 a_14320_15434.t1 9.05295
R20322 a_14320_57556.t0 a_14320_57556.t1 6.71904
R20323 a_14320_21149.t0 a_14320_21149.t1 7.18327
R20324 a_20810_42171.t0 a_20810_42171.t1 7.5582
R20325 a_20810_8501.t0 a_20810_8501.t1 8.49538
R20326 a_1248_11958.t0 a_1248_11958.t1 6.66648
R20327 a_14320_61063.t0 a_14320_61063.t1 6.38524
R20328 a_154_54328.t0 a_154_54328.t1 13.9628
R20329 a_110_54416.t0 a_110_54416.t1 19.5535
R20330 a_20810_5395.t0 a_20810_5395.t1 7.18213
R20331 BIT_SEL[1].t0 BIT_SEL[1] 116.918
R20332 BIT_SEL[1] BIT_SEL[1].n0 11.2682
R20333 BIT_SEL[1] BIT_SEL[1].n0 1.36014
R20334 BIT_SEL[1] BIT_SEL[1].n1 11.2682
R20335 BIT_SEL[1].n1 BIT_SEL[1] 1.36014
R20336 BIT_SEL[1] BIT_SEL[1].n2 11.2682
R20337 BIT_SEL[1].n2 BIT_SEL[1] 1.36014
R20338 BIT_SEL[1] BIT_SEL[1].n3 11.2682
R20339 BIT_SEL[1].n3 BIT_SEL[1] 1.36014
R20340 BIT_SEL[1] BIT_SEL[1].n4 11.2682
R20341 BIT_SEL[1].n4 BIT_SEL[1] 1.36014
R20342 BIT_SEL[1] BIT_SEL[1].n5 11.2682
R20343 BIT_SEL[1].n5 BIT_SEL[1] 1.36014
R20344 BIT_SEL[1] BIT_SEL[1].n6 11.2682
R20345 BIT_SEL[1].n6 BIT_SEL[1] 1.36014
R20346 BIT_SEL[1].t4 BIT_SEL[1].n6 115.558
R20347 BIT_SEL[1].t7 BIT_SEL[1].n5 115.558
R20348 BIT_SEL[1].t3 BIT_SEL[1].n4 115.558
R20349 BIT_SEL[1].t5 BIT_SEL[1].n3 115.558
R20350 BIT_SEL[1].t2 BIT_SEL[1].n2 115.558
R20351 BIT_SEL[1].n1 BIT_SEL[1].t1 115.558
R20352 BIT_SEL[1].n0 BIT_SEL[1].t6 115.558
R20353 a_1340_3154.t0 a_1340_3154.t1 6.02155
R20354 a_154_48056.t0 a_154_48056.t1 13.9628
R20355 a_110_48144.t0 a_110_48144.t1 19.5535
R20356 a_14320_36903.t0 a_14320_36903.t1 7.18213
R20357 a_7830_36535.t0 a_7830_36535.t1 8.02156
R20358 a_154_20356.t0 a_154_20356.t1 13.9628
R20359 a_110_20444.t0 a_110_20444.t1 19.5535
R20360 COL_PROG_N[1] COL_PROG_N[1].n0 0.0965
R20361 COL_PROG_N[1].n0 COL_PROG_N[1].n1 0.3065
R20362 COL_PROG_N[1].n1 COL_PROG_N[1].n2 0.3065
R20363 COL_PROG_N[1].n2 COL_PROG_N[1].t1 292.788
R20364 COL_PROG_N[1].n2 COL_PROG_N[1].t3 292.481
R20365 COL_PROG_N[1].n1 COL_PROG_N[1].t0 292.481
R20366 COL_PROG_N[1].n0 COL_PROG_N[1].t2 292.481
R20367 a_20810_16010.t0 a_20810_16010.t1 9.52407
R20368 a_14320_24783.t0 a_14320_24783.t1 7.42442
R20369 a_14320_46942.t0 a_14320_46942.t1 9.05295
R20370 a_20810_24255.t0 a_20810_24255.t1 8.49538
R20371 a_14320_6660.t0 a_14320_6660.t1 6.95418
R20372 a_1248_43466.t0 a_1248_43466.t1 6.66648
R20373 a_14320_40537.t0 a_14320_40537.t1 7.42442
R20374 a_20810_32660.t0 a_20810_32660.t1 7.42442
R20375 a_20810_31764.t0 a_20810_31764.t1 9.52407
R20376 a_1340_8133.t0 a_1340_8133.t1 9.52293
R20377 a_1340_54451.t0 a_1340_54451.t1 8.02427
R20378 a_14320_50416.t0 a_14320_50416.t1 6.02155
R20379 a_1340_25520.t0 a_1340_25520.t1 5.92075
R20380 a_7830_2786.t0 a_7830_2786.t1 7.5582
R20381 a_7830_50048.t0 a_7830_50048.t1 7.5582
R20382 a_20810_30820.t0 a_20810_30820.t1 8.02468
R20383 a_7830_34294.t0 a_7830_34294.t1 7.5582
R20384 a_7738_4081.t0 a_7738_4081.t1 6.66648
R20385 a_20810_10294.t0 a_20810_10294.t1 6.71904
R20386 a_7830_34662.t0 a_7830_34662.t1 6.02155
R20387 COL_PROG_N[3] COL_PROG_N[3].n0 0.0965
R20388 COL_PROG_N[3].n0 COL_PROG_N[3].n1 0.3065
R20389 COL_PROG_N[3].n1 COL_PROG_N[3].n2 0.3065
R20390 COL_PROG_N[3].n2 COL_PROG_N[3].t2 292.788
R20391 COL_PROG_N[3].n2 COL_PROG_N[3].t0 292.481
R20392 COL_PROG_N[3].n1 COL_PROG_N[3].t3 292.481
R20393 COL_PROG_N[3].n0 COL_PROG_N[3].t1 292.481
R20394 a_1340_7189.t0 a_1340_7189.t1 8.02468
R20395 a_20810_46574.t0 a_20810_46574.t1 8.02468
R20396 a_1340_39641.t0 a_1340_39641.t1 9.52407
R20397 a_14320_29923.t0 a_14320_29923.t1 5.92611
R20398 a_7830_13272.t0 a_7830_13272.t1 7.18327
R20399 a_20810_61799.t0 a_20810_61799.t1 6.9546
R20400 a_20810_26048.t0 a_20810_26048.t1 6.71904
R20401 a_14320_5924.t0 a_14320_5924.t1 6.38524
R20402 a_20810_47518.t0 a_20810_47518.t1 9.52293
R20403 COL_PROG_N[5] COL_PROG_N[5].n0 0.0965
R20404 COL_PROG_N[5].n0 COL_PROG_N[5].n1 0.3065
R20405 COL_PROG_N[5].n1 COL_PROG_N[5].n2 0.3065
R20406 COL_PROG_N[5].n2 COL_PROG_N[5].t2 292.788
R20407 COL_PROG_N[5].n2 COL_PROG_N[5].t0 292.481
R20408 COL_PROG_N[5].n1 COL_PROG_N[5].t3 292.481
R20409 COL_PROG_N[5].n0 COL_PROG_N[5].t1 292.481
R20410 a_1340_9766.t0 a_1340_9766.t1 5.92075
R20411 a_7830_6292.t0 a_7830_6292.t1 5.92569
R20412 a_20810_1152.t0 a_20810_1152.t1 7.42442
R20413 a_154_21476.t0 a_154_21476.t1 13.9628
R20414 a_110_21564.t0 a_110_21564.t1 19.5535
R20415 a_14320_624.t0 a_14320_624.t1 8.49538
R20416 a_14320_5395.t0 a_14320_5395.t1 7.18327
R20417 a_20810_47886.t0 a_20810_47886.t1 8.49425
R20418 a_20810_41802.t0 a_20810_41802.t1 6.71945
R20419 a_14320_32660.t0 a_14320_32660.t1 7.42556
R20420 COL_PROG_N[7] COL_PROG_N[7].n0 0.0965
R20421 COL_PROG_N[7].n0 COL_PROG_N[7].n1 0.3065
R20422 COL_PROG_N[7].n1 COL_PROG_N[7].n2 0.3065
R20423 COL_PROG_N[7].n2 COL_PROG_N[7].t2 292.788
R20424 COL_PROG_N[7].n2 COL_PROG_N[7].t0 292.481
R20425 COL_PROG_N[7].n1 COL_PROG_N[7].t3 292.481
R20426 COL_PROG_N[7].n0 COL_PROG_N[7].t1 292.481
R20427 a_110_5362.t0 a_110_5362.t1 19.5535
R20428 a_154_5274.t0 a_154_5274.t1 13.9628
R20429 a_1340_29555.t0 a_1340_29555.t1 6.38524
R20430 a_7830_55763.t0 a_7830_55763.t1 8.49425
R20431 a_7738_51343.t0 a_7738_51343.t1 6.66648
R20432 a_1340_41274.t0 a_1340_41274.t1 5.92075
R20433 a_7830_56660.t0 a_7830_56660.t1 6.39662
R20434 BIT_SEL[28].n6 BIT_SEL[28] 7.2005
R20435 BIT_SEL[28] BIT_SEL[28].n6 5.42782
R20436 BIT_SEL[28].n6 BIT_SEL[28].t7 117.832
R20437 BIT_SEL[28] BIT_SEL[28].n0 5.42782
R20438 BIT_SEL[28].n0 BIT_SEL[28] 7.2005
R20439 BIT_SEL[28] BIT_SEL[28].n1 5.42782
R20440 BIT_SEL[28].n1 BIT_SEL[28] 7.2005
R20441 BIT_SEL[28] BIT_SEL[28].n2 5.42782
R20442 BIT_SEL[28].n2 BIT_SEL[28] 7.2005
R20443 BIT_SEL[28] BIT_SEL[28].n3 5.42782
R20444 BIT_SEL[28].n3 BIT_SEL[28] 7.2005
R20445 BIT_SEL[28] BIT_SEL[28].n4 5.42782
R20446 BIT_SEL[28].n4 BIT_SEL[28] 7.2005
R20447 BIT_SEL[28] BIT_SEL[28].n5 5.42782
R20448 BIT_SEL[28].n5 BIT_SEL[28] 7.2005
R20449 BIT_SEL[28].t4 BIT_SEL[28] 123.258
R20450 BIT_SEL[28].t1 BIT_SEL[28].n5 117.832
R20451 BIT_SEL[28].t3 BIT_SEL[28].n4 117.832
R20452 BIT_SEL[28].t0 BIT_SEL[28].n3 117.832
R20453 BIT_SEL[28].t2 BIT_SEL[28].n2 117.832
R20454 BIT_SEL[28].t6 BIT_SEL[28].n1 117.832
R20455 BIT_SEL[28].t5 BIT_SEL[28].n0 117.832
R20456 a_7830_38697.t0 a_7830_38697.t1 8.02468
R20457 a_20810_6660.t0 a_20810_6660.t1 6.95418
R20458 a_20810_15066.t0 a_20810_15066.t1 8.02468
R20459 a_20810_30291.t0 a_20810_30291.t1 6.9546
R20460 a_154_52984.t0 a_154_52984.t1 13.9628
R20461 a_110_53072.t0 a_110_53072.t1 19.5535
R20462 a_7830_18171.t0 a_7830_18171.t1 6.71904
R20463 a_14228_59220.t0 a_14228_59220.t1 6.66648
R20464 a_1340_39065.t0 a_1340_39065.t1 9.05337
R20465 a_20810_15434.t0 a_20810_15434.t1 9.05337
R20466 a_14320_26785.t0 a_14320_26785.t1 6.02155
R20467 a_1340_18908.t0 a_1340_18908.t1 6.02155
R20468 a_154_37678.t0 a_154_37678.t1 13.9628
R20469 a_110_37766.t0 a_110_37766.t1 19.5535
R20470 BIT_SEL[8] BIT_SEL[8].n0 3.98621
R20471 BIT_SEL[8] BIT_SEL[8].n0 8.64211
R20472 BIT_SEL[8] BIT_SEL[8].n1 3.98621
R20473 BIT_SEL[8].n1 BIT_SEL[8] 8.64211
R20474 BIT_SEL[8] BIT_SEL[8].n2 3.98621
R20475 BIT_SEL[8].n2 BIT_SEL[8] 8.64211
R20476 BIT_SEL[8] BIT_SEL[8].n3 3.98621
R20477 BIT_SEL[8].n3 BIT_SEL[8] 8.64211
R20478 BIT_SEL[8] BIT_SEL[8].n4 3.98621
R20479 BIT_SEL[8].n4 BIT_SEL[8] 8.64211
R20480 BIT_SEL[8] BIT_SEL[8].n5 3.98621
R20481 BIT_SEL[8].n5 BIT_SEL[8] 8.64211
R20482 BIT_SEL[8] BIT_SEL[8].n6 3.98621
R20483 BIT_SEL[8].n6 BIT_SEL[8] 8.64211
R20484 BIT_SEL[8].t3 BIT_SEL[8] 120.995
R20485 BIT_SEL[8].t5 BIT_SEL[8].n6 117.008
R20486 BIT_SEL[8].t2 BIT_SEL[8].n5 117.008
R20487 BIT_SEL[8].t1 BIT_SEL[8].n4 117.008
R20488 BIT_SEL[8].t7 BIT_SEL[8].n3 117.008
R20489 BIT_SEL[8].t6 BIT_SEL[8].n2 117.008
R20490 BIT_SEL[8].n1 BIT_SEL[8].t4 117.008
R20491 BIT_SEL[8].n0 BIT_SEL[8].t0 117.008
R20492 a_1340_6292.t0 a_1340_6292.t1 5.92611
R20493 a_20810_48783.t0 a_20810_48783.t1 6.39548
R20494 a_7830_33925.t0 a_7830_33925.t1 6.71904
R20495 a_7830_40009.t0 a_7830_40009.t1 8.49425
R20496 a_20810_61063.t0 a_20810_61063.t1 6.38524
R20497 BIT_SEL[30].n6 BIT_SEL[30] 6.60907
R20498 BIT_SEL[30] BIT_SEL[30].n6 6.01925
R20499 BIT_SEL[30].n6 BIT_SEL[30].t7 118.243
R20500 BIT_SEL[30] BIT_SEL[30].n0 6.01925
R20501 BIT_SEL[30].n0 BIT_SEL[30] 6.60907
R20502 BIT_SEL[30] BIT_SEL[30].n1 6.01925
R20503 BIT_SEL[30].n1 BIT_SEL[30] 6.60907
R20504 BIT_SEL[30] BIT_SEL[30].n2 6.01925
R20505 BIT_SEL[30].n2 BIT_SEL[30] 6.60907
R20506 BIT_SEL[30] BIT_SEL[30].n3 6.01925
R20507 BIT_SEL[30].n3 BIT_SEL[30] 6.60907
R20508 BIT_SEL[30] BIT_SEL[30].n4 6.01925
R20509 BIT_SEL[30].n4 BIT_SEL[30] 6.60907
R20510 BIT_SEL[30] BIT_SEL[30].n5 6.01925
R20511 BIT_SEL[30].n5 BIT_SEL[30] 6.60907
R20512 BIT_SEL[30].t5 BIT_SEL[30] 124.261
R20513 BIT_SEL[30].t0 BIT_SEL[30].n5 118.243
R20514 BIT_SEL[30].t3 BIT_SEL[30].n4 118.243
R20515 BIT_SEL[30].t1 BIT_SEL[30].n3 118.243
R20516 BIT_SEL[30].t6 BIT_SEL[30].n2 118.243
R20517 BIT_SEL[30].t4 BIT_SEL[30].n1 118.243
R20518 BIT_SEL[30].t2 BIT_SEL[30].n0 118.243
R20519 a_7830_54819.t0 a_7830_54819.t1 9.05295
R20520 a_14320_42539.t0 a_14320_42539.t1 6.02155
R20521 a_14320_57028.t0 a_14320_57028.t1 5.92075
R20522 a_1340_50416.t0 a_1340_50416.t1 6.02155
R20523 a_14320_23311.t0 a_14320_23311.t1 9.05295
R20524 a_1340_21678.t0 a_1340_21678.t1 6.38524
R20525 a_20810_24783.t0 a_20810_24783.t1 7.42442
R20526 a_20810_46942.t0 a_20810_46942.t1 9.05337
R20527 a_14320_23887.t0 a_14320_23887.t1 9.52407
R20528 a_20810_40537.t0 a_20810_40537.t1 7.42442
R20529 a_1340_37432.t0 a_1340_37432.t1 6.38524
R20530 a_20810_50416.t0 a_20810_50416.t1 6.02155
R20531 a_7830_49679.t0 a_7830_49679.t1 6.71904
R20532 a_7830_1889.t0 a_7830_1889.t1 5.92117
R20533 a_1340_44412.t0 a_1340_44412.t1 8.02269
R20534 a_14320_48783.t0 a_14320_48783.t1 6.39662
R20535 a_7830_53186.t0 a_7830_53186.t1 6.38524
R20536 a_20810_57925.t0 a_20810_57925.t1 7.5582
R20537 a_14320_55395.t0 a_14320_55395.t1 9.52407
R20538 a_20810_29026.t0 a_20810_29026.t1 7.18213
R20539 a_20810_29923.t0 a_20810_29923.t1 5.92569
R20540 a_7830_53554.t0 a_7830_53554.t1 5.92611
R20541 a_1340_14537.t0 a_1340_14537.t1 6.9546
R20542 a_7830_16906.t0 a_7830_16906.t1 7.42442
R20543 a_14320_55763.t0 a_14320_55763.t1 8.49425
R20544 a_20810_44780.t0 a_20810_44780.t1 7.18213
R20545 a_1340_18540.t0 a_1340_18540.t1 7.55862
R20546 a_1340_41802.t0 a_1340_41802.t1 6.71904
R20547 a_1340_30291.t0 a_1340_30291.t1 6.9546
R20548 BIT_SEL[31].n6 BIT_SEL[31] 6.01764
R20549 BIT_SEL[31] BIT_SEL[31].n6 6.61068
R20550 BIT_SEL[31] BIT_SEL[31].t6 124.466
R20551 BIT_SEL[31].n6 BIT_SEL[31].t7 118.448
R20552 BIT_SEL[31] BIT_SEL[31].n0 6.61068
R20553 BIT_SEL[31].n0 BIT_SEL[31] 6.01764
R20554 BIT_SEL[31] BIT_SEL[31].n1 6.61068
R20555 BIT_SEL[31].n1 BIT_SEL[31] 6.01764
R20556 BIT_SEL[31] BIT_SEL[31].n2 6.61068
R20557 BIT_SEL[31].n2 BIT_SEL[31] 6.01764
R20558 BIT_SEL[31] BIT_SEL[31].n3 6.61068
R20559 BIT_SEL[31].n3 BIT_SEL[31] 6.01764
R20560 BIT_SEL[31] BIT_SEL[31].n4 6.61068
R20561 BIT_SEL[31].n4 BIT_SEL[31] 6.01764
R20562 BIT_SEL[31] BIT_SEL[31].n5 6.61068
R20563 BIT_SEL[31].n5 BIT_SEL[31] 6.01764
R20564 BIT_SEL[31].t3 BIT_SEL[31].n5 118.448
R20565 BIT_SEL[31].t1 BIT_SEL[31].n4 118.448
R20566 BIT_SEL[31].t0 BIT_SEL[31].n3 118.448
R20567 BIT_SEL[31].t5 BIT_SEL[31].n2 118.448
R20568 BIT_SEL[31].t2 BIT_SEL[31].n1 118.448
R20569 BIT_SEL[31].t4 BIT_SEL[31].n0 118.448
R20570 a_154_24425.t0 a_154_24425.t1 13.9628
R20571 a_110_24513.t0 a_110_24513.t1 19.5535
R20572 a_7830_2417.t0 a_7830_2417.t1 6.71904
R20573 a_7830_62328.t0 a_7830_62328.t1 8.02468
R20574 a_1340_46045.t0 a_1340_46045.t1 6.9546
R20575 a_20810_2786.t0 a_20810_2786.t1 7.5582
R20576 a_20718_4081.t0 a_20718_4081.t1 6.66648
R20577 a_110_8311.t0 a_110_8311.t1 19.5535
R20578 a_154_8223.t0 a_154_8223.t1 13.9628
R20579 a_14320_57925.t0 a_14320_57925.t1 7.55862
R20580 a_7830_22046.t0 a_7830_22046.t1 5.92611
R20581 a_14320_29026.t0 a_14320_29026.t1 7.18327
R20582 a_7830_28658.t0 a_7830_28658.t1 8.02156
R20583 a_20810_9029.t0 a_20810_9029.t1 7.42442
R20584 a_20718_59220.t0 a_20718_59220.t1 6.66648
R20585 a_14320_44780.t0 a_14320_44780.t1 7.18327
R20586 a_154_55933.t0 a_154_55933.t1 13.9628
R20587 a_110_56021.t0 a_110_56021.t1 19.5535
R20588 a_1340_52657.t0 a_1340_52657.t1 7.18327
R20589 OUT[5] OUT[5].n0 9.0005
R20590 OUT[5].n0 OUT[5].t1 8.56064
R20591 OUT[5].n0 OUT[5].t0 4.38216
R20592 a_1340_10294.t0 a_1340_10294.t1 6.71904
R20593 a_7830_10663.t0 a_7830_10663.t1 7.5582
R20594 a_20810_23887.t0 a_20810_23887.t1 9.52407
R20595 a_7830_11031.t0 a_7830_11031.t1 6.02155
R20596 a_20810_57028.t0 a_20810_57028.t1 5.92075
R20597 a_20810_23311.t0 a_20810_23311.t1 9.05337
R20598 a_1340_60166.t0 a_1340_60166.t1 8.02269
R20599 a_7830_624.t0 a_7830_624.t1 8.49425
R20600 a_14320_2786.t0 a_14320_2786.t1 7.5582
R20601 a_154_14943.t0 a_154_14943.t1 13.9628
R20602 a_110_15031.t0 a_110_15031.t1 19.5535
R20603 a_7830_53922.t0 a_7830_53922.t1 6.9546
R20604 COL_PROG_N[2] COL_PROG_N[2].n0 0.0965
R20605 COL_PROG_N[2].n0 COL_PROG_N[2].n1 0.3065
R20606 COL_PROG_N[2].n1 COL_PROG_N[2].n2 0.3065
R20607 COL_PROG_N[2].n2 COL_PROG_N[2].t2 292.788
R20608 COL_PROG_N[2].n2 COL_PROG_N[2].t0 292.481
R20609 COL_PROG_N[2].n1 COL_PROG_N[2].t3 292.481
R20610 COL_PROG_N[2].n0 COL_PROG_N[2].t1 292.481
R20611 a_7830_42171.t0 a_7830_42171.t1 7.5582
R20612 a_1340_20781.t0 a_1340_20781.t1 8.02269
R20613 a_14228_27712.t0 a_14228_27712.t1 6.66648
R20614 OUT[1] OUT[1].n0 9.0005
R20615 OUT[1].n0 OUT[1].t1 8.56064
R20616 OUT[1].n0 OUT[1].t0 4.38216
R20617 a_20810_5027.t0 a_20810_5027.t1 8.02269
R20618 COL_PROG_N[6] COL_PROG_N[6].n0 0.0965
R20619 COL_PROG_N[6].n0 COL_PROG_N[6].n1 0.3065
R20620 COL_PROG_N[6].n1 COL_PROG_N[6].n2 0.3065
R20621 COL_PROG_N[6].n2 COL_PROG_N[6].t2 292.788
R20622 COL_PROG_N[6].n2 COL_PROG_N[6].t0 292.481
R20623 COL_PROG_N[6].n1 COL_PROG_N[6].t3 292.481
R20624 COL_PROG_N[6].n0 COL_PROG_N[6].t1 292.481
R20625 a_1340_36903.t0 a_1340_36903.t1 7.18327
R20626 a_7830_9029.t0 a_7830_9029.t1 7.42442
R20627 a_1340_15434.t0 a_1340_15434.t1 9.05337
R20628 a_1340_48414.t0 a_1340_48414.t1 7.42556
R20629 a_7830_30820.t0 a_7830_30820.t1 8.02468
R20630 a_14320_62696.t0 a_14320_62696.t1 9.05295
R20631 a_14320_33029.t0 a_14320_33029.t1 6.39662
R20632 a_7830_56291.t0 a_7830_56291.t1 7.42442
R20633 a_7830_46574.t0 a_7830_46574.t1 8.02468
R20634 a_7830_61799.t0 a_7830_61799.t1 6.9546
R20635 a_1340_26417.t0 a_1340_26417.t1 7.55862
R20636 a_7830_26048.t0 a_7830_26048.t1 6.71904
R20637 a_1340_46942.t0 a_1340_46942.t1 9.05295
R20638 a_7830_47518.t0 a_7830_47518.t1 9.52407
R20639 a_154_45555.t0 a_154_45555.t1 13.9628
R20640 a_110_45643.t0 a_110_45643.t1 19.5535
R20641 a_14320_37800.t0 a_14320_37800.t1 5.92611
R20642 a_14320_3154.t0 a_14320_3154.t1 6.02155
R20643 a_7830_3154.t0 a_7830_3154.t1 6.02155
R20644 a_1340_13801.t0 a_1340_13801.t1 6.38524
R20645 a_1340_21149.t0 a_1340_21149.t1 7.18327
R20646 a_7830_16378.t0 a_7830_16378.t1 8.49425
R20647 a_14320_16010.t0 a_14320_16010.t1 9.52407
R20648 a_14320_31188.t0 a_14320_31188.t1 9.05295
R20649 a_7830_17275.t0 a_7830_17275.t1 6.39662
R20650 a_1340_57556.t0 a_1340_57556.t1 6.71904
R20651 a_7830_32132.t0 a_7830_32132.t1 8.49425
R20652 a_14228_19835.t0 a_14228_19835.t1 6.66648
R20653 a_20810_62696.t0 a_20810_62696.t1 9.05337
R20654 a_1340_58293.t0 a_1340_58293.t1 6.02155
R20655 a_154_39731.t0 a_154_39731.t1 13.9628
R20656 a_110_39819.t0 a_110_39819.t1 19.5535
R20657 a_7830_33029.t0 a_7830_33029.t1 6.39548
R20658 a_14320_31764.t0 a_14320_31764.t1 9.52407
R20659 a_7830_15066.t0 a_7830_15066.t1 8.02468
R20660 a_20810_2417.t0 a_20810_2417.t1 6.71904
R20661 a_1340_45309.t0 a_1340_45309.t1 6.38524
R20662 a_14320_17275.t0 a_14320_17275.t1 6.39662
R20663 a_14228_35589.t0 a_14228_35589.t1 6.66648
R20664 a_20810_256.t0 a_20810_256.t1 9.52407
R20665 a_154_14047.t0 a_154_14047.t1 13.9628
R20666 a_110_14135.t0 a_110_14135.t1 19.5535
R20667 a_14320_7189.t0 a_14320_7189.t1 8.02468
R20668 a_14320_17643.t0 a_14320_17643.t1 5.92075
R20669 a_20810_624.t0 a_20810_624.t1 8.49538
R20670 a_20718_27712.t0 a_20718_27712.t1 6.66648
R20671 a_20810_28658.t0 a_20810_28658.t1 8.02269
R20672 a_7830_24783.t0 a_7830_24783.t1 7.42442
R20673 a_1340_1152.t0 a_1340_1152.t1 7.42442
R20674 a_1340_34294.t0 a_1340_34294.t1 7.55862
R20675 a_7830_40537.t0 a_7830_40537.t1 7.42442
R20676 a_7830_50416.t0 a_7830_50416.t1 6.02155
R20677 a_1340_62328.t0 a_1340_62328.t1 8.02468
R20678 a_14320_52289.t0 a_14320_52289.t1 8.02156
R20679 a_20810_18540.t0 a_20810_18540.t1 7.5582
R20680 a_1340_256.t0 a_1340_256.t1 9.52293
R20681 a_20810_33029.t0 a_20810_33029.t1 6.39548
R20682 a_1340_5027.t0 a_1340_5027.t1 8.02269
R20683 a_7830_57925.t0 a_7830_57925.t1 7.5582
R20684 a_154_59741.t0 a_154_59741.t1 13.9628
R20685 a_110_59829.t0 a_110_59829.t1 19.5535
R20686 a_7830_29026.t0 a_7830_29026.t1 7.18327
R20687 a_14320_33397.t0 a_14320_33397.t1 5.92075
R20688 a_1340_9398.t0 a_1340_9398.t1 6.39548
R20689 a_154_28905.t0 a_154_28905.t1 13.9628
R20690 a_110_28993.t0 a_110_28993.t1 19.5535
R20691 a_14320_6292.t0 a_14320_6292.t1 5.92611
R20692 a_7830_49151.t0 a_7830_49151.t1 5.92117
R20693 a_7830_22943.t0 a_7830_22943.t1 8.02468
R20694 a_154_44659.t0 a_154_44659.t1 13.9628
R20695 a_110_44747.t0 a_110_44747.t1 19.5535
R20696 a_14320_18540.t0 a_14320_18540.t1 7.5582
R20697 a_20810_31188.t0 a_20810_31188.t1 9.05337
R20698 a_14320_8133.t0 a_14320_8133.t1 9.52293
R20699 a_1340_12904.t0 a_1340_12904.t1 8.02269
R20700 a_20810_17275.t0 a_20810_17275.t1 6.39548
R20701 a_7738_59220.t0 a_7738_59220.t1 6.66648
R20702 a_20718_35589.t0 a_20718_35589.t1 6.66648
R20703 a_20810_1889.t0 a_20810_1889.t1 5.92075
R20704 a_20810_17643.t0 a_20810_17643.t1 5.92075
R20705 a_154_13151.t0 a_154_13151.t1 13.9628
R20706 a_110_13239.t0 a_110_13239.t1 19.5535
R20707 a_1340_8501.t0 a_1340_8501.t1 8.49538
R20708 a_20810_56660.t0 a_20810_56660.t1 6.39548
R20709 a_7830_57028.t0 a_7830_57028.t1 5.92117
R20710 a_154_39022.t0 a_154_39022.t1 13.9628
R20711 a_110_39110.t0 a_110_39110.t1 19.5535
R20712 a_1340_60534.t0 a_1340_60534.t1 7.18327
R20713 a_7830_5924.t0 a_7830_5924.t1 6.38524
R20714 a_154_30697.t0 a_154_30697.t1 13.9628
R20715 a_110_30785.t0 a_110_30785.t1 19.5535
R20716 a_7830_7557.t0 a_7830_7557.t1 9.05295
R20717 a_14320_38168.t0 a_14320_38168.t1 6.9546
R20718 a_14320_56660.t0 a_14320_56660.t1 6.39662
R20719 a_7830_55395.t0 a_7830_55395.t1 9.52407
R20720 a_1340_34662.t0 a_1340_34662.t1 6.02155
R20721 a_154_53432.t0 a_154_53432.t1 13.9628
R20722 a_110_53520.t0 a_110_53520.t1 19.5535
R20723 a_20810_33397.t0 a_20810_33397.t1 5.92075
R20724 a_1340_53554.t0 a_1340_53554.t1 5.92569
R20725 a_154_40179.t0 a_154_40179.t1 13.9628
R20726 a_110_40267.t0 a_110_40267.t1 19.5535
R20727 a_14228_11958.t0 a_14228_11958.t1 6.66648
R20728 a_1340_16378.t0 a_1340_16378.t1 8.49425
R20729 a_7830_24255.t0 a_7830_24255.t1 8.49425
R20730 a_154_62205.t0 a_154_62205.t1 13.9628
R20731 a_110_62293.t0 a_110_62293.t1 19.5535
R20732 a_20810_1521.t0 a_20810_1521.t1 6.39548
R20733 a_7830_32660.t0 a_7830_32660.t1 7.42442
R20734 a_154_46899.t0 a_154_46899.t1 13.9628
R20735 a_110_46987.t0 a_110_46987.t1 19.5535
R20736 a_14228_43466.t0 a_14228_43466.t1 6.66648
R20737 a_1340_10663.t0 a_1340_10663.t1 7.55862
R20738 a_154_56381.t0 a_154_56381.t1 13.9628
R20739 a_110_56469.t0 a_110_56469.t1 19.5535
R20740 a_1340_38697.t0 a_1340_38697.t1 8.02468
R20741 a_154_21924.t0 a_154_21924.t1 13.9628
R20742 a_110_22012.t0 a_110_22012.t1 19.5535
R20743 a_14320_25520.t0 a_14320_25520.t1 5.92075
R20744 a_1340_40009.t0 a_1340_40009.t1 8.49538
R20745 a_20810_36535.t0 a_20810_36535.t1 8.02269
R20746 a_1340_54819.t0 a_1340_54819.t1 9.05337
R20747 a_154_15391.t0 a_154_15391.t1 13.9628
R20748 a_110_15479.t0 a_110_15479.t1 19.5535
R20749 a_1340_42171.t0 a_1340_42171.t1 7.55862
R20750 a_1340_47518.t0 a_1340_47518.t1 9.52293
R20751 a_14320_9766.t0 a_14320_9766.t1 5.92117
R20752 a_154_38126.t0 a_154_38126.t1 13.9628
R20753 a_110_38214.t0 a_110_38214.t1 19.5535
R20754 a_14320_29555.t0 a_14320_29555.t1 6.38524
R20755 a_1340_53186.t0 a_1340_53186.t1 6.38524
R20756 a_154_36782.t0 a_154_36782.t1 13.9628
R20757 a_110_36870.t0 a_110_36870.t1 19.5535
R20758 a_1340_16906.t0 a_1340_16906.t1 7.42442
R20759 a_20718_11958.t0 a_20718_11958.t1 6.66648
R20760 a_14320_26417.t0 a_14320_26417.t1 7.5582
R20761 a_7830_62696.t0 a_7830_62696.t1 9.05295
R20762 a_1340_56291.t0 a_1340_56291.t1 7.42442
R20763 a_1248_4081.t0 a_1248_4081.t1 6.66648
R20764 a_20718_43466.t0 a_20718_43466.t1 6.66648
R20765 a_14320_37432.t0 a_14320_37432.t1 6.38524
R20766 a_20810_25520.t0 a_20810_25520.t1 5.92075
R20767 a_14320_1152.t0 a_14320_1152.t1 7.42442
R20768 a_7738_35589.t0 a_7738_35589.t1 6.66648
R20769 a_1340_53922.t0 a_1340_53922.t1 6.9546
R20770 a_20810_29555.t0 a_20810_29555.t1 6.38524
R20771 a_14320_52657.t0 a_14320_52657.t1 7.18327
R20772 a_1340_30820.t0 a_1340_30820.t1 8.02468
R20773 a_1340_46574.t0 a_1340_46574.t1 8.02468
R20774 a_7830_7189.t0 a_7830_7189.t1 8.02468
R20775 a_1340_26048.t0 a_1340_26048.t1 6.71904
R20776 a_20810_44412.t0 a_20810_44412.t1 8.02269
R20777 a_1340_15066.t0 a_1340_15066.t1 8.02468
C0 BIT_SEL[30] BIT_SEL[20] 0.2588f
C1 BIT_SEL[28] BIT_SEL[22] 0.22524f
C2 BIT_SEL[60] BIT_SEL[56] 0.24265f
C3 BIT_SEL[26] BIT_SEL[24] 2.44362f
C4 BIT_SEL[62] BIT_SEL[54] 0.26043f
C5 BIT_SEL[58] BIT_SEL[57] 25.7303f
C6 BIT_SEL[54] BIT_SEL[53] 25.7241f
C7 BIT_SEL[60] BIT_SEL[59] 25.7374f
C8 BIT_SEL[56] BIT_SEL[55] 25.7007f
C9 BIT_SEL[62] BIT_SEL[61] 25.7364f
C10 BIT_SEL[28] BIT_SEL[29] 25.7382f
C11 BIT_SEL[30] BIT_SEL[31] 28.6814f
C12 BIT_SEL[20] BIT_SEL[21] 25.7102f
C13 BIT_SEL[22] BIT_SEL[23] 25.7222f
C14 BIT_SEL[24] BIT_SEL[25] 25.7235f
C15 BIT_SEL[26] BIT_SEL[27] 25.7092f
C16 PRESET_N SENSE 27.1755f
C17 BIT_SEL[16] BIT_SEL[33] 0.01882f
C18 BIT_SEL[21] BIT_SEL[31] 0.28174f
C19 BIT_SEL[55] BIT_SEL[59] 0.28253f
C20 BIT_SEL[23] BIT_SEL[29] 0.27378f
C21 BIT_SEL[25] BIT_SEL[27] 2.58494f
C22 BIT_SEL[53] BIT_SEL[61] 0.26342f
C23 VDD BIT_SEL[60] 0.21883f
C24 BIT_SEL[60] BIT_SEL[32] 0.01882f
C25 BIT_SEL[38] BIT_SEL[54] 1.34627f
C26 BIT_SEL[26] BIT_SEL[0] 0.01882f
C27 BIT_SEL[12] SENSE 0.01155f
C28 VDD BIT_SEL[55] 0.22284f
C29 BIT_SEL[32] BIT_SEL[55] 0.01882f
C30 SENSE BIT_SEL[7] 0.02325f
C31 BIT_SEL[3] BIT_SEL[5] 1.51263f
C32 BIT_SEL[0] BIT_SEL[25] 0.01882f
C33 BIT_SEL[12] BIT_SEL[28] 1.34627f
C34 BIT_SEL[45] BIT_SEL[61] 1.34627f
C35 BIT_SEL[56] BIT_SEL[49] 0.25472f
C36 BIT_SEL[2] BIT_SEL[0] 1.02325f
C37 BIT_SEL[22] BIT_SEL[17] 0.2966f
C38 BIT_SEL[36] BIT_SEL[32] 0.27877f
C39 BIT_SEL[58] BIT_SEL[51] 0.25545f
C40 BIT_SEL[24] BIT_SEL[19] 0.23548f
C41 BIT_SEL[49] BIT_SEL[59] 0.29183f
C42 BIT_SEL[17] BIT_SEL[29] 0.28574f
C43 BIT_SEL[51] BIT_SEL[57] 0.21768f
C44 BIT_SEL[7] BIT_SEL[23] 1.34627f
C45 BIT_SEL[19] BIT_SEL[27] 0.25726f
C46 BIT_SEL[32] BIT_SEL[47] 0.28034f
C47 BIT_SEL[42] BIT_SEL[40] 2.44362f
C48 BIT_SEL[44] BIT_SEL[38] 0.22524f
C49 BIT_SEL[46] BIT_SEL[36] 0.2588f
C50 BIT_SEL[12] BIT_SEL[4] 0.23829f
C51 BIT_SEL[10] BIT_SEL[6] 0.27079f
C52 BIT_SEL[14] BIT_SEL[2] 0.2614f
C53 VDD BIT_SEL[49] 0.26125f
C54 BIT_SEL[32] BIT_SEL[49] 0.01882f
C55 BIT_SEL[40] BIT_SEL[41] 25.7235f
C56 BIT_SEL[36] BIT_SEL[37] 25.7102f
C57 BIT_SEL[44] BIT_SEL[45] 25.7382f
C58 BIT_SEL[38] BIT_SEL[39] 25.7222f
C59 BIT_SEL[46] BIT_SEL[47] 28.6814f
C60 BIT_SEL[42] BIT_SEL[43] 25.7092f
C61 BIT_SEL[6] BIT_SEL[9] 0.26576f
C62 BIT_SEL[10] BIT_SEL[13] 0.2575f
C63 BIT_SEL[8] BIT_SEL[11] 0.23092f
C64 BIT_SEL[0] BIT_SEL[19] 0.01882f
C65 BIT_SEL[4] BIT_SEL[7] 0.25036f
C66 BIT_SEL[12] BIT_SEL[15] 0.35892f
C67 BIT_SEL[39] BIT_SEL[45] 0.27378f
C68 BIT_SEL[37] BIT_SEL[47] 0.28174f
C69 BIT_SEL[7] BIT_SEL[15] 0.29084f
C70 BIT_SEL[9] BIT_SEL[13] 0.28151f
C71 BIT_SEL[41] BIT_SEL[43] 2.58494f
C72 BIT_SEL[42] BIT_SEL[16] 0.01882f
C73 COL_PROG_N[7] COL_PROG_N[6] 0.13261f
C74 BIT_SEL[16] BIT_SEL[41] 0.01882f
C75 VDD OUT[6] 0.257f
C76 BIT_SEL[28] BIT_SEL[44] 1.34627f
C77 VDD BIT_SEL[2] 0.01126f
C78 BIT_SEL[18] BIT_SEL[16] 1.02325f
C79 BIT_SEL[52] BIT_SEL[48] 0.27877f
C80 BIT_SEL[40] BIT_SEL[35] 0.23548f
C81 BIT_SEL[6] BIT_SEL[3] 0.27726f
C82 BIT_SEL[4] BIT_SEL[1] 0.28401f
C83 BIT_SEL[8] BIT_SEL[5] 0.22247f
C84 BIT_SEL[38] BIT_SEL[33] 0.2966f
C85 VDD COL_PROG_N[6] 3.59445f
C86 BIT_SEL[23] BIT_SEL[39] 1.34627f
C87 BIT_SEL[35] BIT_SEL[43] 0.25726f
C88 BIT_SEL[1] BIT_SEL[15] 0.30282f
C89 BIT_SEL[48] BIT_SEL[63] 0.28034f
C90 BIT_SEL[3] BIT_SEL[13] 0.24884f
C91 BIT_SEL[5] BIT_SEL[11] 0.27685f
C92 BIT_SEL[33] BIT_SEL[45] 0.28574f
C93 VDD OUT[4] 0.257f
C94 BIT_SEL[60] BIT_SEL[54] 0.22524f
C95 BIT_SEL[28] BIT_SEL[20] 0.23829f
C96 BIT_SEL[58] BIT_SEL[56] 2.44362f
C97 BIT_SEL[62] BIT_SEL[52] 0.2588f
C98 BIT_SEL[26] BIT_SEL[22] 0.27079f
C99 BIT_SEL[30] BIT_SEL[18] 0.2614f
C100 BIT_SEL[60] BIT_SEL[61] 25.7382f
C101 BIT_SEL[54] BIT_SEL[55] 25.7222f
C102 BIT_SEL[1] BIT_SEL[17] 1.33981f
C103 BIT_SEL[58] BIT_SEL[59] 25.7092f
C104 BIT_SEL[56] BIT_SEL[57] 25.7235f
C105 BIT_SEL[52] BIT_SEL[53] 25.7102f
C106 BIT_SEL[24] BIT_SEL[27] 0.23092f
C107 BIT_SEL[18] BIT_SEL[21] 0.23368f
C108 BIT_SEL[20] BIT_SEL[23] 0.25036f
C109 BIT_SEL[26] BIT_SEL[29] 0.2575f
C110 BIT_SEL[28] BIT_SEL[31] 0.35892f
C111 BIT_SEL[22] BIT_SEL[25] 0.26576f
C112 BIT_SEL[62] BIT_SEL[63] 28.6814f
C113 BIT_SEL[16] BIT_SEL[35] 0.01882f
C114 VDD COL_PROG_N[4] 3.59445f
C115 BIT_SEL[53] BIT_SEL[63] 0.28174f
C116 BIT_SEL[25] BIT_SEL[29] 0.28151f
C117 BIT_SEL[55] BIT_SEL[61] 0.27378f
C118 BIT_SEL[23] BIT_SEL[31] 0.29084f
C119 BIT_SEL[57] BIT_SEL[59] 2.58494f
C120 VDD BIT_SEL[58] 0.21883f
C121 BIT_SEL[10] SENSE 0.01069f
C122 BIT_SEL[58] BIT_SEL[32] 0.01882f
C123 BIT_SEL[24] BIT_SEL[0] 0.01882f
C124 VDD OUT[2] 0.257f
C125 BIT_SEL[4] BIT_SEL[20] 1.34627f
C126 VDD BIT_SEL[57] 0.22141f
C127 BIT_SEL[0] BIT_SEL[27] 0.01882f
C128 SENSE BIT_SEL[9] 0.01999f
C129 BIT_SEL[32] BIT_SEL[57] 0.01882f
C130 PRESET_N OUT[6] 0.01765f
C131 BIT_SEL[48] COL_PROG_N[5] 0.06116f
C132 BIT_SEL[44] BIT_SEL[60] 1.34627f
C133 VDD COL_PROG_N[2] 3.59445f
C134 BIT_SEL[15] BIT_SEL[31] 1.34627f
C135 BIT_SEL[20] BIT_SEL[17] 0.28401f
C136 VDD OUT[0] 0.257f
C137 BIT_SEL[56] BIT_SEL[51] 0.23548f
C138 BIT_SEL[22] BIT_SEL[19] 0.27726f
C139 BIT_SEL[54] BIT_SEL[49] 0.2966f
C140 BIT_SEL[34] BIT_SEL[32] 1.02325f
C141 BIT_SEL[51] BIT_SEL[59] 0.25726f
C142 BIT_SEL[17] BIT_SEL[31] 0.30282f
C143 BIT_SEL[49] BIT_SEL[61] 0.28574f
C144 BIT_SEL[19] BIT_SEL[29] 0.24884f
C145 BIT_SEL[39] BIT_SEL[55] 1.34627f
C146 BIT_SEL[44] BIT_SEL[36] 0.23829f
C147 BIT_SEL[8] BIT_SEL[6] 2.05426f
C148 BIT_SEL[42] BIT_SEL[38] 0.27079f
C149 PRESET_N OUT[4] 0.01765f
C150 BIT_SEL[46] BIT_SEL[34] 0.2614f
C151 BIT_SEL[48] COL_PROG_N[3] 0.06116f
C152 BIT_SEL[10] BIT_SEL[4] 0.27323f
C153 BIT_SEL[12] BIT_SEL[2] 0.24323f
C154 BIT_SEL[14] BIT_SEL[0] 0.23787f
C155 VDD COL_PROG_N[0] 3.59535f
C156 VDD BIT_SEL[51] 0.2352f
C157 BIT_SEL[8] BIT_SEL[13] 0.25358f
C158 BIT_SEL[10] BIT_SEL[15] 0.35033f
C159 BIT_SEL[2] BIT_SEL[7] 0.24224f
C160 BIT_SEL[40] BIT_SEL[43] 0.23092f
C161 BIT_SEL[36] BIT_SEL[39] 0.25036f
C162 BIT_SEL[42] BIT_SEL[45] 0.2575f
C163 BIT_SEL[44] BIT_SEL[47] 0.35892f
C164 BIT_SEL[4] BIT_SEL[9] 0.25414f
C165 BIT_SEL[38] BIT_SEL[41] 0.26576f
C166 BIT_SEL[32] BIT_SEL[51] 0.01882f
C167 BIT_SEL[34] BIT_SEL[37] 0.23368f
C168 BIT_SEL[17] BIT_SEL[33] 1.33981f
C169 BIT_SEL[6] BIT_SEL[11] 0.24182f
C170 BIT_SEL[41] BIT_SEL[45] 0.28151f
C171 BIT_SEL[39] BIT_SEL[47] 0.29084f
C172 BIT_SEL[11] BIT_SEL[13] 2.17343f
C173 BIT_SEL[9] BIT_SEL[15] 0.31315f
C174 SENSE OUT[5] 0.05922f
C175 BIT_SEL[20] BIT_SEL[36] 1.34627f
C176 BIT_SEL[40] BIT_SEL[16] 0.01882f
C177 PRESET_N OUT[2] 0.01765f
C178 BIT_SEL[48] COL_PROG_N[1] 0.06116f
C179 BIT_SEL[16] BIT_SEL[43] 0.01882f
C180 BIT_SEL[5] BIT_SEL[21] 1.34627f
C181 BIT_SEL[31] BIT_SEL[47] 1.34627f
C182 SENSE OUT[3] 0.05922f
C183 BIT_SEL[38] BIT_SEL[35] 0.27726f
C184 BIT_SEL[2] BIT_SEL[1] 25.7321f
C185 BIT_SEL[6] BIT_SEL[5] 25.7241f
C186 BIT_SEL[50] BIT_SEL[48] 1.02325f
C187 BIT_SEL[4] BIT_SEL[3] 25.7336f
C188 BIT_SEL[36] BIT_SEL[33] 0.28401f
C189 PRESET_N OUT[0] 0.01765f
C190 BIT_SEL[3] BIT_SEL[15] 0.2831f
C191 BIT_SEL[33] BIT_SEL[47] 0.30282f
C192 BIT_SEL[5] BIT_SEL[13] 0.26342f
C193 BIT_SEL[35] BIT_SEL[45] 0.24884f
C194 BIT_SEL[58] BIT_SEL[54] 0.27079f
C195 BIT_SEL[28] BIT_SEL[18] 0.24323f
C196 BIT_SEL[24] BIT_SEL[22] 2.05426f
C197 BIT_SEL[60] BIT_SEL[52] 0.23829f
C198 BIT_SEL[62] BIT_SEL[50] 0.2614f
C199 BIT_SEL[26] BIT_SEL[20] 0.27323f
C200 BIT_SEL[30] BIT_SEL[16] 0.23787f
C201 SENSE OUT[1] 0.05922f
C202 VDD OUT[7] 0.257f
C203 BIT_SEL[52] BIT_SEL[55] 0.25036f
C204 BIT_SEL[18] BIT_SEL[23] 0.24224f
C205 BIT_SEL[16] BIT_SEL[21] 0.229f
C206 BIT_SEL[24] BIT_SEL[29] 0.25358f
C207 BIT_SEL[56] BIT_SEL[59] 0.23092f
C208 BIT_SEL[33] BIT_SEL[49] 1.33981f
C209 BIT_SEL[22] BIT_SEL[27] 0.24182f
C210 BIT_SEL[60] BIT_SEL[63] 0.35892f
C211 BIT_SEL[20] BIT_SEL[25] 0.25414f
C212 BIT_SEL[58] BIT_SEL[61] 0.2575f
C213 BIT_SEL[54] BIT_SEL[57] 0.26576f
C214 BIT_SEL[50] BIT_SEL[53] 0.23368f
C215 BIT_SEL[26] BIT_SEL[31] 0.35033f
C216 VDD COL_PROG_N[7] 3.45446f
C217 BIT_SEL[55] BIT_SEL[63] 0.29084f
C218 BIT_SEL[27] BIT_SEL[29] 2.17343f
C219 BIT_SEL[57] BIT_SEL[61] 0.28151f
C220 BIT_SEL[25] BIT_SEL[31] 0.31315f
C221 VDD BIT_SEL[56] 0.2843f
C222 BIT_SEL[56] BIT_SEL[32] 0.01882f
C223 BIT_SEL[8] SENSE 0.0229f
C224 BIT_SEL[22] BIT_SEL[0] 0.01882f
C225 BIT_SEL[36] BIT_SEL[52] 1.34627f
C226 BIT_SEL[30] BIT_SEL[21] 0.23012f
C227 VDD BIT_SEL[59] 0.29023f
C228 SENSE BIT_SEL[11] 0.02295f
C229 BIT_SEL[0] BIT_SEL[29] 0.01882f
C230 BIT_SEL[32] BIT_SEL[59] 0.01882f
C231 BIT_SEL[10] BIT_SEL[26] 1.34627f
C232 BIT_SEL[47] BIT_SEL[63] 1.34627f
C233 BIT_SEL[52] BIT_SEL[49] 0.28401f
C234 BIT_SEL[54] BIT_SEL[51] 0.27726f
C235 BIT_SEL[20] BIT_SEL[19] 25.7336f
C236 BIT_SEL[18] BIT_SEL[17] 25.7321f
C237 BIT_SEL[9] BIT_SEL[25] 1.34627f
C238 BIT_SEL[51] BIT_SEL[61] 0.24884f
C239 BIT_SEL[49] BIT_SEL[63] 0.30282f
C240 BIT_SEL[19] BIT_SEL[31] 0.2831f
C241 BIT_SEL[42] BIT_SEL[36] 0.27323f
C242 BIT_SEL[44] BIT_SEL[34] 0.24323f
C243 BIT_SEL[46] BIT_SEL[32] 0.23787f
C244 BIT_SEL[12] BIT_SEL[0] 0.22623f
C245 BIT_SEL[10] BIT_SEL[2] 0.27106f
C246 BIT_SEL[8] BIT_SEL[4] 0.27301f
C247 BIT_SEL[40] BIT_SEL[38] 2.05426f
C248 BIT_SEL[0] BIT_SEL[7] 0.24037f
C249 BIT_SEL[6] BIT_SEL[13] 0.25287f
C250 BIT_SEL[36] BIT_SEL[41] 0.25414f
C251 BIT_SEL[8] BIT_SEL[15] 0.31694f
C252 BIT_SEL[32] BIT_SEL[37] 0.229f
C253 BIT_SEL[38] BIT_SEL[43] 0.24182f
C254 BIT_SEL[42] BIT_SEL[47] 0.35033f
C255 PRESET_N OUT[7] 0.01765f
C256 BIT_SEL[2] BIT_SEL[9] 0.24873f
C257 BIT_SEL[4] BIT_SEL[11] 0.2329f
C258 BIT_SEL[34] BIT_SEL[39] 0.24224f
C259 BIT_SEL[40] BIT_SEL[45] 0.25358f
C260 BIT_SEL[14] BIT_SEL[12] 3.17801f
C261 BIT_SEL[11] BIT_SEL[15] 0.3627f
C262 BIT_SEL[43] BIT_SEL[45] 2.17343f
C263 BIT_SEL[41] BIT_SEL[47] 0.31315f
C264 BIT_SEL[46] BIT_SEL[37] 0.23012f
C265 BIT_SEL[38] BIT_SEL[16] 0.01882f
C266 BIT_SEL[14] BIT_SEL[7] 0.22988f
C267 BIT_SEL[16] BIT_SEL[45] 0.01882f
C268 BIT_SEL[26] BIT_SEL[42] 1.34627f
C269 VDD PRESET_N 18.9795f
C270 BIT_SEL[0] BIT_SEL[1] 25.8271f
C271 BIT_SEL[34] BIT_SEL[33] 25.7321f
C272 BIT_SEL[2] BIT_SEL[3] 25.7305f
C273 BIT_SEL[4] BIT_SEL[5] 25.7102f
C274 BIT_SEL[36] BIT_SEL[35] 25.7336f
C275 BIT_SEL[35] BIT_SEL[47] 0.2831f
C276 BIT_SEL[25] BIT_SEL[41] 1.34627f
C277 BIT_SEL[5] BIT_SEL[15] 0.28174f
C278 BIT_SEL[24] BIT_SEL[20] 0.27301f
C279 BIT_SEL[60] BIT_SEL[50] 0.24323f
C280 BIT_SEL[56] BIT_SEL[54] 2.05426f
C281 BIT_SEL[58] BIT_SEL[52] 0.27323f
C282 BIT_SEL[62] BIT_SEL[48] 0.23787f
C283 BIT_SEL[26] BIT_SEL[18] 0.27106f
C284 BIT_SEL[14] BIT_SEL[1] 0.25111f
C285 BIT_SEL[28] BIT_SEL[16] 0.22623f
C286 VDD BIT_SEL[7] 0.01085f
C287 BIT_SEL[20] BIT_SEL[27] 0.2329f
C288 BIT_SEL[3] BIT_SEL[19] 1.34627f
C289 BIT_SEL[58] BIT_SEL[63] 0.35033f
C290 BIT_SEL[18] BIT_SEL[25] 0.24873f
C291 BIT_SEL[22] BIT_SEL[29] 0.25287f
C292 BIT_SEL[24] BIT_SEL[31] 0.31694f
C293 BIT_SEL[48] BIT_SEL[53] 0.229f
C294 BIT_SEL[56] BIT_SEL[61] 0.25358f
C295 BIT_SEL[50] BIT_SEL[55] 0.24224f
C296 BIT_SEL[54] BIT_SEL[59] 0.24182f
C297 BIT_SEL[52] BIT_SEL[57] 0.25414f
C298 BIT_SEL[16] BIT_SEL[23] 0.24037f
C299 BIT_SEL[30] BIT_SEL[28] 3.17801f
C300 BIT_SEL[27] BIT_SEL[31] 0.3627f
C301 BIT_SEL[59] BIT_SEL[61] 2.17343f
C302 BIT_SEL[57] BIT_SEL[63] 0.31315f
C303 VDD BIT_SEL[54] 0.22372f
C304 COL_PROG_N[6] COL_PROG_N[5] 0.13261f
C305 BIT_SEL[28] BIT_SEL[21] 0.25476f
C306 BIT_SEL[62] BIT_SEL[53] 0.23012f
C307 BIT_SEL[20] BIT_SEL[0] 0.01882f
C308 BIT_SEL[6] SENSE 0.02324f
C309 BIT_SEL[30] BIT_SEL[23] 0.22988f
C310 BIT_SEL[54] BIT_SEL[32] 0.01882f
C311 BIT_SEL[2] BIT_SEL[18] 1.34627f
C312 VDD BIT_SEL[61] 0.22385f
C313 BIT_SEL[21] BIT_SEL[23] 1.38186f
C314 SENSE BIT_SEL[13] 0.0227f
C315 BIT_SEL[0] BIT_SEL[31] 0.01882f
C316 BIT_SEL[32] BIT_SEL[61] 0.01882f
C317 BIT_SEL[42] BIT_SEL[58] 1.34627f
C318 BIT_SEL[18] BIT_SEL[19] 25.7305f
C319 BIT_SEL[52] BIT_SEL[51] 25.7336f
C320 BIT_SEL[16] BIT_SEL[17] 25.8271f
C321 BIT_SEL[50] BIT_SEL[49] 25.7321f
C322 COL_PROG_N[5] COL_PROG_N[4] 0.13261f
C323 BIT_SEL[51] BIT_SEL[63] 0.2831f
C324 BIT_SEL[41] BIT_SEL[57] 1.34627f
C325 BIT_SEL[6] BIT_SEL[4] 1.21257f
C326 BIT_SEL[8] BIT_SEL[2] 0.27227f
C327 BIT_SEL[30] BIT_SEL[17] 0.25111f
C328 BIT_SEL[44] BIT_SEL[32] 0.22623f
C329 BIT_SEL[42] BIT_SEL[34] 0.27106f
C330 BIT_SEL[10] BIT_SEL[0] 0.25042f
C331 BIT_SEL[40] BIT_SEL[36] 0.27301f
C332 BIT_SEL[40] BIT_SEL[47] 0.31694f
C333 BIT_SEL[38] BIT_SEL[45] 0.25287f
C334 BIT_SEL[36] BIT_SEL[43] 0.2329f
C335 BIT_SEL[0] BIT_SEL[9] 0.24167f
C336 BIT_SEL[6] BIT_SEL[15] 0.30037f
C337 BIT_SEL[32] BIT_SEL[39] 0.24037f
C338 BIT_SEL[34] BIT_SEL[41] 0.24873f
C339 BIT_SEL[17] BIT_SEL[21] 0.30911f
C340 BIT_SEL[2] BIT_SEL[11] 0.22817f
C341 BIT_SEL[4] BIT_SEL[13] 0.24463f
C342 BIT_SEL[19] BIT_SEL[35] 1.34627f
C343 COL_PROG_N[4] COL_PROG_N[3] 0.13261f
C344 BIT_SEL[46] BIT_SEL[44] 3.17801f
C345 BIT_SEL[14] BIT_SEL[10] 0.27077f
C346 BIT_SEL[13] BIT_SEL[15] 3.44717f
C347 BIT_SEL[43] BIT_SEL[47] 0.3627f
C348 BIT_SEL[44] BIT_SEL[37] 0.25476f
C349 BIT_SEL[36] BIT_SEL[16] 0.01882f
C350 BIT_SEL[14] BIT_SEL[9] 0.23081f
C351 BIT_SEL[46] BIT_SEL[39] 0.22988f
C352 BIT_SEL[12] BIT_SEL[7] 0.26185f
C353 BIT_SEL[18] BIT_SEL[34] 1.34627f
C354 BIT_SEL[37] BIT_SEL[39] 1.38186f
C355 BIT_SEL[16] BIT_SEL[47] 0.01882f
C356 COL_PROG_N[3] COL_PROG_N[2] 0.13261f
C357 BIT_SEL[2] BIT_SEL[5] 0.23368f
C358 BIT_SEL[32] BIT_SEL[33] 25.8271f
C359 BIT_SEL[34] BIT_SEL[35] 25.7305f
C360 BIT_SEL[0] BIT_SEL[3] 0.25101f
C361 COL_PROG_N[2] COL_PROG_N[1] 0.13261f
C362 BIT_SEL[26] BIT_SEL[16] 0.25042f
C363 BIT_SEL[56] BIT_SEL[52] 0.27301f
C364 BIT_SEL[22] BIT_SEL[20] 1.21257f
C365 BIT_SEL[14] BIT_SEL[3] 0.23152f
C366 BIT_SEL[12] BIT_SEL[1] 0.29412f
C367 BIT_SEL[24] BIT_SEL[18] 0.27227f
C368 BIT_SEL[58] BIT_SEL[50] 0.27106f
C369 BIT_SEL[60] BIT_SEL[48] 0.22623f
C370 BIT_SEL[46] BIT_SEL[33] 0.25111f
C371 BIT_SEL[20] BIT_SEL[29] 0.24463f
C372 BIT_SEL[16] BIT_SEL[25] 0.24167f
C373 BIT_SEL[56] BIT_SEL[63] 0.31694f
C374 BIT_SEL[54] BIT_SEL[61] 0.25287f
C375 BIT_SEL[50] BIT_SEL[57] 0.24873f
C376 BIT_SEL[22] BIT_SEL[31] 0.30037f
C377 BIT_SEL[48] BIT_SEL[55] 0.24037f
C378 BIT_SEL[33] BIT_SEL[37] 0.30911f
C379 BIT_SEL[35] BIT_SEL[51] 1.34627f
C380 BIT_SEL[1] BIT_SEL[7] 0.29767f
C381 BIT_SEL[18] BIT_SEL[27] 0.22817f
C382 BIT_SEL[52] BIT_SEL[59] 0.2329f
C383 BIT_SEL[62] BIT_SEL[60] 3.17801f
C384 BIT_SEL[30] BIT_SEL[26] 0.27077f
C385 BIT_SEL[59] BIT_SEL[63] 0.3627f
C386 BIT_SEL[29] BIT_SEL[31] 3.44717f
C387 VDD BIT_SEL[52] 0.23144f
C388 COL_PROG_N[1] COL_PROG_N[0] 0.13261f
C389 BIT_SEL[26] BIT_SEL[21] 0.23973f
C390 BIT_SEL[4] SENSE 0.01076f
C391 BIT_SEL[60] BIT_SEL[53] 0.25476f
C392 BIT_SEL[34] BIT_SEL[50] 1.34627f
C393 BIT_SEL[28] BIT_SEL[23] 0.26185f
C394 BIT_SEL[30] BIT_SEL[25] 0.23081f
C395 BIT_SEL[18] BIT_SEL[0] 0.01882f
C396 BIT_SEL[62] BIT_SEL[55] 0.22988f
C397 BIT_SEL[52] BIT_SEL[32] 0.01882f
C398 VDD BIT_SEL[63] 0.24979f
C399 BIT_SEL[32] BIT_SEL[63] 0.01882f
C400 BIT_SEL[21] BIT_SEL[25] 0.23468f
C401 BIT_SEL[53] BIT_SEL[55] 1.38186f
C402 BIT_SEL[8] BIT_SEL[24] 1.34627f
C403 BIT_SEL[16] BIT_SEL[19] 0.25101f
C404 BIT_SEL[50] BIT_SEL[51] 25.7305f
C405 BIT_SEL[48] BIT_SEL[49] 25.8271f
C406 VDD OUT[5] 0.257f
C407 BIT_SEL[11] BIT_SEL[27] 1.34627f
C408 BIT_SEL[8] BIT_SEL[0] 0.24444f
C409 BIT_SEL[38] BIT_SEL[36] 1.21257f
C410 BIT_SEL[40] BIT_SEL[34] 0.27227f
C411 BIT_SEL[6] BIT_SEL[2] 0.2473f
C412 BIT_SEL[28] BIT_SEL[17] 0.29412f
C413 BIT_SEL[42] BIT_SEL[32] 0.25042f
C414 BIT_SEL[30] BIT_SEL[19] 0.23152f
C415 BIT_SEL[62] BIT_SEL[49] 0.25111f
C416 BIT_SEL[36] BIT_SEL[45] 0.24463f
C417 BIT_SEL[2] BIT_SEL[13] 0.24013f
C418 BIT_SEL[19] BIT_SEL[21] 1.51263f
C419 BIT_SEL[49] BIT_SEL[53] 0.30911f
C420 BIT_SEL[4] BIT_SEL[15] 0.30114f
C421 BIT_SEL[38] BIT_SEL[47] 0.30037f
C422 BIT_SEL[17] BIT_SEL[23] 0.29767f
C423 BIT_SEL[32] BIT_SEL[41] 0.24167f
C424 BIT_SEL[34] BIT_SEL[43] 0.22817f
C425 BIT_SEL[0] BIT_SEL[11] 0.22736f
C426 VDD COL_PROG_N[5] 3.59445f
C427 BIT_SEL[12] BIT_SEL[10] 1.9907f
C428 BIT_SEL[46] BIT_SEL[42] 0.27077f
C429 BIT_SEL[14] BIT_SEL[8] 0.26507f
C430 BIT_SEL[45] BIT_SEL[47] 3.44717f
C431 VDD OUT[3] 0.257f
C432 BIT_SEL[44] BIT_SEL[39] 0.26185f
C433 BIT_SEL[42] BIT_SEL[37] 0.23973f
C434 BIT_SEL[46] BIT_SEL[41] 0.23081f
C435 BIT_SEL[14] BIT_SEL[11] 0.26348f
C436 BIT_SEL[34] BIT_SEL[16] 0.01882f
C437 BIT_SEL[10] BIT_SEL[7] 0.24953f
C438 BIT_SEL[12] BIT_SEL[9] 0.27368f
C439 BIT_SEL[37] BIT_SEL[41] 0.23468f
C440 BIT_SEL[7] BIT_SEL[9] 2.1937f
C441 BIT_SEL[48] COL_PROG_N[6] 0.06116f
C442 VDD COL_PROG_N[3] 3.59445f
C443 BIT_SEL[24] BIT_SEL[40] 1.34627f
C444 VDD OUT[1] 0.257f
C445 BIT_SEL[0] BIT_SEL[5] 0.229f
C446 BIT_SEL[32] BIT_SEL[35] 0.25101f
C447 BIT_SEL[27] BIT_SEL[43] 1.34627f
C448 BIT_SEL[48] COL_PROG_N[4] 0.06116f
C449 PRESET_N OUT[5] 0.01765f
C450 BIT_SEL[12] BIT_SEL[3] 0.27116f
C451 VDD COL_PROG_N[1] 3.59445f
C452 BIT_SEL[10] BIT_SEL[1] 0.27818f
C453 BIT_SEL[24] BIT_SEL[16] 0.24444f
C454 BIT_SEL[58] BIT_SEL[48] 0.25042f
C455 BIT_SEL[14] BIT_SEL[5] 0.23012f
C456 BIT_SEL[44] BIT_SEL[33] 0.29412f
C457 BIT_SEL[54] BIT_SEL[52] 1.21257f
C458 BIT_SEL[56] BIT_SEL[50] 0.27227f
C459 BIT_SEL[46] BIT_SEL[35] 0.23152f
C460 BIT_SEL[22] BIT_SEL[18] 0.2473f
C461 BIT_SEL[33] BIT_SEL[39] 0.29767f
C462 BIT_SEL[1] BIT_SEL[9] 0.25124f
C463 BIT_SEL[20] BIT_SEL[31] 0.30114f
C464 BIT_SEL[48] BIT_SEL[57] 0.24167f
C465 BIT_SEL[3] BIT_SEL[7] 0.26814f
C466 BIT_SEL[52] BIT_SEL[61] 0.24463f
C467 BIT_SEL[50] BIT_SEL[59] 0.22817f
C468 BIT_SEL[16] BIT_SEL[27] 0.22736f
C469 BIT_SEL[18] BIT_SEL[29] 0.24013f
C470 BIT_SEL[35] BIT_SEL[37] 1.51263f
C471 BIT_SEL[54] BIT_SEL[63] 0.30037f
C472 SENSE OUT[6] 0.05922f
C473 BIT_SEL[30] BIT_SEL[24] 0.26507f
C474 BIT_SEL[28] BIT_SEL[26] 1.9907f
C475 BIT_SEL[62] BIT_SEL[58] 0.27077f
C476 BIT_SEL[61] BIT_SEL[63] 3.44717f
C477 BIT_SEL[48] COL_PROG_N[2] 0.06116f
C478 PRESET_N OUT[3] 0.01765f
C479 VDD BIT_SEL[50] 0.24084f
C480 BIT_SEL[26] BIT_SEL[23] 0.24953f
C481 BIT_SEL[58] BIT_SEL[53] 0.23973f
C482 BIT_SEL[30] BIT_SEL[27] 0.26348f
C483 BIT_SEL[60] BIT_SEL[55] 0.26185f
C484 BIT_SEL[2] SENSE 0.02316f
C485 BIT_SEL[50] BIT_SEL[32] 0.01882f
C486 BIT_SEL[62] BIT_SEL[57] 0.23081f
C487 BIT_SEL[0] BIT_SEL[16] 1.35136f
C488 BIT_SEL[24] BIT_SEL[21] 0.22247f
C489 BIT_SEL[28] BIT_SEL[25] 0.27368f
C490 BIT_SEL[23] BIT_SEL[25] 2.1937f
C491 BIT_SEL[53] BIT_SEL[57] 0.23468f
C492 BIT_SEL[21] BIT_SEL[27] 0.27685f
C493 SENSE OUT[4] 0.05922f
C494 BIT_SEL[30] BIT_SEL[0] 0.01882f
C495 BIT_SEL[40] BIT_SEL[56] 1.34627f
C496 BIT_SEL[48] COL_PROG_N[0] 0.06116f
C497 PRESET_N OUT[1] 0.01765f
C498 BIT_SEL[1] BIT_SEL[3] 1.14059f
C499 BIT_SEL[0] BIT_SEL[21] 0.01882f
C500 BIT_SEL[48] BIT_SEL[51] 0.25101f
C501 BIT_SEL[14] BIT_SEL[30] 1.34627f
C502 BIT_SEL[43] BIT_SEL[59] 1.34627f
C503 BIT_SEL[4] BIT_SEL[2] 1.37487f
C504 BIT_SEL[62] BIT_SEL[51] 0.23152f
C505 BIT_SEL[40] BIT_SEL[32] 0.24444f
C506 BIT_SEL[6] BIT_SEL[0] 0.22864f
C507 BIT_SEL[60] BIT_SEL[49] 0.29412f
C508 BIT_SEL[38] BIT_SEL[34] 0.2473f
C509 BIT_SEL[26] BIT_SEL[17] 0.27818f
C510 BIT_SEL[28] BIT_SEL[19] 0.27116f
C511 SENSE OUT[2] 0.05922f
C512 BIT_SEL[19] BIT_SEL[23] 0.26814f
C513 BIT_SEL[0] BIT_SEL[13] 0.23927f
C514 BIT_SEL[49] BIT_SEL[55] 0.29767f
C515 BIT_SEL[36] BIT_SEL[47] 0.30114f
C516 BIT_SEL[34] BIT_SEL[45] 0.24013f
C517 BIT_SEL[2] BIT_SEL[15] 0.30342f
C518 BIT_SEL[51] BIT_SEL[53] 1.51263f
C519 BIT_SEL[17] BIT_SEL[25] 0.25124f
C520 BIT_SEL[32] BIT_SEL[43] 0.22736f
C521 BIT_SEL[44] BIT_SEL[42] 1.9907f
C522 BIT_SEL[12] BIT_SEL[8] 0.24265f
C523 BIT_SEL[46] BIT_SEL[40] 0.26507f
C524 BIT_SEL[14] BIT_SEL[6] 0.26043f
C525 BIT_SEL[8] BIT_SEL[7] 25.7007f
C526 BIT_SEL[10] BIT_SEL[9] 25.7303f
C527 BIT_SEL[12] BIT_SEL[11] 25.7374f
C528 BIT_SEL[44] BIT_SEL[41] 0.27368f
C529 BIT_SEL[42] BIT_SEL[39] 0.24953f
C530 BIT_SEL[46] BIT_SEL[43] 0.26348f
C531 BIT_SEL[16] BIT_SEL[32] 1.35136f
C532 BIT_SEL[14] BIT_SEL[13] 25.7364f
C533 BIT_SEL[40] BIT_SEL[37] 0.22247f
C534 SENSE OUT[0] 0.05922f
C535 BIT_SEL[37] BIT_SEL[43] 0.27685f
C536 BIT_SEL[39] BIT_SEL[41] 2.1937f
C537 BIT_SEL[7] BIT_SEL[11] 0.28253f
C538 BIT_SEL[46] BIT_SEL[16] 0.01882f
C539 BIT_SEL[16] BIT_SEL[37] 0.01882f
C540 BIT_SEL[17] BIT_SEL[19] 1.14059f
C541 BIT_SEL[30] BIT_SEL[46] 1.34627f
C542 COL_PROG_N[7] BIT_SEL[48] 0.06046f
C543 VDD BIT_SEL[6] 0.01062f
C544 BIT_SEL[42] BIT_SEL[33] 0.27818f
C545 BIT_SEL[10] BIT_SEL[3] 0.25545f
C546 BIT_SEL[12] BIT_SEL[5] 0.25476f
C547 BIT_SEL[54] BIT_SEL[50] 0.2473f
C548 BIT_SEL[56] BIT_SEL[48] 0.24444f
C549 BIT_SEL[20] BIT_SEL[18] 1.37487f
C550 BIT_SEL[22] BIT_SEL[16] 0.22864f
C551 BIT_SEL[44] BIT_SEL[35] 0.27116f
C552 BIT_SEL[8] BIT_SEL[1] 0.25472f
C553 BIT_SEL[3] BIT_SEL[9] 0.21768f
C554 BIT_SEL[33] BIT_SEL[41] 0.25124f
C555 BIT_SEL[52] BIT_SEL[63] 0.30114f
C556 BIT_SEL[35] BIT_SEL[39] 0.26814f
C557 BIT_SEL[18] BIT_SEL[31] 0.30342f
C558 BIT_SEL[21] BIT_SEL[37] 1.34627f
C559 BIT_SEL[50] BIT_SEL[61] 0.24013f
C560 BIT_SEL[48] BIT_SEL[59] 0.22736f
C561 BIT_SEL[1] BIT_SEL[11] 0.29183f
C562 BIT_SEL[16] BIT_SEL[29] 0.23927f
C563 BIT_SEL[5] BIT_SEL[7] 1.38186f
C564 BIT_SEL[62] BIT_SEL[56] 0.26507f
C565 BIT_SEL[28] BIT_SEL[24] 0.24265f
C566 BIT_SEL[30] BIT_SEL[22] 0.26043f
C567 BIT_SEL[60] BIT_SEL[58] 1.9907f
C568 VDD BIT_SEL[48] 10.3134f
C569 BIT_SEL[26] BIT_SEL[25] 25.7303f
C570 BIT_SEL[58] BIT_SEL[55] 0.24953f
C571 BIT_SEL[60] BIT_SEL[57] 0.27368f
C572 BIT_SEL[30] BIT_SEL[29] 25.7364f
C573 BIT_SEL[56] BIT_SEL[53] 0.22247f
C574 BIT_SEL[32] BIT_SEL[48] 1.35136f
C575 BIT_SEL[24] BIT_SEL[23] 25.7007f
C576 BIT_SEL[28] BIT_SEL[27] 25.7374f
C577 BIT_SEL[0] SENSE 0.0227f
C578 BIT_SEL[62] BIT_SEL[59] 0.26348f
C579 BIT_SEL[22] BIT_SEL[21] 25.7241f
C580 BIT_SEL[55] BIT_SEL[57] 2.1937f
C581 BIT_SEL[53] BIT_SEL[59] 0.27685f
C582 BIT_SEL[23] BIT_SEL[27] 0.28253f
C583 BIT_SEL[21] BIT_SEL[29] 0.26342f
C584 VDD BIT_SEL[62] 0.21883f
C585 BIT_SEL[14] SENSE 0.0227f
C586 BIT_SEL[6] BIT_SEL[22] 1.34627f
C587 BIT_SEL[28] BIT_SEL[0] 0.01882f
C588 BIT_SEL[62] BIT_SEL[32] 0.01882f
C589 VDD BIT_SEL[53] 0.23295f
C590 BIT_SEL[32] BIT_SEL[53] 0.01882f
C591 SENSE OUT[7] 0.05922f
C592 BIT_SEL[0] BIT_SEL[23] 0.01882f
C593 BIT_SEL[33] BIT_SEL[35] 1.14059f
C594 BIT_SEL[1] BIT_SEL[5] 0.30911f
C595 BIT_SEL[46] BIT_SEL[62] 1.34627f
C596 BIT_SEL[13] BIT_SEL[29] 1.34627f
C597 BIT_SEL[4] BIT_SEL[0] 0.27877f
C598 BIT_SEL[26] BIT_SEL[19] 0.25545f
C599 BIT_SEL[58] BIT_SEL[49] 0.27818f
C600 BIT_SEL[24] BIT_SEL[17] 0.25472f
C601 BIT_SEL[36] BIT_SEL[34] 1.37487f
C602 BIT_SEL[38] BIT_SEL[32] 0.22864f
C603 BIT_SEL[60] BIT_SEL[51] 0.27116f
C604 BIT_SEL[19] BIT_SEL[25] 0.21768f
C605 BIT_SEL[17] BIT_SEL[27] 0.29183f
C606 BIT_SEL[32] BIT_SEL[45] 0.23927f
C607 BIT_SEL[51] BIT_SEL[55] 0.26814f
C608 BIT_SEL[0] BIT_SEL[15] 0.28034f
C609 BIT_SEL[37] BIT_SEL[53] 1.34627f
C610 BIT_SEL[34] BIT_SEL[47] 0.30342f
C611 BIT_SEL[49] BIT_SEL[57] 0.25124f
C612 BIT_SEL[46] BIT_SEL[38] 0.26043f
C613 BIT_SEL[14] BIT_SEL[4] 0.2588f
C614 BIT_SEL[10] BIT_SEL[8] 2.44362f
C615 BIT_SEL[12] BIT_SEL[6] 0.22524f
C616 BIT_SEL[44] BIT_SEL[40] 0.24265f
C617 VDD SENSE 4.89915f
C618 BIT_SEL[40] BIT_SEL[39] 25.7007f
C619 BIT_SEL[38] BIT_SEL[37] 25.7241f
C620 BIT_SEL[6] BIT_SEL[7] 25.7222f
C621 BIT_SEL[46] BIT_SEL[45] 25.7364f
C622 BIT_SEL[14] BIT_SEL[15] 28.6814f
C623 BIT_SEL[0] BIT_SEL[17] 0.01882f
C624 BIT_SEL[10] BIT_SEL[11] 25.7092f
C625 BIT_SEL[44] BIT_SEL[43] 25.7374f
C626 BIT_SEL[42] BIT_SEL[41] 25.7303f
C627 BIT_SEL[8] BIT_SEL[9] 25.7235f
C628 BIT_SEL[12] BIT_SEL[13] 25.7382f
C629 BIT_SEL[37] BIT_SEL[45] 0.26342f
C630 BIT_SEL[9] BIT_SEL[11] 2.58494f
C631 BIT_SEL[39] BIT_SEL[43] 0.28253f
C632 BIT_SEL[7] BIT_SEL[13] 0.27378f
C633 BIT_SEL[44] BIT_SEL[16] 0.01882f
C634 BIT_SEL[22] BIT_SEL[38] 1.34627f
C635 BIT_SEL[16] BIT_SEL[39] 0.01882f
C636 BIT_SEL[49] BIT_SEL[51] 1.14059f
C637 BIT_SEL[29] BIT_SEL[45] 1.34627f
C638 BIT_SEL[6] BIT_SEL[1] 0.2966f
C639 BIT_SEL[42] BIT_SEL[35] 0.25545f
C640 BIT_SEL[54] BIT_SEL[48] 0.22864f
C641 BIT_SEL[20] BIT_SEL[16] 0.27877f
C642 BIT_SEL[8] BIT_SEL[3] 0.23548f
C643 BIT_SEL[10] BIT_SEL[5] 0.23973f
C644 BIT_SEL[40] BIT_SEL[33] 0.25472f
C645 BIT_SEL[52] BIT_SEL[50] 1.37487f
C646 VDD BIT_SEL[15] 0.01196f
C647 BIT_SEL[48] BIT_SEL[61] 0.23927f
C648 BIT_SEL[35] BIT_SEL[41] 0.21768f
C649 BIT_SEL[33] BIT_SEL[43] 0.29183f
C650 BIT_SEL[3] BIT_SEL[11] 0.25726f
C651 BIT_SEL[5] BIT_SEL[9] 0.23468f
C652 BIT_SEL[50] BIT_SEL[63] 0.30342f
C653 BIT_SEL[16] BIT_SEL[31] 0.28034f
C654 BIT_SEL[1] BIT_SEL[13] 0.28574f
C655 OUT[0] VSS 0.24364f
C656 COL_PROG_N[0] VSS 0.31996f
C657 OUT[1] VSS 0.24364f
C658 COL_PROG_N[1] VSS 0.26368f
C659 OUT[2] VSS 0.24364f
C660 COL_PROG_N[2] VSS 0.26368f
C661 OUT[3] VSS 0.24364f
C662 COL_PROG_N[3] VSS 0.26368f
C663 OUT[4] VSS 0.24364f
C664 COL_PROG_N[4] VSS 0.26368f
C665 OUT[5] VSS 0.24364f
C666 COL_PROG_N[5] VSS 0.26368f
C667 OUT[6] VSS 0.24364f
C668 COL_PROG_N[6] VSS 0.26368f
C669 BIT_SEL[63] VSS 77.63976f
C670 BIT_SEL[47] VSS 77.67365f
C671 BIT_SEL[31] VSS 77.67365f
C672 BIT_SEL[15] VSS 78.10236f
C673 BIT_SEL[61] VSS 76.1151f
C674 BIT_SEL[45] VSS 76.1583f
C675 BIT_SEL[29] VSS 76.1583f
C676 BIT_SEL[13] VSS 76.4484f
C677 BIT_SEL[59] VSS 75.1795f
C678 BIT_SEL[43] VSS 75.2761f
C679 BIT_SEL[27] VSS 75.2761f
C680 BIT_SEL[11] VSS 75.5839f
C681 BIT_SEL[57] VSS 74.6701f
C682 BIT_SEL[41] VSS 74.7218f
C683 BIT_SEL[25] VSS 74.7218f
C684 BIT_SEL[9] VSS 75.02949f
C685 BIT_SEL[55] VSS 74.37981f
C686 BIT_SEL[39] VSS 74.43552f
C687 BIT_SEL[23] VSS 74.43552f
C688 BIT_SEL[7] VSS 74.75763f
C689 BIT_SEL[53] VSS 73.46686f
C690 BIT_SEL[37] VSS 73.53016f
C691 BIT_SEL[21] VSS 73.53016f
C692 OUT[7] VSS 0.24364f
C693 BIT_SEL[5] VSS 73.82256f
C694 BIT_SEL[51] VSS 72.99814f
C695 BIT_SEL[35] VSS 73.09554f
C696 BIT_SEL[19] VSS 73.09544f
C697 BIT_SEL[3] VSS 73.40794f
C698 BIT_SEL[49] VSS 73.35287f
C699 BIT_SEL[33] VSS 73.53497f
C700 BIT_SEL[17] VSS 73.53497f
C701 BIT_SEL[1] VSS 73.88026f
C702 SENSE VSS 12.642f
C703 PRESET_N VSS 23.65587f
C704 BIT_SEL[48] VSS 70.54855f
C705 BIT_SEL[32] VSS 83.42216f
C706 BIT_SEL[16] VSS 83.42216f
C707 BIT_SEL[0] VSS 83.71227f
C708 BIT_SEL[50] VSS 73.15499f
C709 BIT_SEL[34] VSS 73.27539f
C710 BIT_SEL[18] VSS 73.27539f
C711 BIT_SEL[2] VSS 73.5981f
C712 BIT_SEL[52] VSS 73.74922f
C713 BIT_SEL[36] VSS 73.83221f
C714 BIT_SEL[20] VSS 73.83221f
C715 BIT_SEL[4] VSS 74.22492f
C716 BIT_SEL[54] VSS 74.19282f
C717 BIT_SEL[38] VSS 74.25162f
C718 BIT_SEL[22] VSS 74.25162f
C719 BIT_SEL[6] VSS 74.57222f
C720 BIT_SEL[56] VSS 74.74476f
C721 BIT_SEL[40] VSS 74.83517f
C722 BIT_SEL[24] VSS 74.83517f
C723 BIT_SEL[8] VSS 75.13598f
C724 BIT_SEL[58] VSS 75.03268f
C725 BIT_SEL[42] VSS 75.08308f
C726 BIT_SEL[26] VSS 75.08308f
C727 BIT_SEL[10] VSS 75.46397f
C728 BIT_SEL[60] VSS 75.76613f
C729 BIT_SEL[44] VSS 75.80943f
C730 BIT_SEL[28] VSS 75.80943f
C731 BIT_SEL[12] VSS 76.19472f
C732 BIT_SEL[62] VSS 76.81227f
C733 BIT_SEL[46] VSS 76.85559f
C734 BIT_SEL[30] VSS 76.85559f
C735 BIT_SEL[14] VSS 77.14569f
C736 COL_PROG_N[7] VSS 0.48031f
C737 VDD VSS 0.36167p
C738 a_1340_15066.t0 VSS 4.06398f
C739 a_1340_15066.t1 VSS 2.23602f
C740 a_20810_44412.t0 VSS 4.30649f
C741 a_20810_44412.t1 VSS 1.69351f
C742 a_1340_26048.t0 VSS 4.3173f
C743 a_1340_26048.t1 VSS 1.6827f
C744 a_7830_7189.t0 VSS 4.06398f
C745 a_7830_7189.t1 VSS 2.23602f
C746 a_1340_46574.t0 VSS 4.06398f
C747 a_1340_46574.t1 VSS 2.23602f
C748 a_1340_30820.t0 VSS 4.06398f
C749 a_1340_30820.t1 VSS 2.23602f
C750 a_14320_52657.t0 VSS 4.27849f
C751 a_14320_52657.t1 VSS 1.72151f
C752 a_20810_29555.t0 VSS 4.25498f
C753 a_20810_29555.t1 VSS 1.74502f
C754 a_1340_53922.t0 VSS 4.08932f
C755 a_1340_53922.t1 VSS 1.91068f
C756 a_7738_35589.t0 VSS 1.47655f
C757 a_7738_35589.t1 VSS 4.52345f
C758 a_14320_1152.t0 VSS 4.01916f
C759 a_14320_1152.t1 VSS 1.98084f
C760 a_20810_25520.t0 VSS 4.30261f
C761 a_20810_25520.t1 VSS 1.69739f
C762 a_14320_37432.t0 VSS 4.25498f
C763 a_14320_37432.t1 VSS 1.74502f
C764 a_20718_43466.t0 VSS 1.47655f
C765 a_20718_43466.t1 VSS 4.52345f
C766 a_1248_4081.t0 VSS 4.52345f
C767 a_1248_4081.t1 VSS 1.47655f
C768 a_1340_56291.t0 VSS 4.01916f
C769 a_1340_56291.t1 VSS 1.98084f
C770 a_7830_62696.t0 VSS 2.354f
C771 a_7830_62696.t1 VSS 3.746f
C772 a_14320_26417.t0 VSS 4.34773f
C773 a_14320_26417.t1 VSS 1.65227f
C774 a_20718_11958.t0 VSS 1.47655f
C775 a_20718_11958.t1 VSS 4.52345f
C776 a_1340_16906.t0 VSS 4.01916f
C777 a_1340_16906.t1 VSS 1.98084f
C778 a_1340_53186.t0 VSS 4.25498f
C779 a_1340_53186.t1 VSS 1.74502f
C780 a_14320_29555.t0 VSS 4.25498f
C781 a_14320_29555.t1 VSS 1.74502f
C782 a_14320_9766.t0 VSS 1.69725f
C783 a_14320_9766.t1 VSS 4.30275f
C784 a_1340_47518.t0 VSS 3.68292f
C785 a_1340_47518.t1 VSS 2.41708f
C786 a_1340_42171.t0 VSS 1.6522f
C787 a_1340_42171.t1 VSS 4.3478f
C788 a_1340_54819.t0 VSS 3.74618f
C789 a_1340_54819.t1 VSS 2.35382f
C790 a_20810_36535.t0 VSS 4.30649f
C791 a_20810_36535.t1 VSS 1.69351f
C792 a_1340_40009.t0 VSS 2.23454f
C793 a_1340_40009.t1 VSS 3.86546f
C794 a_14320_25520.t0 VSS 4.30261f
C795 a_14320_25520.t1 VSS 1.69739f
C796 a_1340_38697.t0 VSS 4.06398f
C797 a_1340_38697.t1 VSS 2.23602f
C798 a_1340_10663.t0 VSS 1.6522f
C799 a_1340_10663.t1 VSS 4.3478f
C800 a_14228_43466.t0 VSS 4.52345f
C801 a_14228_43466.t1 VSS 1.47655f
C802 a_7830_32660.t0 VSS 4.01916f
C803 a_7830_32660.t1 VSS 1.98084f
C804 a_20810_1521.t0 VSS 4.20807f
C805 a_20810_1521.t1 VSS 1.79193f
C806 a_7830_24255.t0 VSS 3.86539f
C807 a_7830_24255.t1 VSS 2.23461f
C808 a_1340_16378.t0 VSS 3.86539f
C809 a_1340_16378.t1 VSS 2.23461f
C810 a_14228_11958.t0 VSS 4.52345f
C811 a_14228_11958.t1 VSS 1.47655f
C812 a_1340_53554.t0 VSS 2.33483f
C813 a_1340_53554.t1 VSS 3.66517f
C814 a_20810_33397.t0 VSS 4.30261f
C815 a_20810_33397.t1 VSS 1.69739f
C816 a_1340_34662.t0 VSS 1.39007f
C817 a_1340_34662.t1 VSS 4.60993f
C818 a_7830_55395.t0 VSS 2.41699f
C819 a_7830_55395.t1 VSS 3.68301f
C820 a_14320_56660.t0 VSS 1.79192f
C821 a_14320_56660.t1 VSS 4.20808f
C822 a_14320_38168.t0 VSS 4.08932f
C823 a_14320_38168.t1 VSS 1.91068f
C824 a_7830_7557.t0 VSS 2.354f
C825 a_7830_7557.t1 VSS 3.746f
C826 a_7830_5924.t0 VSS 4.25498f
C827 a_7830_5924.t1 VSS 1.74502f
C828 a_1340_60534.t0 VSS 4.27849f
C829 a_1340_60534.t1 VSS 1.72151f
C830 a_7830_57028.t0 VSS 1.69725f
C831 a_7830_57028.t1 VSS 4.30275f
C832 a_20810_56660.t0 VSS 4.20807f
C833 a_20810_56660.t1 VSS 1.79193f
C834 a_1340_8501.t0 VSS 2.23454f
C835 a_1340_8501.t1 VSS 3.86546f
C836 a_20810_17643.t0 VSS 4.30261f
C837 a_20810_17643.t1 VSS 1.69739f
C838 a_20810_1889.t0 VSS 4.30261f
C839 a_20810_1889.t1 VSS 1.69739f
C840 a_20718_35589.t0 VSS 1.47655f
C841 a_20718_35589.t1 VSS 4.52345f
C842 a_7738_59220.t0 VSS 4.52345f
C843 a_7738_59220.t1 VSS 1.47655f
C844 a_20810_17275.t0 VSS 4.20807f
C845 a_20810_17275.t1 VSS 1.79193f
C846 a_1340_12904.t0 VSS 4.30649f
C847 a_1340_12904.t1 VSS 1.69351f
C848 a_14320_8133.t0 VSS 3.68292f
C849 a_14320_8133.t1 VSS 2.41708f
C850 a_20810_31188.t0 VSS 3.74618f
C851 a_20810_31188.t1 VSS 2.35382f
C852 a_14320_18540.t0 VSS 4.34773f
C853 a_14320_18540.t1 VSS 1.65227f
C854 a_7830_22943.t0 VSS 4.06398f
C855 a_7830_22943.t1 VSS 2.23602f
C856 a_7830_49151.t0 VSS 1.69725f
C857 a_7830_49151.t1 VSS 4.30275f
C858 a_14320_6292.t0 VSS 3.66536f
C859 a_14320_6292.t1 VSS 2.33464f
C860 a_1340_9398.t0 VSS 4.20807f
C861 a_1340_9398.t1 VSS 1.79193f
C862 a_14320_33397.t0 VSS 4.30261f
C863 a_14320_33397.t1 VSS 1.69739f
C864 a_7830_29026.t0 VSS 4.27849f
C865 a_7830_29026.t1 VSS 1.72151f
C866 a_7830_57925.t0 VSS 4.34773f
C867 a_7830_57925.t1 VSS 1.65227f
C868 a_1340_5027.t0 VSS 4.30649f
C869 a_1340_5027.t1 VSS 1.69351f
C870 a_20810_33029.t0 VSS 4.20807f
C871 a_20810_33029.t1 VSS 1.79193f
C872 a_1340_256.t0 VSS 3.68292f
C873 a_1340_256.t1 VSS 2.41708f
C874 a_20810_18540.t0 VSS 4.34773f
C875 a_20810_18540.t1 VSS 1.65227f
C876 a_14320_52289.t0 VSS 1.69351f
C877 a_14320_52289.t1 VSS 4.30649f
C878 a_1340_62328.t0 VSS 4.06398f
C879 a_1340_62328.t1 VSS 2.23602f
C880 a_7830_50416.t0 VSS 1.39007f
C881 a_7830_50416.t1 VSS 4.60993f
C882 a_7830_40537.t0 VSS 4.01916f
C883 a_7830_40537.t1 VSS 1.98084f
C884 a_1340_34294.t0 VSS 1.6522f
C885 a_1340_34294.t1 VSS 4.3478f
C886 a_1340_1152.t0 VSS 4.01916f
C887 a_1340_1152.t1 VSS 1.98084f
C888 a_7830_24783.t0 VSS 4.01916f
C889 a_7830_24783.t1 VSS 1.98084f
C890 a_20810_28658.t0 VSS 4.30649f
C891 a_20810_28658.t1 VSS 1.69351f
C892 a_20718_27712.t0 VSS 1.47655f
C893 a_20718_27712.t1 VSS 4.52345f
C894 a_20810_624.t0 VSS 2.23454f
C895 a_20810_624.t1 VSS 3.86546f
C896 a_14320_17643.t0 VSS 4.30261f
C897 a_14320_17643.t1 VSS 1.69739f
C898 a_14320_7189.t0 VSS 4.06398f
C899 a_14320_7189.t1 VSS 2.23602f
C900 a_20810_256.t0 VSS 2.41699f
C901 a_20810_256.t1 VSS 3.68301f
C902 a_14228_35589.t0 VSS 4.52345f
C903 a_14228_35589.t1 VSS 1.47655f
C904 a_14320_17275.t0 VSS 1.79192f
C905 a_14320_17275.t1 VSS 4.20808f
C906 a_1340_45309.t0 VSS 4.25498f
C907 a_1340_45309.t1 VSS 1.74502f
C908 a_20810_2417.t0 VSS 4.3173f
C909 a_20810_2417.t1 VSS 1.6827f
C910 a_7830_15066.t0 VSS 4.06398f
C911 a_7830_15066.t1 VSS 2.23602f
C912 a_14320_31764.t0 VSS 2.41699f
C913 a_14320_31764.t1 VSS 3.68301f
C914 a_7830_33029.t0 VSS 4.20807f
C915 a_7830_33029.t1 VSS 1.79193f
C916 a_1340_58293.t0 VSS 1.39007f
C917 a_1340_58293.t1 VSS 4.60993f
C918 a_20810_62696.t0 VSS 3.74618f
C919 a_20810_62696.t1 VSS 2.35382f
C920 a_14228_19835.t0 VSS 4.52345f
C921 a_14228_19835.t1 VSS 1.47655f
C922 a_7830_32132.t0 VSS 3.86539f
C923 a_7830_32132.t1 VSS 2.23461f
C924 a_1340_57556.t0 VSS 4.3173f
C925 a_1340_57556.t1 VSS 1.6827f
C926 a_7830_17275.t0 VSS 1.79192f
C927 a_7830_17275.t1 VSS 4.20808f
C928 a_14320_31188.t0 VSS 2.354f
C929 a_14320_31188.t1 VSS 3.746f
C930 a_14320_16010.t0 VSS 2.41699f
C931 a_14320_16010.t1 VSS 3.68301f
C932 a_7830_16378.t0 VSS 3.86539f
C933 a_7830_16378.t1 VSS 2.23461f
C934 a_1340_21149.t0 VSS 4.27849f
C935 a_1340_21149.t1 VSS 1.72151f
C936 a_1340_13801.t0 VSS 4.25498f
C937 a_1340_13801.t1 VSS 1.74502f
C938 a_7830_3154.t0 VSS 1.39007f
C939 a_7830_3154.t1 VSS 4.60993f
C940 a_14320_3154.t0 VSS 4.60993f
C941 a_14320_3154.t1 VSS 1.39007f
C942 a_14320_37800.t0 VSS 3.66536f
C943 a_14320_37800.t1 VSS 2.33464f
C944 a_7830_47518.t0 VSS 2.41699f
C945 a_7830_47518.t1 VSS 3.68301f
C946 a_1340_46942.t0 VSS 2.354f
C947 a_1340_46942.t1 VSS 3.746f
C948 a_7830_26048.t0 VSS 4.3173f
C949 a_7830_26048.t1 VSS 1.6827f
C950 a_1340_26417.t0 VSS 1.6522f
C951 a_1340_26417.t1 VSS 4.3478f
C952 a_7830_61799.t0 VSS 4.08932f
C953 a_7830_61799.t1 VSS 1.91068f
C954 a_7830_46574.t0 VSS 4.06398f
C955 a_7830_46574.t1 VSS 2.23602f
C956 a_7830_56291.t0 VSS 4.01916f
C957 a_7830_56291.t1 VSS 1.98084f
C958 a_14320_33029.t0 VSS 1.79192f
C959 a_14320_33029.t1 VSS 4.20808f
C960 a_14320_62696.t0 VSS 2.354f
C961 a_14320_62696.t1 VSS 3.746f
C962 a_7830_30820.t0 VSS 4.06398f
C963 a_7830_30820.t1 VSS 2.23602f
C964 a_1340_48414.t0 VSS 1.98079f
C965 a_1340_48414.t1 VSS 4.01921f
C966 a_1340_15434.t0 VSS 3.74618f
C967 a_1340_15434.t1 VSS 2.35382f
C968 a_7830_9029.t0 VSS 4.01916f
C969 a_7830_9029.t1 VSS 1.98084f
C970 a_1340_36903.t0 VSS 4.27849f
C971 a_1340_36903.t1 VSS 1.72151f
C972 COL_PROG_N[6].t1 VSS 1.10931f
C973 COL_PROG_N[6].n0 VSS 0.38563f
C974 COL_PROG_N[6].t3 VSS 1.10931f
C975 COL_PROG_N[6].n1 VSS 0.39369f
C976 COL_PROG_N[6].t0 VSS 1.10931f
C977 COL_PROG_N[6].n2 VSS 0.77937f
C978 COL_PROG_N[6].t2 VSS 1.10971f
C979 a_20810_5027.t0 VSS 4.30649f
C980 a_20810_5027.t1 VSS 1.69351f
C981 a_14228_27712.t0 VSS 4.52345f
C982 a_14228_27712.t1 VSS 1.47655f
C983 a_1340_20781.t0 VSS 4.30649f
C984 a_1340_20781.t1 VSS 1.69351f
C985 a_7830_42171.t0 VSS 4.34773f
C986 a_7830_42171.t1 VSS 1.65227f
C987 COL_PROG_N[2].t1 VSS 1.10931f
C988 COL_PROG_N[2].n0 VSS 0.38563f
C989 COL_PROG_N[2].t3 VSS 1.10931f
C990 COL_PROG_N[2].n1 VSS 0.39369f
C991 COL_PROG_N[2].t0 VSS 1.10931f
C992 COL_PROG_N[2].n2 VSS 0.77937f
C993 COL_PROG_N[2].t2 VSS 1.10971f
C994 a_7830_53922.t0 VSS 4.08932f
C995 a_7830_53922.t1 VSS 1.91068f
C996 a_14320_2786.t0 VSS 4.34773f
C997 a_14320_2786.t1 VSS 1.65227f
C998 a_7830_624.t0 VSS 3.86539f
C999 a_7830_624.t1 VSS 2.23461f
C1000 a_1340_60166.t0 VSS 4.30649f
C1001 a_1340_60166.t1 VSS 1.69351f
C1002 a_20810_23311.t0 VSS 3.74618f
C1003 a_20810_23311.t1 VSS 2.35382f
C1004 a_20810_57028.t0 VSS 4.30261f
C1005 a_20810_57028.t1 VSS 1.69739f
C1006 a_7830_11031.t0 VSS 4.60993f
C1007 a_7830_11031.t1 VSS 1.39007f
C1008 a_20810_23887.t0 VSS 2.41699f
C1009 a_20810_23887.t1 VSS 3.68301f
C1010 a_7830_10663.t0 VSS 4.34773f
C1011 a_7830_10663.t1 VSS 1.65227f
C1012 a_1340_10294.t0 VSS 4.3173f
C1013 a_1340_10294.t1 VSS 1.6827f
C1014 a_1340_52657.t0 VSS 4.27849f
C1015 a_1340_52657.t1 VSS 1.72151f
C1016 a_14320_44780.t0 VSS 4.27849f
C1017 a_14320_44780.t1 VSS 1.72151f
C1018 a_20718_59220.t0 VSS 1.47655f
C1019 a_20718_59220.t1 VSS 4.52345f
C1020 a_20810_9029.t0 VSS 4.01916f
C1021 a_20810_9029.t1 VSS 1.98084f
C1022 a_7830_28658.t0 VSS 1.69351f
C1023 a_7830_28658.t1 VSS 4.30649f
C1024 a_14320_29026.t0 VSS 4.27849f
C1025 a_14320_29026.t1 VSS 1.72151f
C1026 a_7830_22046.t0 VSS 3.66536f
C1027 a_7830_22046.t1 VSS 2.33464f
C1028 a_14320_57925.t0 VSS 1.6522f
C1029 a_14320_57925.t1 VSS 4.3478f
C1030 a_20718_4081.t0 VSS 1.47655f
C1031 a_20718_4081.t1 VSS 4.52345f
C1032 a_20810_2786.t0 VSS 4.34773f
C1033 a_20810_2786.t1 VSS 1.65227f
C1034 a_1340_46045.t0 VSS 4.08932f
C1035 a_1340_46045.t1 VSS 1.91068f
C1036 a_7830_62328.t0 VSS 4.06398f
C1037 a_7830_62328.t1 VSS 2.23602f
C1038 a_7830_2417.t0 VSS 4.3173f
C1039 a_7830_2417.t1 VSS 1.6827f
C1040 BIT_SEL[31].t4 VSS 3.1518f
C1041 BIT_SEL[31].n0 VSS 5.61038f
C1042 BIT_SEL[31].t2 VSS 3.1518f
C1043 BIT_SEL[31].n1 VSS 5.61038f
C1044 BIT_SEL[31].t5 VSS 3.1518f
C1045 BIT_SEL[31].n2 VSS 5.61038f
C1046 BIT_SEL[31].t0 VSS 3.1518f
C1047 BIT_SEL[31].n3 VSS 5.61038f
C1048 BIT_SEL[31].t1 VSS 3.1518f
C1049 BIT_SEL[31].n4 VSS 5.61038f
C1050 BIT_SEL[31].t3 VSS 3.1518f
C1051 BIT_SEL[31].n5 VSS 5.61038f
C1052 BIT_SEL[31].t7 VSS 3.1518f
C1053 BIT_SEL[31].n6 VSS 5.61038f
C1054 BIT_SEL[31].t6 VSS 3.38636f
C1055 a_1340_30291.t0 VSS 4.08932f
C1056 a_1340_30291.t1 VSS 1.91068f
C1057 a_1340_41802.t0 VSS 4.3173f
C1058 a_1340_41802.t1 VSS 1.6827f
C1059 a_1340_18540.t0 VSS 1.6522f
C1060 a_1340_18540.t1 VSS 4.3478f
C1061 a_20810_44780.t0 VSS 1.7215f
C1062 a_20810_44780.t1 VSS 4.2785f
C1063 a_14320_55763.t0 VSS 3.86539f
C1064 a_14320_55763.t1 VSS 2.23461f
C1065 a_7830_16906.t0 VSS 4.01916f
C1066 a_7830_16906.t1 VSS 1.98084f
C1067 a_1340_14537.t0 VSS 4.08932f
C1068 a_1340_14537.t1 VSS 1.91068f
C1069 a_7830_53554.t0 VSS 3.66536f
C1070 a_7830_53554.t1 VSS 2.33464f
C1071 a_20810_29923.t0 VSS 2.33483f
C1072 a_20810_29923.t1 VSS 3.66517f
C1073 a_20810_29026.t0 VSS 1.7215f
C1074 a_20810_29026.t1 VSS 4.2785f
C1075 a_14320_55395.t0 VSS 2.41699f
C1076 a_14320_55395.t1 VSS 3.68301f
C1077 a_20810_57925.t0 VSS 4.34773f
C1078 a_20810_57925.t1 VSS 1.65227f
C1079 a_7830_53186.t0 VSS 4.25498f
C1080 a_7830_53186.t1 VSS 1.74502f
C1081 a_14320_48783.t0 VSS 1.79192f
C1082 a_14320_48783.t1 VSS 4.20808f
C1083 a_1340_44412.t0 VSS 4.30649f
C1084 a_1340_44412.t1 VSS 1.69351f
C1085 a_7830_1889.t0 VSS 1.69725f
C1086 a_7830_1889.t1 VSS 4.30275f
C1087 a_7830_49679.t0 VSS 4.3173f
C1088 a_7830_49679.t1 VSS 1.6827f
C1089 a_20810_50416.t0 VSS 4.60993f
C1090 a_20810_50416.t1 VSS 1.39007f
C1091 a_1340_37432.t0 VSS 4.25498f
C1092 a_1340_37432.t1 VSS 1.74502f
C1093 a_20810_40537.t0 VSS 4.01916f
C1094 a_20810_40537.t1 VSS 1.98084f
C1095 a_14320_23887.t0 VSS 2.41699f
C1096 a_14320_23887.t1 VSS 3.68301f
C1097 a_20810_46942.t0 VSS 3.74618f
C1098 a_20810_46942.t1 VSS 2.35382f
C1099 a_20810_24783.t0 VSS 4.01916f
C1100 a_20810_24783.t1 VSS 1.98084f
C1101 a_1340_21678.t0 VSS 4.25498f
C1102 a_1340_21678.t1 VSS 1.74502f
C1103 a_14320_23311.t0 VSS 2.354f
C1104 a_14320_23311.t1 VSS 3.746f
C1105 a_1340_50416.t0 VSS 1.39007f
C1106 a_1340_50416.t1 VSS 4.60993f
C1107 a_14320_57028.t0 VSS 4.30261f
C1108 a_14320_57028.t1 VSS 1.69739f
C1109 a_14320_42539.t0 VSS 4.60993f
C1110 a_14320_42539.t1 VSS 1.39007f
C1111 a_7830_54819.t0 VSS 2.354f
C1112 a_7830_54819.t1 VSS 3.746f
C1113 BIT_SEL[30].t2 VSS 4.1517f
C1114 BIT_SEL[30].n0 VSS 7.36453f
C1115 BIT_SEL[30].t4 VSS 4.1517f
C1116 BIT_SEL[30].n1 VSS 7.36453f
C1117 BIT_SEL[30].t6 VSS 4.1517f
C1118 BIT_SEL[30].n2 VSS 7.36453f
C1119 BIT_SEL[30].t1 VSS 4.1517f
C1120 BIT_SEL[30].n3 VSS 7.36453f
C1121 BIT_SEL[30].t3 VSS 4.1517f
C1122 BIT_SEL[30].n4 VSS 7.36453f
C1123 BIT_SEL[30].t0 VSS 4.1517f
C1124 BIT_SEL[30].n5 VSS 7.36453f
C1125 BIT_SEL[30].t5 VSS 4.45988f
C1126 BIT_SEL[30].t7 VSS 4.1517f
C1127 BIT_SEL[30].n6 VSS 7.36453f
C1128 a_20810_61063.t0 VSS 4.25498f
C1129 a_20810_61063.t1 VSS 1.74502f
C1130 a_7830_40009.t0 VSS 3.86539f
C1131 a_7830_40009.t1 VSS 2.23461f
C1132 a_7830_33925.t0 VSS 4.3173f
C1133 a_7830_33925.t1 VSS 1.6827f
C1134 a_20810_48783.t0 VSS 4.20807f
C1135 a_20810_48783.t1 VSS 1.79193f
C1136 a_1340_6292.t0 VSS 3.66536f
C1137 a_1340_6292.t1 VSS 2.33464f
C1138 BIT_SEL[8].t0 VSS 4.14071f
C1139 BIT_SEL[8].n0 VSS 7.18434f
C1140 BIT_SEL[8].t4 VSS 4.14071f
C1141 BIT_SEL[8].n1 VSS 7.18434f
C1142 BIT_SEL[8].t6 VSS 4.14071f
C1143 BIT_SEL[8].n2 VSS 7.18434f
C1144 BIT_SEL[8].t7 VSS 4.14071f
C1145 BIT_SEL[8].n3 VSS 7.18434f
C1146 BIT_SEL[8].t1 VSS 4.14071f
C1147 BIT_SEL[8].n4 VSS 7.18434f
C1148 BIT_SEL[8].t2 VSS 4.14071f
C1149 BIT_SEL[8].n5 VSS 7.18434f
C1150 BIT_SEL[8].t5 VSS 4.14071f
C1151 BIT_SEL[8].n6 VSS 7.18434f
C1152 BIT_SEL[8].t3 VSS 4.31483f
C1153 a_1340_18908.t0 VSS 1.39007f
C1154 a_1340_18908.t1 VSS 4.60993f
C1155 a_14320_26785.t0 VSS 4.60993f
C1156 a_14320_26785.t1 VSS 1.39007f
C1157 a_20810_15434.t0 VSS 3.74618f
C1158 a_20810_15434.t1 VSS 2.35382f
C1159 a_1340_39065.t0 VSS 3.74618f
C1160 a_1340_39065.t1 VSS 2.35382f
C1161 a_14228_59220.t0 VSS 4.52345f
C1162 a_14228_59220.t1 VSS 1.47655f
C1163 a_7830_18171.t0 VSS 4.3173f
C1164 a_7830_18171.t1 VSS 1.6827f
C1165 a_20810_30291.t0 VSS 4.08932f
C1166 a_20810_30291.t1 VSS 1.91068f
C1167 a_20810_15066.t0 VSS 4.06398f
C1168 a_20810_15066.t1 VSS 2.23602f
C1169 a_20810_6660.t0 VSS 1.91084f
C1170 a_20810_6660.t1 VSS 4.08916f
C1171 a_7830_38697.t0 VSS 4.06398f
C1172 a_7830_38697.t1 VSS 2.23602f
C1173 BIT_SEL[28].t5 VSS 4.12331f
C1174 BIT_SEL[28].n0 VSS 7.26213f
C1175 BIT_SEL[28].t6 VSS 4.12331f
C1176 BIT_SEL[28].n1 VSS 7.26213f
C1177 BIT_SEL[28].t2 VSS 4.12331f
C1178 BIT_SEL[28].n2 VSS 7.26213f
C1179 BIT_SEL[28].t0 VSS 4.12331f
C1180 BIT_SEL[28].n3 VSS 7.26213f
C1181 BIT_SEL[28].t3 VSS 4.12331f
C1182 BIT_SEL[28].n4 VSS 7.26213f
C1183 BIT_SEL[28].t1 VSS 4.12331f
C1184 BIT_SEL[28].n5 VSS 7.26213f
C1185 BIT_SEL[28].t4 VSS 4.3879f
C1186 BIT_SEL[28].t7 VSS 4.12331f
C1187 BIT_SEL[28].n6 VSS 7.26213f
C1188 a_7830_56660.t0 VSS 1.79192f
C1189 a_7830_56660.t1 VSS 4.20808f
C1190 a_1340_41274.t0 VSS 4.30261f
C1191 a_1340_41274.t1 VSS 1.69739f
C1192 a_7738_51343.t0 VSS 1.47655f
C1193 a_7738_51343.t1 VSS 4.52345f
C1194 a_7830_55763.t0 VSS 3.86539f
C1195 a_7830_55763.t1 VSS 2.23461f
C1196 a_1340_29555.t0 VSS 4.25498f
C1197 a_1340_29555.t1 VSS 1.74502f
C1198 COL_PROG_N[7].t1 VSS 1.09082f
C1199 COL_PROG_N[7].n0 VSS 0.3792f
C1200 COL_PROG_N[7].t3 VSS 1.09082f
C1201 COL_PROG_N[7].n1 VSS 0.38712f
C1202 COL_PROG_N[7].t0 VSS 1.09082f
C1203 COL_PROG_N[7].n2 VSS 0.76638f
C1204 COL_PROG_N[7].t2 VSS 1.09122f
C1205 a_14320_32660.t0 VSS 1.98079f
C1206 a_14320_32660.t1 VSS 4.01921f
C1207 a_20810_41802.t0 VSS 1.6826f
C1208 a_20810_41802.t1 VSS 4.3174f
C1209 a_20810_47886.t0 VSS 3.86539f
C1210 a_20810_47886.t1 VSS 2.23461f
C1211 a_14320_5395.t0 VSS 4.27849f
C1212 a_14320_5395.t1 VSS 1.72151f
C1213 a_14320_624.t0 VSS 2.23454f
C1214 a_14320_624.t1 VSS 3.86546f
C1215 a_20810_1152.t0 VSS 4.01916f
C1216 a_20810_1152.t1 VSS 1.98084f
C1217 a_7830_6292.t0 VSS 2.33483f
C1218 a_7830_6292.t1 VSS 3.66517f
C1219 a_1340_9766.t0 VSS 4.30261f
C1220 a_1340_9766.t1 VSS 1.69739f
C1221 COL_PROG_N[5].t1 VSS 1.10931f
C1222 COL_PROG_N[5].n0 VSS 0.38563f
C1223 COL_PROG_N[5].t3 VSS 1.10931f
C1224 COL_PROG_N[5].n1 VSS 0.39369f
C1225 COL_PROG_N[5].t0 VSS 1.10931f
C1226 COL_PROG_N[5].n2 VSS 0.77937f
C1227 COL_PROG_N[5].t2 VSS 1.10971f
C1228 a_20810_47518.t0 VSS 3.68292f
C1229 a_20810_47518.t1 VSS 2.41708f
C1230 a_14320_5924.t0 VSS 4.25498f
C1231 a_14320_5924.t1 VSS 1.74502f
C1232 a_20810_26048.t0 VSS 4.3173f
C1233 a_20810_26048.t1 VSS 1.6827f
C1234 a_20810_61799.t0 VSS 4.08932f
C1235 a_20810_61799.t1 VSS 1.91068f
C1236 a_7830_13272.t0 VSS 4.27849f
C1237 a_7830_13272.t1 VSS 1.72151f
C1238 a_14320_29923.t0 VSS 3.66536f
C1239 a_14320_29923.t1 VSS 2.33464f
C1240 a_1340_39641.t0 VSS 2.41699f
C1241 a_1340_39641.t1 VSS 3.68301f
C1242 a_20810_46574.t0 VSS 4.06398f
C1243 a_20810_46574.t1 VSS 2.23602f
C1244 a_1340_7189.t0 VSS 4.06398f
C1245 a_1340_7189.t1 VSS 2.23602f
C1246 COL_PROG_N[3].t1 VSS 1.10931f
C1247 COL_PROG_N[3].n0 VSS 0.38563f
C1248 COL_PROG_N[3].t3 VSS 1.10931f
C1249 COL_PROG_N[3].n1 VSS 0.39369f
C1250 COL_PROG_N[3].t0 VSS 1.10931f
C1251 COL_PROG_N[3].n2 VSS 0.77937f
C1252 COL_PROG_N[3].t2 VSS 1.10971f
C1253 a_7830_34662.t0 VSS 4.60993f
C1254 a_7830_34662.t1 VSS 1.39007f
C1255 a_20810_10294.t0 VSS 4.3173f
C1256 a_20810_10294.t1 VSS 1.6827f
C1257 a_7738_4081.t0 VSS 1.47655f
C1258 a_7738_4081.t1 VSS 4.52345f
C1259 a_7830_34294.t0 VSS 4.34773f
C1260 a_7830_34294.t1 VSS 1.65227f
C1261 a_20810_30820.t0 VSS 4.06398f
C1262 a_20810_30820.t1 VSS 2.23602f
C1263 a_7830_50048.t0 VSS 4.34773f
C1264 a_7830_50048.t1 VSS 1.65227f
C1265 a_7830_2786.t0 VSS 4.34773f
C1266 a_7830_2786.t1 VSS 1.65227f
C1267 a_1340_25520.t0 VSS 4.30261f
C1268 a_1340_25520.t1 VSS 1.69739f
C1269 a_14320_50416.t0 VSS 4.60993f
C1270 a_14320_50416.t1 VSS 1.39007f
C1271 a_1340_54451.t0 VSS 2.2362f
C1272 a_1340_54451.t1 VSS 4.0638f
C1273 a_1340_8133.t0 VSS 3.68292f
C1274 a_1340_8133.t1 VSS 2.41708f
C1275 a_20810_31764.t0 VSS 2.41699f
C1276 a_20810_31764.t1 VSS 3.68301f
C1277 a_20810_32660.t0 VSS 4.01916f
C1278 a_20810_32660.t1 VSS 1.98084f
C1279 a_14320_40537.t0 VSS 4.01916f
C1280 a_14320_40537.t1 VSS 1.98084f
C1281 a_1248_43466.t0 VSS 1.47655f
C1282 a_1248_43466.t1 VSS 4.52345f
C1283 a_14320_6660.t0 VSS 1.91084f
C1284 a_14320_6660.t1 VSS 4.08916f
C1285 a_20810_24255.t0 VSS 2.23454f
C1286 a_20810_24255.t1 VSS 3.86546f
C1287 a_14320_46942.t0 VSS 2.354f
C1288 a_14320_46942.t1 VSS 3.746f
C1289 a_14320_24783.t0 VSS 4.01916f
C1290 a_14320_24783.t1 VSS 1.98084f
C1291 a_20810_16010.t0 VSS 2.41699f
C1292 a_20810_16010.t1 VSS 3.68301f
C1293 COL_PROG_N[1].t2 VSS 1.10931f
C1294 COL_PROG_N[1].n0 VSS 0.38563f
C1295 COL_PROG_N[1].t0 VSS 1.10931f
C1296 COL_PROG_N[1].n1 VSS 0.39369f
C1297 COL_PROG_N[1].t3 VSS 1.10931f
C1298 COL_PROG_N[1].n2 VSS 0.77937f
C1299 COL_PROG_N[1].t1 VSS 1.10971f
C1300 a_7830_36535.t0 VSS 1.69351f
C1301 a_7830_36535.t1 VSS 4.30649f
C1302 a_14320_36903.t0 VSS 1.7215f
C1303 a_14320_36903.t1 VSS 4.2785f
C1304 a_1340_3154.t0 VSS 1.39007f
C1305 a_1340_3154.t1 VSS 4.60993f
C1306 BIT_SEL[1].t6 VSS 4.07792f
C1307 BIT_SEL[1].n0 VSS 6.88058f
C1308 BIT_SEL[1].t1 VSS 4.07792f
C1309 BIT_SEL[1].n1 VSS 6.88058f
C1310 BIT_SEL[1].t2 VSS 4.07792f
C1311 BIT_SEL[1].n2 VSS 6.88058f
C1312 BIT_SEL[1].t5 VSS 4.07792f
C1313 BIT_SEL[1].n3 VSS 6.88058f
C1314 BIT_SEL[1].t3 VSS 4.07792f
C1315 BIT_SEL[1].n4 VSS 6.88058f
C1316 BIT_SEL[1].t7 VSS 4.07792f
C1317 BIT_SEL[1].n5 VSS 6.88058f
C1318 BIT_SEL[1].t4 VSS 4.07792f
C1319 BIT_SEL[1].n6 VSS 6.88058f
C1320 BIT_SEL[1].t0 VSS 4.12246f
C1321 a_20810_5395.t0 VSS 1.7215f
C1322 a_20810_5395.t1 VSS 4.2785f
C1323 a_14320_61063.t0 VSS 4.25498f
C1324 a_14320_61063.t1 VSS 1.74502f
C1325 a_1248_11958.t0 VSS 1.47655f
C1326 a_1248_11958.t1 VSS 4.52345f
C1327 a_20810_8501.t0 VSS 2.23454f
C1328 a_20810_8501.t1 VSS 3.86546f
C1329 a_20810_42171.t0 VSS 4.34773f
C1330 a_20810_42171.t1 VSS 1.65227f
C1331 a_14320_21149.t0 VSS 4.27849f
C1332 a_14320_21149.t1 VSS 1.72151f
C1333 a_14320_57556.t0 VSS 4.3173f
C1334 a_14320_57556.t1 VSS 1.6827f
C1335 a_14320_15434.t0 VSS 2.354f
C1336 a_14320_15434.t1 VSS 3.746f
C1337 a_20810_53922.t0 VSS 4.08932f
C1338 a_20810_53922.t1 VSS 1.91068f
C1339 a_14320_256.t0 VSS 2.41699f
C1340 a_14320_256.t1 VSS 3.68301f
C1341 a_1340_45677.t0 VSS 2.33483f
C1342 a_1340_45677.t1 VSS 3.66517f
C1343 a_7830_46045.t0 VSS 4.08932f
C1344 a_7830_46045.t1 VSS 1.91068f
C1345 a_14320_30291.t0 VSS 4.08932f
C1346 a_14320_30291.t1 VSS 1.91068f
C1347 a_1340_56660.t0 VSS 4.20807f
C1348 a_1340_56660.t1 VSS 1.79193f
C1349 a_14320_15066.t0 VSS 2.2362f
C1350 a_14320_15066.t1 VSS 4.0638f
C1351 a_20810_11031.t0 VSS 1.39007f
C1352 a_20810_11031.t1 VSS 4.60993f
C1353 a_1340_38168.t0 VSS 4.08932f
C1354 a_1340_38168.t1 VSS 1.91068f
C1355 a_1340_29923.t0 VSS 3.66536f
C1356 a_1340_29923.t1 VSS 2.33464f
C1357 a_7830_12904.t0 VSS 1.69351f
C1358 a_7830_12904.t1 VSS 4.30649f
C1359 a_7830_30291.t0 VSS 1.91084f
C1360 a_7830_30291.t1 VSS 4.08916f
C1361 a_20810_10663.t0 VSS 1.6522f
C1362 a_20810_10663.t1 VSS 4.3478f
C1363 a_1340_22414.t0 VSS 4.08932f
C1364 a_1340_22414.t1 VSS 1.91068f
C1365 a_7830_256.t0 VSS 2.41699f
C1366 a_7830_256.t1 VSS 3.68301f
C1367 a_20810_22414.t0 VSS 4.08932f
C1368 a_20810_22414.t1 VSS 1.91068f
C1369 a_7830_61431.t0 VSS 3.66536f
C1370 a_7830_61431.t1 VSS 2.33464f
C1371 a_20810_37800.t0 VSS 2.33483f
C1372 a_20810_37800.t1 VSS 3.66517f
C1373 a_1340_49679.t0 VSS 1.6826f
C1374 a_1340_49679.t1 VSS 4.3174f
C1375 a_7830_60534.t0 VSS 4.27849f
C1376 a_7830_60534.t1 VSS 1.72151f
C1377 a_1340_14169.t0 VSS 3.66536f
C1378 a_1340_14169.t1 VSS 2.33464f
C1379 a_14320_41802.t0 VSS 1.6826f
C1380 a_14320_41802.t1 VSS 4.3174f
C1381 a_14320_47886.t0 VSS 3.86539f
C1382 a_14320_47886.t1 VSS 2.23461f
C1383 a_7830_14537.t0 VSS 1.91084f
C1384 a_7830_14537.t1 VSS 4.08916f
C1385 BIT_SEL[41].t3 VSS 4.14534f
C1386 BIT_SEL[41].n0 VSS 7.22001f
C1387 BIT_SEL[41].t5 VSS 4.14534f
C1388 BIT_SEL[41].n1 VSS 7.22001f
C1389 BIT_SEL[41].t1 VSS 4.14534f
C1390 BIT_SEL[41].n2 VSS 7.22001f
C1391 BIT_SEL[41].t7 VSS 4.14534f
C1392 BIT_SEL[41].n3 VSS 7.22001f
C1393 BIT_SEL[41].t2 VSS 4.14534f
C1394 BIT_SEL[41].n4 VSS 7.22001f
C1395 BIT_SEL[41].t4 VSS 4.14534f
C1396 BIT_SEL[41].n5 VSS 7.22001f
C1397 BIT_SEL[41].t6 VSS 4.14534f
C1398 BIT_SEL[41].n6 VSS 7.22001f
C1399 BIT_SEL[41].t0 VSS 4.32038f
C1400 a_20810_22046.t0 VSS 2.33483f
C1401 a_20810_22046.t1 VSS 3.66517f
C1402 a_20810_9766.t0 VSS 4.30261f
C1403 a_20810_9766.t1 VSS 1.69739f
C1404 a_14320_26048.t0 VSS 1.6826f
C1405 a_14320_26048.t1 VSS 4.3174f
C1406 a_7830_46942.t0 VSS 3.74618f
C1407 a_7830_46942.t1 VSS 2.35382f
C1408 a_20810_48414.t0 VSS 4.01916f
C1409 a_20810_48414.t1 VSS 1.98084f
C1410 a_7830_45309.t0 VSS 4.25498f
C1411 a_7830_45309.t1 VSS 1.74502f
C1412 a_14320_61799.t0 VSS 1.91084f
C1413 a_14320_61799.t1 VSS 4.08916f
C1414 a_14320_46574.t0 VSS 2.2362f
C1415 a_14320_46574.t1 VSS 4.0638f
C1416 a_1248_51343.t0 VSS 4.52345f
C1417 a_1248_51343.t1 VSS 1.47655f
C1418 a_7830_31188.t0 VSS 3.74618f
C1419 a_7830_31188.t1 VSS 2.35382f
C1420 a_1340_36535.t0 VSS 4.30649f
C1421 a_1340_36535.t1 VSS 1.69351f
C1422 a_1340_2417.t0 VSS 4.3173f
C1423 a_1340_2417.t1 VSS 1.6827f
C1424 a_1340_57925.t0 VSS 1.6522f
C1425 a_1340_57925.t1 VSS 4.3478f
C1426 a_14320_10294.t0 VSS 1.6826f
C1427 a_14320_10294.t1 VSS 4.3174f
C1428 a_20810_39641.t0 VSS 3.68292f
C1429 a_20810_39641.t1 VSS 2.41708f
C1430 a_14320_30820.t0 VSS 4.06398f
C1431 a_14320_30820.t1 VSS 2.23602f
C1432 a_7830_48414.t0 VSS 4.01916f
C1433 a_7830_48414.t1 VSS 1.98084f
C1434 a_1340_47886.t0 VSS 2.23454f
C1435 a_1340_47886.t1 VSS 3.86546f
C1436 a_7830_15434.t0 VSS 3.74618f
C1437 a_7830_15434.t1 VSS 2.35382f
C1438 a_20810_39065.t0 VSS 3.74618f
C1439 a_20810_39065.t1 VSS 2.35382f
C1440 a_20810_16906.t0 VSS 4.01916f
C1441 a_20810_16906.t1 VSS 1.98084f
C1442 BIT_SEL[59].t0 VSS 4.11768f
C1443 BIT_SEL[59].n0 VSS 7.22573f
C1444 BIT_SEL[59].t3 VSS 4.11768f
C1445 BIT_SEL[59].n1 VSS 7.22573f
C1446 BIT_SEL[59].t6 VSS 4.11768f
C1447 BIT_SEL[59].n2 VSS 7.22573f
C1448 BIT_SEL[59].t4 VSS 4.11768f
C1449 BIT_SEL[59].n3 VSS 7.22573f
C1450 BIT_SEL[59].t1 VSS 4.11768f
C1451 BIT_SEL[59].n4 VSS 7.22573f
C1452 BIT_SEL[59].t5 VSS 4.11768f
C1453 BIT_SEL[59].n5 VSS 7.22573f
C1454 BIT_SEL[59].t7 VSS 4.11768f
C1455 BIT_SEL[59].n6 VSS 7.22573f
C1456 BIT_SEL[59].t2 VSS 4.3277f
C1457 a_20810_22943.t0 VSS 4.06398f
C1458 a_20810_22943.t1 VSS 2.23602f
C1459 a_7830_13801.t0 VSS 1.745f
C1460 a_7830_13801.t1 VSS 4.255f
C1461 a_20810_53554.t0 VSS 2.33483f
C1462 a_20810_53554.t1 VSS 3.66517f
C1463 a_7830_1152.t0 VSS 4.01916f
C1464 a_7830_1152.t1 VSS 1.98084f
C1465 BIT_SEL[27].t1 VSS 4.11768f
C1466 BIT_SEL[27].n0 VSS 7.22573f
C1467 BIT_SEL[27].t4 VSS 4.11768f
C1468 BIT_SEL[27].n1 VSS 7.22573f
C1469 BIT_SEL[27].t7 VSS 4.11768f
C1470 BIT_SEL[27].n2 VSS 7.22573f
C1471 BIT_SEL[27].t5 VSS 4.11768f
C1472 BIT_SEL[27].n3 VSS 7.22573f
C1473 BIT_SEL[27].t2 VSS 4.11768f
C1474 BIT_SEL[27].n4 VSS 7.22573f
C1475 BIT_SEL[27].t6 VSS 4.11768f
C1476 BIT_SEL[27].n5 VSS 7.22573f
C1477 BIT_SEL[27].t3 VSS 4.11768f
C1478 BIT_SEL[27].n6 VSS 7.22573f
C1479 BIT_SEL[27].t0 VSS 4.3277f
C1480 a_14320_24255.t0 VSS 3.86539f
C1481 a_14320_24255.t1 VSS 2.23461f
C1482 a_20810_49151.t0 VSS 4.30261f
C1483 a_20810_49151.t1 VSS 1.69739f
C1484 a_20810_53186.t0 VSS 1.745f
C1485 a_20810_53186.t1 VSS 4.255f
C1486 a_14320_18908.t0 VSS 4.60993f
C1487 a_14320_18908.t1 VSS 1.39007f
C1488 a_20810_49679.t0 VSS 4.3173f
C1489 a_20810_49679.t1 VSS 1.6827f
C1490 BIT_SEL[53].t7 VSS 4.01572f
C1491 BIT_SEL[53].n0 VSS 6.88525f
C1492 BIT_SEL[53].t5 VSS 4.01572f
C1493 BIT_SEL[53].n1 VSS 6.88525f
C1494 BIT_SEL[53].t1 VSS 4.01572f
C1495 BIT_SEL[53].n2 VSS 6.88525f
C1496 BIT_SEL[53].t3 VSS 4.01572f
C1497 BIT_SEL[53].n3 VSS 6.88525f
C1498 BIT_SEL[53].t6 VSS 4.01572f
C1499 BIT_SEL[53].n4 VSS 6.88525f
C1500 BIT_SEL[53].t0 VSS 4.01572f
C1501 BIT_SEL[53].n5 VSS 6.88525f
C1502 BIT_SEL[53].t2 VSS 4.01572f
C1503 BIT_SEL[53].n6 VSS 6.88525f
C1504 BIT_SEL[53].t4 VSS 4.11021f
C1505 a_14320_8501.t0 VSS 3.86539f
C1506 a_14320_8501.t1 VSS 2.23461f
C1507 a_14320_1889.t0 VSS 4.30261f
C1508 a_14320_1889.t1 VSS 1.69739f
C1509 a_1340_61063.t0 VSS 4.25498f
C1510 a_1340_61063.t1 VSS 1.74502f
C1511 a_14320_42171.t0 VSS 4.34773f
C1512 a_14320_42171.t1 VSS 1.65227f
C1513 a_1340_32132.t0 VSS 3.86539f
C1514 a_1340_32132.t1 VSS 2.23461f
C1515 a_7830_41274.t0 VSS 1.69725f
C1516 a_7830_41274.t1 VSS 4.30275f
C1517 a_1340_33397.t0 VSS 4.30261f
C1518 a_1340_33397.t1 VSS 1.69739f
C1519 a_14320_53922.t0 VSS 1.91084f
C1520 a_14320_53922.t1 VSS 4.08916f
C1521 a_14320_7557.t0 VSS 2.354f
C1522 a_14320_7557.t1 VSS 3.746f
C1523 a_14320_47518.t0 VSS 2.41699f
C1524 a_14320_47518.t1 VSS 3.68301f
C1525 a_7830_1521.t0 VSS 1.79192f
C1526 a_7830_1521.t1 VSS 4.20808f
C1527 a_20810_21678.t0 VSS 1.745f
C1528 a_20810_21678.t1 VSS 4.255f
C1529 a_14320_11031.t0 VSS 1.39007f
C1530 a_14320_11031.t1 VSS 4.60993f
C1531 a_20810_54819.t0 VSS 3.74618f
C1532 a_20810_54819.t1 VSS 2.35382f
C1533 a_20810_40009.t0 VSS 3.86539f
C1534 a_20810_40009.t1 VSS 2.23461f
C1535 BIT_SEL[61].t3 VSS 4.14801f
C1536 BIT_SEL[61].n0 VSS 7.33197f
C1537 BIT_SEL[61].t5 VSS 4.14801f
C1538 BIT_SEL[61].n1 VSS 7.33197f
C1539 BIT_SEL[61].t7 VSS 4.14801f
C1540 BIT_SEL[61].n2 VSS 7.33197f
C1541 BIT_SEL[61].t0 VSS 4.14801f
C1542 BIT_SEL[61].n3 VSS 7.33197f
C1543 BIT_SEL[61].t2 VSS 4.14801f
C1544 BIT_SEL[61].n4 VSS 7.33197f
C1545 BIT_SEL[61].t4 VSS 4.14801f
C1546 BIT_SEL[61].n5 VSS 7.33197f
C1547 BIT_SEL[61].t1 VSS 4.14801f
C1548 BIT_SEL[61].n6 VSS 7.33197f
C1549 BIT_SEL[61].t6 VSS 4.41496f
C1550 a_1340_52289.t0 VSS 1.69351f
C1551 a_1340_52289.t1 VSS 4.30649f
C1552 a_7830_58293.t0 VSS 1.39007f
C1553 a_7830_58293.t1 VSS 4.60993f
C1554 a_14320_10663.t0 VSS 1.6522f
C1555 a_14320_10663.t1 VSS 4.3478f
C1556 a_1340_2786.t0 VSS 1.6522f
C1557 a_1340_2786.t1 VSS 4.3478f
C1558 a_20810_33925.t0 VSS 1.6826f
C1559 a_20810_33925.t1 VSS 4.3174f
C1560 a_7830_57556.t0 VSS 4.3173f
C1561 a_7830_57556.t1 VSS 1.6827f
C1562 a_14320_44412.t0 VSS 1.69351f
C1563 a_14320_44412.t1 VSS 4.30649f
C1564 a_14320_9029.t0 VSS 4.01916f
C1565 a_14320_9029.t1 VSS 1.98084f
C1566 a_7830_21149.t0 VSS 4.27849f
C1567 a_7830_21149.t1 VSS 1.72151f
C1568 a_20810_54451.t0 VSS 4.06398f
C1569 a_20810_54451.t1 VSS 2.23602f
C1570 a_14320_22414.t0 VSS 4.08932f
C1571 a_14320_22414.t1 VSS 1.91068f
C1572 a_1340_49151.t0 VSS 4.30261f
C1573 a_1340_49151.t1 VSS 1.69739f
C1574 a_20810_18171.t0 VSS 1.6826f
C1575 a_20810_18171.t1 VSS 4.3174f
C1576 a_20810_18908.t0 VSS 1.39007f
C1577 a_20810_18908.t1 VSS 4.60993f
C1578 a_7830_42539.t0 VSS 1.39007f
C1579 a_7830_42539.t1 VSS 4.60993f
C1580 a_7830_5395.t0 VSS 4.27849f
C1581 a_7830_5395.t1 VSS 1.72151f
C1582 a_14320_28658.t0 VSS 1.69351f
C1583 a_14320_28658.t1 VSS 4.30649f
C1584 a_7830_39641.t0 VSS 2.41699f
C1585 a_7830_39641.t1 VSS 3.68301f
C1586 a_7738_19835.t0 VSS 1.47655f
C1587 a_7738_19835.t1 VSS 4.52345f
C1588 a_7830_8501.t0 VSS 3.86539f
C1589 a_7830_8501.t1 VSS 2.23461f
C1590 BIT_SEL[29].t3 VSS 4.14801f
C1591 BIT_SEL[29].n0 VSS 7.33197f
C1592 BIT_SEL[29].t5 VSS 4.14801f
C1593 BIT_SEL[29].n1 VSS 7.33197f
C1594 BIT_SEL[29].t6 VSS 4.14801f
C1595 BIT_SEL[29].n2 VSS 7.33197f
C1596 BIT_SEL[29].t1 VSS 4.14801f
C1597 BIT_SEL[29].n3 VSS 7.33197f
C1598 BIT_SEL[29].t2 VSS 4.14801f
C1599 BIT_SEL[29].n4 VSS 7.33197f
C1600 BIT_SEL[29].t4 VSS 4.14801f
C1601 BIT_SEL[29].n5 VSS 7.33197f
C1602 BIT_SEL[29].t0 VSS 4.14801f
C1603 BIT_SEL[29].n6 VSS 7.33197f
C1604 BIT_SEL[29].t7 VSS 4.41496f
C1605 a_14320_22046.t0 VSS 3.66536f
C1606 a_14320_22046.t1 VSS 2.33464f
C1607 a_20810_38697.t0 VSS 4.06398f
C1608 a_20810_38697.t1 VSS 2.23602f
C1609 a_20718_51343.t0 VSS 1.47655f
C1610 a_20718_51343.t1 VSS 4.52345f
C1611 a_7830_26785.t0 VSS 1.39007f
C1612 a_7830_26785.t1 VSS 4.60993f
C1613 a_7830_23887.t0 VSS 2.41699f
C1614 a_7830_23887.t1 VSS 3.68301f
C1615 a_14320_48414.t0 VSS 4.01916f
C1616 a_14320_48414.t1 VSS 1.98084f
C1617 a_14320_50048.t0 VSS 1.6522f
C1618 a_14320_50048.t1 VSS 4.3478f
C1619 a_7830_26417.t0 VSS 4.34773f
C1620 a_7830_26417.t1 VSS 1.65227f
C1621 a_1340_17643.t0 VSS 4.30261f
C1622 a_1340_17643.t1 VSS 1.69739f
C1623 a_20810_32132.t0 VSS 2.23454f
C1624 a_20810_32132.t1 VSS 3.86546f
C1625 BIT_SEL[26].t1 VSS 4.02969f
C1626 BIT_SEL[26].n0 VSS 7.04511f
C1627 BIT_SEL[26].t3 VSS 4.02969f
C1628 BIT_SEL[26].n1 VSS 7.04511f
C1629 BIT_SEL[26].t6 VSS 4.02969f
C1630 BIT_SEL[26].n2 VSS 7.04511f
C1631 BIT_SEL[26].t0 VSS 4.02969f
C1632 BIT_SEL[26].n3 VSS 7.04511f
C1633 BIT_SEL[26].t2 VSS 4.02969f
C1634 BIT_SEL[26].n4 VSS 7.04511f
C1635 BIT_SEL[26].t4 VSS 4.02969f
C1636 BIT_SEL[26].n5 VSS 7.04511f
C1637 BIT_SEL[26].t5 VSS 4.2344f
C1638 BIT_SEL[26].t7 VSS 4.02969f
C1639 BIT_SEL[26].n6 VSS 7.04511f
C1640 a_7830_40906.t0 VSS 1.79192f
C1641 a_7830_40906.t1 VSS 4.20808f
C1642 a_7830_54451.t0 VSS 4.06398f
C1643 a_7830_54451.t1 VSS 2.23602f
C1644 a_14320_39641.t0 VSS 3.68292f
C1645 a_14320_39641.t1 VSS 2.41708f
C1646 BIT_SEL[47].t4 VSS 3.1518f
C1647 BIT_SEL[47].n0 VSS 5.61038f
C1648 BIT_SEL[47].t2 VSS 3.1518f
C1649 BIT_SEL[47].n1 VSS 5.61038f
C1650 BIT_SEL[47].t5 VSS 3.1518f
C1651 BIT_SEL[47].n2 VSS 5.61038f
C1652 BIT_SEL[47].t0 VSS 3.1518f
C1653 BIT_SEL[47].n3 VSS 5.61038f
C1654 BIT_SEL[47].t1 VSS 3.1518f
C1655 BIT_SEL[47].n4 VSS 5.61038f
C1656 BIT_SEL[47].t3 VSS 3.1518f
C1657 BIT_SEL[47].n5 VSS 5.61038f
C1658 BIT_SEL[47].t6 VSS 3.1518f
C1659 BIT_SEL[47].n6 VSS 5.61038f
C1660 BIT_SEL[47].t7 VSS 3.38636f
C1661 a_14320_56291.t0 VSS 4.01916f
C1662 a_14320_56291.t1 VSS 1.98084f
C1663 a_7830_8133.t0 VSS 3.68292f
C1664 a_7830_8133.t1 VSS 2.41708f
C1665 a_1248_35589.t0 VSS 4.52345f
C1666 a_1248_35589.t1 VSS 1.47655f
C1667 a_1340_17275.t0 VSS 4.20807f
C1668 a_1340_17275.t1 VSS 1.79193f
C1669 a_20810_16378.t0 VSS 3.86539f
C1670 a_20810_16378.t1 VSS 2.23461f
C1671 a_14320_39065.t0 VSS 2.354f
C1672 a_14320_39065.t1 VSS 3.746f
C1673 a_1340_31764.t0 VSS 3.68292f
C1674 a_1340_31764.t1 VSS 2.41708f
C1675 a_14320_16906.t0 VSS 4.01916f
C1676 a_14320_16906.t1 VSS 1.98084f
C1677 BIT_SEL[43].t0 VSS 4.11768f
C1678 BIT_SEL[43].n0 VSS 7.22573f
C1679 BIT_SEL[43].t3 VSS 4.11768f
C1680 BIT_SEL[43].n1 VSS 7.22573f
C1681 BIT_SEL[43].t6 VSS 4.11768f
C1682 BIT_SEL[43].n2 VSS 7.22573f
C1683 BIT_SEL[43].t4 VSS 4.11768f
C1684 BIT_SEL[43].n3 VSS 7.22573f
C1685 BIT_SEL[43].t1 VSS 4.11768f
C1686 BIT_SEL[43].n4 VSS 7.22573f
C1687 BIT_SEL[43].t5 VSS 4.11768f
C1688 BIT_SEL[43].n5 VSS 7.22573f
C1689 BIT_SEL[43].t2 VSS 4.11768f
C1690 BIT_SEL[43].n6 VSS 7.22573f
C1691 BIT_SEL[43].t7 VSS 4.3277f
C1692 a_20810_13272.t0 VSS 1.7215f
C1693 a_20810_13272.t1 VSS 4.2785f
C1694 a_1248_19835.t0 VSS 4.52345f
C1695 a_1248_19835.t1 VSS 1.47655f
C1696 a_7830_36903.t0 VSS 4.27849f
C1697 a_7830_36903.t1 VSS 1.72151f
C1698 a_7830_52289.t0 VSS 1.69351f
C1699 a_7830_52289.t1 VSS 4.30649f
C1700 a_14320_22943.t0 VSS 4.06398f
C1701 a_14320_22943.t1 VSS 2.23602f
C1702 a_20810_34662.t0 VSS 1.39007f
C1703 a_20810_34662.t1 VSS 4.60993f
C1704 a_1340_16010.t0 VSS 3.68292f
C1705 a_1340_16010.t1 VSS 2.41708f
C1706 a_1340_31188.t0 VSS 3.74618f
C1707 a_1340_31188.t1 VSS 2.35382f
C1708 a_14320_49151.t0 VSS 1.69725f
C1709 a_14320_49151.t1 VSS 4.30275f
C1710 a_7830_9766.t0 VSS 1.69725f
C1711 a_7830_9766.t1 VSS 4.30275f
C1712 a_14320_53186.t0 VSS 1.745f
C1713 a_14320_53186.t1 VSS 4.255f
C1714 a_20810_34294.t0 VSS 4.34773f
C1715 a_20810_34294.t1 VSS 1.65227f
C1716 a_20810_50048.t0 VSS 4.34773f
C1717 a_20810_50048.t1 VSS 1.65227f
C1718 a_14320_49679.t0 VSS 4.3173f
C1719 a_14320_49679.t1 VSS 1.6827f
C1720 a_7830_9398.t0 VSS 1.79192f
C1721 a_7830_9398.t1 VSS 4.20808f
C1722 a_20810_46045.t0 VSS 4.08932f
C1723 a_20810_46045.t1 VSS 1.91068f
C1724 a_1340_37800.t0 VSS 3.66536f
C1725 a_1340_37800.t1 VSS 2.33464f
C1726 a_7830_20781.t0 VSS 1.69351f
C1727 a_7830_20781.t1 VSS 4.30649f
C1728 a_7830_37432.t0 VSS 1.745f
C1729 a_7830_37432.t1 VSS 4.255f
C1730 a_20810_56291.t0 VSS 1.98079f
C1731 a_20810_56291.t1 VSS 4.01921f
C1732 a_7830_38168.t0 VSS 1.91084f
C1733 a_7830_38168.t1 VSS 4.08916f
C1734 a_1340_48783.t0 VSS 4.20807f
C1735 a_1340_48783.t1 VSS 1.79193f
C1736 a_20810_55395.t0 VSS 3.68292f
C1737 a_20810_55395.t1 VSS 2.41708f
C1738 a_7830_5027.t0 VSS 1.69351f
C1739 a_7830_5027.t1 VSS 4.30649f
C1740 BIT_SEL[6].t0 VSS 4.07324f
C1741 BIT_SEL[6].n0 VSS 7.01202f
C1742 BIT_SEL[6].t3 VSS 4.07324f
C1743 BIT_SEL[6].n1 VSS 7.01202f
C1744 BIT_SEL[6].t5 VSS 4.07324f
C1745 BIT_SEL[6].n2 VSS 7.01202f
C1746 BIT_SEL[6].t1 VSS 4.07324f
C1747 BIT_SEL[6].n3 VSS 7.01202f
C1748 BIT_SEL[6].t2 VSS 4.07324f
C1749 BIT_SEL[6].n4 VSS 7.01202f
C1750 BIT_SEL[6].t4 VSS 4.07324f
C1751 BIT_SEL[6].n5 VSS 7.01202f
C1752 BIT_SEL[6].t6 VSS 4.07324f
C1753 BIT_SEL[6].n6 VSS 7.01202f
C1754 BIT_SEL[6].t7 VSS 4.21129f
C1755 a_7830_21678.t0 VSS 1.745f
C1756 a_7830_21678.t1 VSS 4.255f
C1757 a_1340_22046.t0 VSS 2.33483f
C1758 a_1340_22046.t1 VSS 3.66517f
C1759 a_20810_60166.t0 VSS 4.30649f
C1760 a_20810_60166.t1 VSS 1.69351f
C1761 a_7830_22414.t0 VSS 1.91084f
C1762 a_7830_22414.t1 VSS 4.08916f
C1763 a_14320_21678.t0 VSS 4.25498f
C1764 a_14320_21678.t1 VSS 1.74502f
C1765 a_14320_2417.t0 VSS 4.3173f
C1766 a_14320_2417.t1 VSS 1.6827f
C1767 BIT_SEL[37].t7 VSS 4.01572f
C1768 BIT_SEL[37].n0 VSS 6.88525f
C1769 BIT_SEL[37].t5 VSS 4.01572f
C1770 BIT_SEL[37].n1 VSS 6.88525f
C1771 BIT_SEL[37].t2 VSS 4.01572f
C1772 BIT_SEL[37].n2 VSS 6.88525f
C1773 BIT_SEL[37].t4 VSS 4.01572f
C1774 BIT_SEL[37].n3 VSS 6.88525f
C1775 BIT_SEL[37].t6 VSS 4.01572f
C1776 BIT_SEL[37].n4 VSS 6.88525f
C1777 BIT_SEL[37].t1 VSS 4.01572f
C1778 BIT_SEL[37].n5 VSS 6.88525f
C1779 BIT_SEL[37].t3 VSS 4.01572f
C1780 BIT_SEL[37].n6 VSS 6.88525f
C1781 BIT_SEL[37].t0 VSS 4.11021f
C1782 a_1340_5395.t0 VSS 4.27849f
C1783 a_1340_5395.t1 VSS 1.72151f
C1784 BIT_SEL[4].t7 VSS 4.02347f
C1785 BIT_SEL[4].n0 VSS 6.87043f
C1786 BIT_SEL[4].t5 VSS 4.02347f
C1787 BIT_SEL[4].n1 VSS 6.87043f
C1788 BIT_SEL[4].t1 VSS 4.02347f
C1789 BIT_SEL[4].n2 VSS 6.87043f
C1790 BIT_SEL[4].t3 VSS 4.02347f
C1791 BIT_SEL[4].n3 VSS 6.87043f
C1792 BIT_SEL[4].t2 VSS 4.02347f
C1793 BIT_SEL[4].n4 VSS 6.87043f
C1794 BIT_SEL[4].t4 VSS 4.02347f
C1795 BIT_SEL[4].n5 VSS 6.87043f
C1796 BIT_SEL[4].t6 VSS 4.11755f
C1797 BIT_SEL[4].t0 VSS 4.02347f
C1798 BIT_SEL[4].n6 VSS 6.87043f
C1799 a_7830_60166.t0 VSS 1.69351f
C1800 a_7830_60166.t1 VSS 4.30649f
C1801 a_1340_624.t0 VSS 2.23454f
C1802 a_1340_624.t1 VSS 3.86546f
C1803 a_1340_33029.t0 VSS 4.20807f
C1804 a_1340_33029.t1 VSS 1.79193f
C1805 a_1340_62696.t0 VSS 3.74618f
C1806 a_1340_62696.t1 VSS 2.35382f
C1807 a_20810_14537.t0 VSS 4.08932f
C1808 a_20810_14537.t1 VSS 1.91068f
C1809 a_14320_54819.t0 VSS 2.354f
C1810 a_14320_54819.t1 VSS 3.746f
C1811 BIT_SEL[46].t2 VSS 4.1517f
C1812 BIT_SEL[46].n0 VSS 7.36453f
C1813 BIT_SEL[46].t4 VSS 4.1517f
C1814 BIT_SEL[46].n1 VSS 7.36453f
C1815 BIT_SEL[46].t6 VSS 4.1517f
C1816 BIT_SEL[46].n2 VSS 7.36453f
C1817 BIT_SEL[46].t1 VSS 4.1517f
C1818 BIT_SEL[46].n3 VSS 7.36453f
C1819 BIT_SEL[46].t3 VSS 4.1517f
C1820 BIT_SEL[46].n4 VSS 7.36453f
C1821 BIT_SEL[46].t0 VSS 4.1517f
C1822 BIT_SEL[46].n5 VSS 7.36453f
C1823 BIT_SEL[46].t5 VSS 4.45988f
C1824 BIT_SEL[46].t7 VSS 4.1517f
C1825 BIT_SEL[46].n6 VSS 7.36453f
C1826 a_14320_33925.t0 VSS 1.6826f
C1827 a_14320_33925.t1 VSS 4.3174f
C1828 a_14320_40009.t0 VSS 3.86539f
C1829 a_14320_40009.t1 VSS 2.23461f
C1830 BIT_SEL[45].t2 VSS 4.14801f
C1831 BIT_SEL[45].n0 VSS 7.33197f
C1832 BIT_SEL[45].t4 VSS 4.14801f
C1833 BIT_SEL[45].n1 VSS 7.33197f
C1834 BIT_SEL[45].t5 VSS 4.14801f
C1835 BIT_SEL[45].n2 VSS 7.33197f
C1836 BIT_SEL[45].t0 VSS 4.14801f
C1837 BIT_SEL[45].n3 VSS 7.33197f
C1838 BIT_SEL[45].t1 VSS 4.14801f
C1839 BIT_SEL[45].n4 VSS 7.33197f
C1840 BIT_SEL[45].t3 VSS 4.14801f
C1841 BIT_SEL[45].n5 VSS 7.33197f
C1842 BIT_SEL[45].t6 VSS 4.14801f
C1843 BIT_SEL[45].n6 VSS 7.33197f
C1844 BIT_SEL[45].t7 VSS 4.41496f
C1845 a_20810_14169.t0 VSS 2.33483f
C1846 a_20810_14169.t1 VSS 3.66517f
C1847 a_7830_10294.t0 VSS 4.3173f
C1848 a_7830_10294.t1 VSS 1.6827f
C1849 a_1340_5924.t0 VSS 1.745f
C1850 a_1340_5924.t1 VSS 4.255f
C1851 a_1340_40537.t0 VSS 4.01916f
C1852 a_1340_40537.t1 VSS 1.98084f
C1853 a_7830_37800.t0 VSS 2.33483f
C1854 a_7830_37800.t1 VSS 3.66517f
C1855 BIT_SEL[24].t3 VSS 4.14071f
C1856 BIT_SEL[24].n0 VSS 7.18434f
C1857 BIT_SEL[24].t5 VSS 4.14071f
C1858 BIT_SEL[24].n1 VSS 7.18434f
C1859 BIT_SEL[24].t6 VSS 4.14071f
C1860 BIT_SEL[24].n2 VSS 7.18434f
C1861 BIT_SEL[24].t0 VSS 4.14071f
C1862 BIT_SEL[24].n3 VSS 7.18434f
C1863 BIT_SEL[24].t1 VSS 4.14071f
C1864 BIT_SEL[24].n4 VSS 7.18434f
C1865 BIT_SEL[24].t4 VSS 4.14071f
C1866 BIT_SEL[24].n5 VSS 7.18434f
C1867 BIT_SEL[24].t2 VSS 4.31483f
C1868 BIT_SEL[24].t7 VSS 4.14071f
C1869 BIT_SEL[24].n6 VSS 7.18434f
C1870 a_14320_54451.t0 VSS 4.06398f
C1871 a_14320_54451.t1 VSS 2.23602f
C1872 a_7830_39065.t0 VSS 2.354f
C1873 a_7830_39065.t1 VSS 3.746f
C1874 a_14320_18171.t0 VSS 1.6826f
C1875 a_14320_18171.t1 VSS 4.3174f
C1876 a_20810_5924.t0 VSS 1.745f
C1877 a_20810_5924.t1 VSS 4.255f
C1878 a_1340_24783.t0 VSS 4.01916f
C1879 a_1340_24783.t1 VSS 1.98084f
C1880 a_14320_5027.t0 VSS 1.69351f
C1881 a_14320_5027.t1 VSS 4.30649f
C1882 a_14320_38697.t0 VSS 4.06398f
C1883 a_14320_38697.t1 VSS 2.23602f
C1884 BIT_SEL[44].t5 VSS 4.12331f
C1885 BIT_SEL[44].n0 VSS 7.26213f
C1886 BIT_SEL[44].t6 VSS 4.12331f
C1887 BIT_SEL[44].n1 VSS 7.26213f
C1888 BIT_SEL[44].t2 VSS 4.12331f
C1889 BIT_SEL[44].n2 VSS 7.26213f
C1890 BIT_SEL[44].t0 VSS 4.12331f
C1891 BIT_SEL[44].n3 VSS 7.26213f
C1892 BIT_SEL[44].t3 VSS 4.12331f
C1893 BIT_SEL[44].n4 VSS 7.26213f
C1894 BIT_SEL[44].t1 VSS 4.12331f
C1895 BIT_SEL[44].n5 VSS 7.26213f
C1896 BIT_SEL[44].t4 VSS 4.3879f
C1897 BIT_SEL[44].t7 VSS 4.12331f
C1898 BIT_SEL[44].n6 VSS 7.26213f
C1899 a_14228_51343.t0 VSS 4.52345f
C1900 a_14228_51343.t1 VSS 1.47655f
C1901 a_1340_61799.t0 VSS 4.08932f
C1902 a_1340_61799.t1 VSS 1.91068f
C1903 a_7830_23311.t0 VSS 3.74618f
C1904 a_7830_23311.t1 VSS 2.35382f
C1905 a_1340_28658.t0 VSS 4.30649f
C1906 a_1340_28658.t1 VSS 1.69351f
C1907 BIT_SEL[2].t7 VSS 4.05315f
C1908 BIT_SEL[2].n0 VSS 6.86345f
C1909 BIT_SEL[2].t5 VSS 4.05315f
C1910 BIT_SEL[2].n1 VSS 6.86345f
C1911 BIT_SEL[2].t3 VSS 4.05315f
C1912 BIT_SEL[2].n2 VSS 6.86345f
C1913 BIT_SEL[2].t0 VSS 4.05315f
C1914 BIT_SEL[2].n3 VSS 6.86345f
C1915 BIT_SEL[2].t1 VSS 4.05315f
C1916 BIT_SEL[2].n4 VSS 6.86345f
C1917 BIT_SEL[2].t2 VSS 4.05315f
C1918 BIT_SEL[2].n5 VSS 6.86345f
C1919 BIT_SEL[2].t4 VSS 4.05315f
C1920 BIT_SEL[2].n6 VSS 6.86345f
C1921 BIT_SEL[2].t6 VSS 4.12109f
C1922 a_20810_12904.t0 VSS 4.30649f
C1923 a_20810_12904.t1 VSS 1.69351f
C1924 COL_PROG_N[4].t3 VSS 1.10931f
C1925 COL_PROG_N[4].n0 VSS 0.38563f
C1926 COL_PROG_N[4].t1 VSS 1.10931f
C1927 COL_PROG_N[4].n1 VSS 0.39369f
C1928 COL_PROG_N[4].t2 VSS 1.10931f
C1929 COL_PROG_N[4].n2 VSS 0.77937f
C1930 COL_PROG_N[4].t0 VSS 1.10971f
C1931 a_1340_50048.t0 VSS 1.6522f
C1932 a_1340_50048.t1 VSS 4.3478f
C1933 BIT_SEL[3].t6 VSS 4.04507f
C1934 BIT_SEL[3].n0 VSS 6.87869f
C1935 BIT_SEL[3].t3 VSS 4.04507f
C1936 BIT_SEL[3].n1 VSS 6.87869f
C1937 BIT_SEL[3].t4 VSS 4.04507f
C1938 BIT_SEL[3].n2 VSS 6.87869f
C1939 BIT_SEL[3].t5 VSS 4.04507f
C1940 BIT_SEL[3].n3 VSS 6.87869f
C1941 BIT_SEL[3].t7 VSS 4.04507f
C1942 BIT_SEL[3].n4 VSS 6.87869f
C1943 BIT_SEL[3].t0 VSS 4.04507f
C1944 BIT_SEL[3].n5 VSS 6.87869f
C1945 BIT_SEL[3].t2 VSS 4.04507f
C1946 BIT_SEL[3].n6 VSS 6.87869f
C1947 BIT_SEL[3].t1 VSS 4.1133f
C1948 a_7830_48783.t0 VSS 1.79192f
C1949 a_7830_48783.t1 VSS 4.20808f
C1950 a_1248_27712.t0 VSS 1.47655f
C1951 a_1248_27712.t1 VSS 4.52345f
C1952 a_7830_47886.t0 VSS 3.86539f
C1953 a_7830_47886.t1 VSS 2.23461f
C1954 a_20810_60534.t0 VSS 1.7215f
C1955 a_20810_60534.t1 VSS 4.2785f
C1956 a_1340_6660.t0 VSS 4.08932f
C1957 a_1340_6660.t1 VSS 1.91068f
C1958 BIT_SEL[10].t0 VSS 4.02969f
C1959 BIT_SEL[10].n0 VSS 7.04511f
C1960 BIT_SEL[10].t2 VSS 4.02969f
C1961 BIT_SEL[10].n1 VSS 7.04511f
C1962 BIT_SEL[10].t4 VSS 4.02969f
C1963 BIT_SEL[10].n2 VSS 7.04511f
C1964 BIT_SEL[10].t7 VSS 4.02969f
C1965 BIT_SEL[10].n3 VSS 7.04511f
C1966 BIT_SEL[10].t1 VSS 4.02969f
C1967 BIT_SEL[10].n4 VSS 7.04511f
C1968 BIT_SEL[10].t3 VSS 4.02969f
C1969 BIT_SEL[10].n5 VSS 7.04511f
C1970 BIT_SEL[10].t5 VSS 4.02969f
C1971 BIT_SEL[10].n6 VSS 7.04511f
C1972 BIT_SEL[10].t6 VSS 4.2344f
C1973 a_14320_32132.t0 VSS 3.86539f
C1974 a_14320_32132.t1 VSS 2.23461f
C1975 a_20810_61431.t0 VSS 2.33483f
C1976 a_20810_61431.t1 VSS 3.66517f
C1977 a_7830_41802.t0 VSS 4.3173f
C1978 a_7830_41802.t1 VSS 1.6827f
C1979 BIT_SEL[21].t1 VSS 4.01572f
C1980 BIT_SEL[21].n0 VSS 6.88525f
C1981 BIT_SEL[21].t7 VSS 4.01572f
C1982 BIT_SEL[21].n1 VSS 6.88525f
C1983 BIT_SEL[21].t4 VSS 4.01572f
C1984 BIT_SEL[21].n2 VSS 6.88525f
C1985 BIT_SEL[21].t6 VSS 4.01572f
C1986 BIT_SEL[21].n3 VSS 6.88525f
C1987 BIT_SEL[21].t0 VSS 4.01572f
C1988 BIT_SEL[21].n4 VSS 6.88525f
C1989 BIT_SEL[21].t2 VSS 4.01572f
C1990 BIT_SEL[21].n5 VSS 6.88525f
C1991 BIT_SEL[21].t5 VSS 4.01572f
C1992 BIT_SEL[21].n6 VSS 6.88525f
C1993 BIT_SEL[21].t3 VSS 4.11021f
C1994 a_20810_45677.t0 VSS 2.33483f
C1995 a_20810_45677.t1 VSS 3.66517f
C1996 a_14320_16378.t0 VSS 2.23454f
C1997 a_14320_16378.t1 VSS 3.86546f
C1998 a_7830_18540.t0 VSS 4.34773f
C1999 a_7830_18540.t1 VSS 1.65227f
C2000 BIT_SEL[19].t3 VSS 4.04507f
C2001 BIT_SEL[19].n0 VSS 6.87869f
C2002 BIT_SEL[19].t0 VSS 4.04507f
C2003 BIT_SEL[19].n1 VSS 6.87869f
C2004 BIT_SEL[19].t1 VSS 4.04507f
C2005 BIT_SEL[19].n2 VSS 6.87869f
C2006 BIT_SEL[19].t2 VSS 4.04507f
C2007 BIT_SEL[19].n3 VSS 6.87869f
C2008 BIT_SEL[19].t4 VSS 4.04507f
C2009 BIT_SEL[19].n4 VSS 6.87869f
C2010 BIT_SEL[19].t5 VSS 4.04507f
C2011 BIT_SEL[19].n5 VSS 6.87869f
C2012 BIT_SEL[19].t7 VSS 4.04507f
C2013 BIT_SEL[19].n6 VSS 6.87869f
C2014 BIT_SEL[19].t6 VSS 4.1133f
C2015 a_1340_18171.t0 VSS 4.3173f
C2016 a_1340_18171.t1 VSS 1.6827f
C2017 a_20810_45309.t0 VSS 1.745f
C2018 a_20810_45309.t1 VSS 4.255f
C2019 a_14320_13272.t0 VSS 4.27849f
C2020 a_14320_13272.t1 VSS 1.72151f
C2021 a_14320_53554.t0 VSS 2.33483f
C2022 a_14320_53554.t1 VSS 3.66517f
C2023 a_14320_34662.t0 VSS 1.39007f
C2024 a_14320_34662.t1 VSS 4.60993f
C2025 BIT_SEL[33].t1 VSS 4.07792f
C2026 BIT_SEL[33].n0 VSS 6.88058f
C2027 BIT_SEL[33].t4 VSS 4.07792f
C2028 BIT_SEL[33].n1 VSS 6.88058f
C2029 BIT_SEL[33].t5 VSS 4.07792f
C2030 BIT_SEL[33].n2 VSS 6.88058f
C2031 BIT_SEL[33].t0 VSS 4.07792f
C2032 BIT_SEL[33].n3 VSS 6.88058f
C2033 BIT_SEL[33].t6 VSS 4.07792f
C2034 BIT_SEL[33].n4 VSS 6.88058f
C2035 BIT_SEL[33].t2 VSS 4.07792f
C2036 BIT_SEL[33].n5 VSS 6.88058f
C2037 BIT_SEL[33].t7 VSS 4.07792f
C2038 BIT_SEL[33].n6 VSS 6.88058f
C2039 BIT_SEL[33].t3 VSS 4.12246f
C2040 a_1340_44780.t0 VSS 1.7215f
C2041 a_1340_44780.t1 VSS 4.2785f
C2042 SENSE.t7 VSS 0.24927f
C2043 SENSE.t3 VSS 0.24927f
C2044 SENSE.n0 VSS 4.53187f
C2045 SENSE.t6 VSS 0.24927f
C2046 SENSE.t0 VSS 0.24927f
C2047 SENSE.n1 VSS 4.53012f
C2048 SENSE.t4 VSS 0.24927f
C2049 SENSE.n2 VSS 4.531f
C2050 SENSE.t2 VSS 0.24927f
C2051 SENSE.n3 VSS 4.531f
C2052 SENSE.t5 VSS 0.24927f
C2053 SENSE.n4 VSS 4.531f
C2054 SENSE.t1 VSS 0.24927f
C2055 SENSE.n5 VSS 4.531f
C2056 a_7830_6660.t0 VSS 1.91084f
C2057 a_7830_6660.t1 VSS 4.08916f
C2058 a_14320_34294.t0 VSS 1.6522f
C2059 a_14320_34294.t1 VSS 4.3478f
C2060 BIT_SEL[35].t1 VSS 4.04507f
C2061 BIT_SEL[35].n0 VSS 6.87869f
C2062 BIT_SEL[35].t6 VSS 4.04507f
C2063 BIT_SEL[35].n1 VSS 6.87869f
C2064 BIT_SEL[35].t7 VSS 4.04507f
C2065 BIT_SEL[35].n2 VSS 6.87869f
C2066 BIT_SEL[35].t0 VSS 4.04507f
C2067 BIT_SEL[35].n3 VSS 6.87869f
C2068 BIT_SEL[35].t2 VSS 4.04507f
C2069 BIT_SEL[35].n4 VSS 6.87869f
C2070 BIT_SEL[35].t4 VSS 4.04507f
C2071 BIT_SEL[35].n5 VSS 6.87869f
C2072 BIT_SEL[35].t5 VSS 4.04507f
C2073 BIT_SEL[35].n6 VSS 6.87869f
C2074 BIT_SEL[35].t3 VSS 4.1133f
C2075 BIT_SEL[0].t4 VSS 3.0317f
C2076 BIT_SEL[0].n0 VSS 5.09227f
C2077 BIT_SEL[0].t6 VSS 3.0317f
C2078 BIT_SEL[0].n1 VSS 5.09227f
C2079 BIT_SEL[0].t1 VSS 3.0317f
C2080 BIT_SEL[0].n2 VSS 5.09227f
C2081 BIT_SEL[0].t2 VSS 3.0317f
C2082 BIT_SEL[0].n3 VSS 5.09227f
C2083 BIT_SEL[0].t5 VSS 3.0317f
C2084 BIT_SEL[0].n4 VSS 5.09227f
C2085 BIT_SEL[0].t3 VSS 3.0317f
C2086 BIT_SEL[0].n5 VSS 5.09227f
C2087 BIT_SEL[0].t0 VSS 3.06458f
C2088 BIT_SEL[0].t7 VSS 3.0317f
C2089 BIT_SEL[0].n6 VSS 5.09227f
C2090 a_1340_24255.t0 VSS 3.86539f
C2091 a_1340_24255.t1 VSS 2.23461f
C2092 a_7830_33397.t0 VSS 1.69725f
C2093 a_7830_33397.t1 VSS 4.30275f
C2094 a_20810_62328.t0 VSS 4.06398f
C2095 a_20810_62328.t1 VSS 2.23602f
C2096 a_7830_44412.t0 VSS 4.30649f
C2097 a_7830_44412.t1 VSS 1.69351f
C2098 BIT_SEL[18].t5 VSS 4.05315f
C2099 BIT_SEL[18].n0 VSS 6.86345f
C2100 BIT_SEL[18].t3 VSS 4.05315f
C2101 BIT_SEL[18].n1 VSS 6.86345f
C2102 BIT_SEL[18].t1 VSS 4.05315f
C2103 BIT_SEL[18].n2 VSS 6.86345f
C2104 BIT_SEL[18].t6 VSS 4.05315f
C2105 BIT_SEL[18].n3 VSS 6.86345f
C2106 BIT_SEL[18].t7 VSS 4.05315f
C2107 BIT_SEL[18].n4 VSS 6.86345f
C2108 BIT_SEL[18].t0 VSS 4.05315f
C2109 BIT_SEL[18].n5 VSS 6.86345f
C2110 BIT_SEL[18].t2 VSS 4.05315f
C2111 BIT_SEL[18].n6 VSS 6.86345f
C2112 BIT_SEL[18].t4 VSS 4.12109f
C2113 a_1340_29026.t0 VSS 1.7215f
C2114 a_1340_29026.t1 VSS 4.2785f
C2115 a_14320_46045.t0 VSS 4.08932f
C2116 a_14320_46045.t1 VSS 1.91068f
C2117 a_20810_13801.t0 VSS 4.25498f
C2118 a_20810_13801.t1 VSS 1.74502f
C2119 a_14320_60534.t0 VSS 4.27849f
C2120 a_14320_60534.t1 VSS 1.72151f
C2121 BIT_SEL[36].t2 VSS 4.02347f
C2122 BIT_SEL[36].n0 VSS 6.87043f
C2123 BIT_SEL[36].t1 VSS 4.02347f
C2124 BIT_SEL[36].n1 VSS 6.87043f
C2125 BIT_SEL[36].t7 VSS 4.02347f
C2126 BIT_SEL[36].n2 VSS 6.87043f
C2127 BIT_SEL[36].t3 VSS 4.02347f
C2128 BIT_SEL[36].n3 VSS 6.87043f
C2129 BIT_SEL[36].t5 VSS 4.02347f
C2130 BIT_SEL[36].n4 VSS 6.87043f
C2131 BIT_SEL[36].t4 VSS 4.02347f
C2132 BIT_SEL[36].n5 VSS 6.87043f
C2133 BIT_SEL[36].t6 VSS 4.02347f
C2134 BIT_SEL[36].n6 VSS 6.87043f
C2135 BIT_SEL[36].t0 VSS 4.11755f
C2136 a_7830_17643.t0 VSS 1.69725f
C2137 a_7830_17643.t1 VSS 4.30275f
C2138 a_20810_8133.t0 VSS 3.68292f
C2139 a_20810_8133.t1 VSS 2.41708f
C2140 BIT_SEL[63].t0 VSS 3.1518f
C2141 BIT_SEL[63].n0 VSS 5.61038f
C2142 BIT_SEL[63].t6 VSS 3.1518f
C2143 BIT_SEL[63].n1 VSS 5.61038f
C2144 BIT_SEL[63].t3 VSS 3.1518f
C2145 BIT_SEL[63].n2 VSS 5.61038f
C2146 BIT_SEL[63].t7 VSS 3.1518f
C2147 BIT_SEL[63].n3 VSS 5.61038f
C2148 BIT_SEL[63].t1 VSS 3.1518f
C2149 BIT_SEL[63].n4 VSS 5.61038f
C2150 BIT_SEL[63].t2 VSS 3.1518f
C2151 BIT_SEL[63].n5 VSS 5.61038f
C2152 BIT_SEL[63].t4 VSS 3.1518f
C2153 BIT_SEL[63].n6 VSS 5.61038f
C2154 BIT_SEL[63].t5 VSS 3.38636f
C2155 a_1340_22943.t0 VSS 4.06398f
C2156 a_1340_22943.t1 VSS 2.23602f
C2157 BIT_SEL[12].t7 VSS 4.12331f
C2158 BIT_SEL[12].n0 VSS 7.26213f
C2159 BIT_SEL[12].t0 VSS 4.12331f
C2160 BIT_SEL[12].n1 VSS 7.26213f
C2161 BIT_SEL[12].t4 VSS 4.12331f
C2162 BIT_SEL[12].n2 VSS 7.26213f
C2163 BIT_SEL[12].t2 VSS 4.12331f
C2164 BIT_SEL[12].n3 VSS 7.26213f
C2165 BIT_SEL[12].t5 VSS 4.12331f
C2166 BIT_SEL[12].n4 VSS 7.26213f
C2167 BIT_SEL[12].t3 VSS 4.12331f
C2168 BIT_SEL[12].n5 VSS 7.26213f
C2169 BIT_SEL[12].t6 VSS 4.3879f
C2170 BIT_SEL[12].t1 VSS 4.12331f
C2171 BIT_SEL[12].n6 VSS 7.26213f
C2172 PRESET_N.t19 VSS 0.25481f
C2173 PRESET_N.n0 VSS 0.52194f
C2174 PRESET_N.t18 VSS 0.25481f
C2175 PRESET_N.n1 VSS 0.52127f
C2176 PRESET_N.t1 VSS 0.2583f
C2177 PRESET_N.n2 VSS 2.6482f
C2178 PRESET_N.t15 VSS 0.25481f
C2179 PRESET_N.n3 VSS 0.52194f
C2180 PRESET_N.t22 VSS 0.25481f
C2181 PRESET_N.n4 VSS 0.52127f
C2182 PRESET_N.t6 VSS 0.2583f
C2183 PRESET_N.n5 VSS 2.6482f
C2184 PRESET_N.t20 VSS 0.25481f
C2185 PRESET_N.n6 VSS 0.52194f
C2186 PRESET_N.t0 VSS 0.25481f
C2187 PRESET_N.n7 VSS 0.52127f
C2188 PRESET_N.t13 VSS 0.2583f
C2189 PRESET_N.n8 VSS 2.6482f
C2190 PRESET_N.t4 VSS 0.25481f
C2191 PRESET_N.n9 VSS 0.52194f
C2192 PRESET_N.t2 VSS 0.25481f
C2193 PRESET_N.n10 VSS 0.52127f
C2194 PRESET_N.t7 VSS 0.2583f
C2195 PRESET_N.n11 VSS 2.6482f
C2196 PRESET_N.t9 VSS 0.25481f
C2197 PRESET_N.n12 VSS 0.52194f
C2198 PRESET_N.t8 VSS 0.25481f
C2199 PRESET_N.n13 VSS 0.52127f
C2200 PRESET_N.t10 VSS 0.2583f
C2201 PRESET_N.n14 VSS 2.6482f
C2202 PRESET_N.t17 VSS 0.25481f
C2203 PRESET_N.n15 VSS 0.52194f
C2204 PRESET_N.t23 VSS 0.25481f
C2205 PRESET_N.n16 VSS 0.52127f
C2206 PRESET_N.t5 VSS 0.2583f
C2207 PRESET_N.n17 VSS 2.6482f
C2208 PRESET_N.t3 VSS 0.25481f
C2209 PRESET_N.n18 VSS 0.52194f
C2210 PRESET_N.t11 VSS 0.25481f
C2211 PRESET_N.n19 VSS 0.52127f
C2212 PRESET_N.t14 VSS 0.2583f
C2213 PRESET_N.n20 VSS 2.6482f
C2214 PRESET_N.t12 VSS 0.25481f
C2215 PRESET_N.n21 VSS 0.51783f
C2216 PRESET_N.t16 VSS 0.25481f
C2217 PRESET_N.n22 VSS 0.52127f
C2218 PRESET_N.t21 VSS 0.2583f
C2219 a_14320_58293.t0 VSS 1.39007f
C2220 a_14320_58293.t1 VSS 4.60993f
C2221 a_14320_60166.t0 VSS 1.69351f
C2222 a_14320_60166.t1 VSS 4.30649f
C2223 a_1340_13272.t0 VSS 4.27849f
C2224 a_1340_13272.t1 VSS 1.72151f
C2225 BIT_SEL[32].t0 VSS 3.0317f
C2226 BIT_SEL[32].n0 VSS 5.09227f
C2227 BIT_SEL[32].t5 VSS 3.0317f
C2228 BIT_SEL[32].n1 VSS 5.09227f
C2229 BIT_SEL[32].t7 VSS 3.0317f
C2230 BIT_SEL[32].n2 VSS 5.09227f
C2231 BIT_SEL[32].t2 VSS 3.0317f
C2232 BIT_SEL[32].n3 VSS 5.09227f
C2233 BIT_SEL[32].t3 VSS 3.0317f
C2234 BIT_SEL[32].n4 VSS 5.09227f
C2235 BIT_SEL[32].t6 VSS 3.0317f
C2236 BIT_SEL[32].n5 VSS 5.09227f
C2237 BIT_SEL[32].t4 VSS 3.0317f
C2238 BIT_SEL[32].n6 VSS 5.09227f
C2239 BIT_SEL[32].t1 VSS 3.06458f
C2240 a_20810_41274.t0 VSS 4.30261f
C2241 a_20810_41274.t1 VSS 1.69739f
C2242 BIT_SEL[55].t4 VSS 4.06977f
C2243 BIT_SEL[55].n0 VSS 7.03381f
C2244 BIT_SEL[55].t6 VSS 4.06977f
C2245 BIT_SEL[55].n1 VSS 7.03381f
C2246 BIT_SEL[55].t7 VSS 4.06977f
C2247 BIT_SEL[55].n2 VSS 7.03381f
C2248 BIT_SEL[55].t0 VSS 4.06977f
C2249 BIT_SEL[55].n3 VSS 7.03381f
C2250 BIT_SEL[55].t5 VSS 4.06977f
C2251 BIT_SEL[55].n4 VSS 7.03381f
C2252 BIT_SEL[55].t2 VSS 4.06977f
C2253 BIT_SEL[55].n5 VSS 7.03381f
C2254 BIT_SEL[55].t1 VSS 4.06977f
C2255 BIT_SEL[55].n6 VSS 7.03381f
C2256 BIT_SEL[55].t3 VSS 4.20835f
C2257 a_14320_36535.t0 VSS 1.69351f
C2258 a_14320_36535.t1 VSS 4.30649f
C2259 a_1340_1521.t0 VSS 4.20807f
C2260 a_1340_1521.t1 VSS 1.79193f
C2261 BIT_SEL[9].t7 VSS 4.14534f
C2262 BIT_SEL[9].n0 VSS 7.22001f
C2263 BIT_SEL[9].t3 VSS 4.14534f
C2264 BIT_SEL[9].n1 VSS 7.22001f
C2265 BIT_SEL[9].t5 VSS 4.14534f
C2266 BIT_SEL[9].n2 VSS 7.22001f
C2267 BIT_SEL[9].t1 VSS 4.14534f
C2268 BIT_SEL[9].n3 VSS 7.22001f
C2269 BIT_SEL[9].t6 VSS 4.14534f
C2270 BIT_SEL[9].n4 VSS 7.22001f
C2271 BIT_SEL[9].t2 VSS 4.14534f
C2272 BIT_SEL[9].n5 VSS 7.22001f
C2273 BIT_SEL[9].t4 VSS 4.14534f
C2274 BIT_SEL[9].n6 VSS 7.22001f
C2275 BIT_SEL[9].t0 VSS 4.32038f
C2276 a_14320_14537.t0 VSS 4.08932f
C2277 a_14320_14537.t1 VSS 1.91068f
C2278 BIT_SEL[42].t0 VSS 4.02969f
C2279 BIT_SEL[42].n0 VSS 7.04511f
C2280 BIT_SEL[42].t2 VSS 4.02969f
C2281 BIT_SEL[42].n1 VSS 7.04511f
C2282 BIT_SEL[42].t5 VSS 4.02969f
C2283 BIT_SEL[42].n2 VSS 7.04511f
C2284 BIT_SEL[42].t7 VSS 4.02969f
C2285 BIT_SEL[42].n3 VSS 7.04511f
C2286 BIT_SEL[42].t1 VSS 4.02969f
C2287 BIT_SEL[42].n4 VSS 7.04511f
C2288 BIT_SEL[42].t3 VSS 4.02969f
C2289 BIT_SEL[42].n5 VSS 7.04511f
C2290 BIT_SEL[42].t4 VSS 4.2344f
C2291 BIT_SEL[42].t6 VSS 4.02969f
C2292 BIT_SEL[42].n6 VSS 7.04511f
C2293 a_1340_33925.t0 VSS 4.3173f
C2294 a_1340_33925.t1 VSS 1.6827f
C2295 BIT_SEL[5].t3 VSS 4.01572f
C2296 BIT_SEL[5].n0 VSS 6.88525f
C2297 BIT_SEL[5].t1 VSS 4.01572f
C2298 BIT_SEL[5].n1 VSS 6.88525f
C2299 BIT_SEL[5].t5 VSS 4.01572f
C2300 BIT_SEL[5].n2 VSS 6.88525f
C2301 BIT_SEL[5].t0 VSS 4.01572f
C2302 BIT_SEL[5].n3 VSS 6.88525f
C2303 BIT_SEL[5].t2 VSS 4.01572f
C2304 BIT_SEL[5].n4 VSS 6.88525f
C2305 BIT_SEL[5].t4 VSS 4.01572f
C2306 BIT_SEL[5].n5 VSS 6.88525f
C2307 BIT_SEL[5].t7 VSS 4.01572f
C2308 BIT_SEL[5].n6 VSS 6.88525f
C2309 BIT_SEL[5].t6 VSS 4.11021f
C2310 a_14320_20781.t0 VSS 1.69351f
C2311 a_14320_20781.t1 VSS 4.30649f
C2312 a_7830_31764.t0 VSS 2.41699f
C2313 a_7830_31764.t1 VSS 3.68301f
C2314 a_7738_11958.t0 VSS 1.47655f
C2315 a_7738_11958.t1 VSS 4.52345f
C2316 BIT_SEL[16].t0 VSS 3.0317f
C2317 BIT_SEL[16].n0 VSS 5.09227f
C2318 BIT_SEL[16].t2 VSS 3.0317f
C2319 BIT_SEL[16].n1 VSS 5.09227f
C2320 BIT_SEL[16].t5 VSS 3.0317f
C2321 BIT_SEL[16].n2 VSS 5.09227f
C2322 BIT_SEL[16].t6 VSS 3.0317f
C2323 BIT_SEL[16].n3 VSS 5.09227f
C2324 BIT_SEL[16].t1 VSS 3.0317f
C2325 BIT_SEL[16].n4 VSS 5.09227f
C2326 BIT_SEL[16].t7 VSS 3.0317f
C2327 BIT_SEL[16].n5 VSS 5.09227f
C2328 BIT_SEL[16].t4 VSS 3.06458f
C2329 BIT_SEL[16].t3 VSS 3.0317f
C2330 BIT_SEL[16].n6 VSS 5.09227f
C2331 a_1340_55763.t0 VSS 3.86539f
C2332 a_1340_55763.t1 VSS 2.23461f
C2333 BIT_SEL[13].t7 VSS 4.14801f
C2334 BIT_SEL[13].n0 VSS 7.33197f
C2335 BIT_SEL[13].t1 VSS 4.14801f
C2336 BIT_SEL[13].n1 VSS 7.33197f
C2337 BIT_SEL[13].t2 VSS 4.14801f
C2338 BIT_SEL[13].n2 VSS 7.33197f
C2339 BIT_SEL[13].t5 VSS 4.14801f
C2340 BIT_SEL[13].n3 VSS 7.33197f
C2341 BIT_SEL[13].t6 VSS 4.14801f
C2342 BIT_SEL[13].n4 VSS 7.33197f
C2343 BIT_SEL[13].t0 VSS 4.14801f
C2344 BIT_SEL[13].n5 VSS 7.33197f
C2345 BIT_SEL[13].t4 VSS 4.14801f
C2346 BIT_SEL[13].n6 VSS 7.33197f
C2347 BIT_SEL[13].t3 VSS 4.41496f
C2348 a_14320_14169.t0 VSS 3.66536f
C2349 a_14320_14169.t1 VSS 2.33464f
C2350 a_20810_6292.t0 VSS 2.33483f
C2351 a_20810_6292.t1 VSS 3.66517f
C2352 BIT_SEL[56].t3 VSS 4.14071f
C2353 BIT_SEL[56].n0 VSS 7.18434f
C2354 BIT_SEL[56].t5 VSS 4.14071f
C2355 BIT_SEL[56].n1 VSS 7.18434f
C2356 BIT_SEL[56].t6 VSS 4.14071f
C2357 BIT_SEL[56].n2 VSS 7.18434f
C2358 BIT_SEL[56].t7 VSS 4.14071f
C2359 BIT_SEL[56].n3 VSS 7.18434f
C2360 BIT_SEL[56].t1 VSS 4.14071f
C2361 BIT_SEL[56].n4 VSS 7.18434f
C2362 BIT_SEL[56].t4 VSS 4.14071f
C2363 BIT_SEL[56].n5 VSS 7.18434f
C2364 BIT_SEL[56].t2 VSS 4.31483f
C2365 BIT_SEL[56].t0 VSS 4.14071f
C2366 BIT_SEL[56].n6 VSS 7.18434f
C2367 a_7830_18908.t0 VSS 4.60993f
C2368 a_7830_18908.t1 VSS 1.39007f
C2369 BIT_SEL[17].t5 VSS 4.07792f
C2370 BIT_SEL[17].n0 VSS 6.88058f
C2371 BIT_SEL[17].t0 VSS 4.07792f
C2372 BIT_SEL[17].n1 VSS 6.88058f
C2373 BIT_SEL[17].t1 VSS 4.07792f
C2374 BIT_SEL[17].n2 VSS 6.88058f
C2375 BIT_SEL[17].t4 VSS 4.07792f
C2376 BIT_SEL[17].n3 VSS 6.88058f
C2377 BIT_SEL[17].t2 VSS 4.07792f
C2378 BIT_SEL[17].n4 VSS 6.88058f
C2379 BIT_SEL[17].t6 VSS 4.07792f
C2380 BIT_SEL[17].n5 VSS 6.88058f
C2381 BIT_SEL[17].t3 VSS 4.07792f
C2382 BIT_SEL[17].n6 VSS 6.88058f
C2383 BIT_SEL[17].t7 VSS 4.12246f
C2384 a_7830_45677.t0 VSS 2.33483f
C2385 a_7830_45677.t1 VSS 3.66517f
C2386 a_7830_16010.t0 VSS 2.41699f
C2387 a_7830_16010.t1 VSS 3.68301f
C2388 a_638_19518.t0 VSS 0.07629f
C2389 a_638_19518.n0 VSS 0.1989f
C2390 a_638_19518.n1 VSS 0.20832f
C2391 a_638_19518.t66 VSS 0.07629f
C2392 a_638_19518.n2 VSS 0.1989f
C2393 a_638_19518.t34 VSS 0.07629f
C2394 a_638_19518.n3 VSS 0.1989f
C2395 a_638_19518.t47 VSS 0.07629f
C2396 a_638_19518.n4 VSS 0.1989f
C2397 a_638_19518.t60 VSS 0.07629f
C2398 a_638_19518.n5 VSS 0.1989f
C2399 a_638_19518.t15 VSS 0.07629f
C2400 a_638_19518.n6 VSS 0.1989f
C2401 a_638_19518.t61 VSS 0.07629f
C2402 a_638_19518.n7 VSS 0.1989f
C2403 a_638_19518.t40 VSS 0.07629f
C2404 a_638_19518.n8 VSS 0.22891f
C2405 a_638_19518.t51 VSS 0.07629f
C2406 a_638_19518.n9 VSS 0.22891f
C2407 a_638_19518.t26 VSS 0.07629f
C2408 a_638_19518.n10 VSS 0.1989f
C2409 a_638_19518.t6 VSS 0.07629f
C2410 a_638_19518.n11 VSS 0.1989f
C2411 a_638_19518.t29 VSS 0.07629f
C2412 a_638_19518.n12 VSS 0.1989f
C2413 a_638_19518.t1 VSS 0.07629f
C2414 a_638_19518.n13 VSS 0.1989f
C2415 a_638_19518.t45 VSS 0.07629f
C2416 a_638_19518.n14 VSS 0.1989f
C2417 a_638_19518.t16 VSS 0.07629f
C2418 a_638_19518.n15 VSS 0.22891f
C2419 a_638_19518.t17 VSS 0.07629f
C2420 a_638_19518.n16 VSS 0.22891f
C2421 a_638_19518.t35 VSS 0.07629f
C2422 a_638_19518.n17 VSS 0.1989f
C2423 a_638_19518.t21 VSS 0.07629f
C2424 a_638_19518.n18 VSS 0.1989f
C2425 a_638_19518.t63 VSS 0.07629f
C2426 a_638_19518.n19 VSS 0.1989f
C2427 a_638_19518.t39 VSS 0.07629f
C2428 a_638_19518.n20 VSS 0.1989f
C2429 a_638_19518.t54 VSS 0.07629f
C2430 a_638_19518.n21 VSS 0.1989f
C2431 a_638_19518.t56 VSS 0.07629f
C2432 a_638_19518.n22 VSS 0.1989f
C2433 a_638_19518.t68 VSS 0.07629f
C2434 a_638_19518.n23 VSS 0.22891f
C2435 a_638_19518.t9 VSS 0.07629f
C2436 a_638_19518.n24 VSS 0.22891f
C2437 a_638_19518.t41 VSS 0.07629f
C2438 a_638_19518.n25 VSS 0.1989f
C2439 a_638_19518.t19 VSS 0.07629f
C2440 a_638_19518.n26 VSS 0.1989f
C2441 a_638_19518.t65 VSS 0.07629f
C2442 a_638_19518.n27 VSS 0.1989f
C2443 a_638_19518.t25 VSS 0.07629f
C2444 a_638_19518.n28 VSS 0.1989f
C2445 a_638_19518.t38 VSS 0.07629f
C2446 a_638_19518.n29 VSS 0.1989f
C2447 a_638_19518.t36 VSS 0.07629f
C2448 a_638_19518.n30 VSS 0.1989f
C2449 a_638_19518.t12 VSS 0.07629f
C2450 a_638_19518.n31 VSS 0.21781f
C2451 a_638_19518.t43 VSS 0.07629f
C2452 a_638_19518.n32 VSS 0.22837f
C2453 a_638_19518.t24 VSS 0.01725f
C2454 a_638_19518.t52 VSS 0.50628f
C2455 a_638_19518.n33 VSS -0.31292f
C2456 a_638_19518.n34 VSS 0.10989f
C2457 a_638_19518.n35 VSS 0.07801f
C2458 a_638_19518.n36 VSS 0.2494f
C2459 a_638_19518.t23 VSS 0.07629f
C2460 a_638_19518.n37 VSS 0.20508f
C2461 a_638_19518.t44 VSS 0.07629f
C2462 a_638_19518.n38 VSS 0.20508f
C2463 a_638_19518.t18 VSS 0.07629f
C2464 a_638_19518.n39 VSS 0.20508f
C2465 a_638_19518.t8 VSS 0.07629f
C2466 a_638_19518.n40 VSS 0.20508f
C2467 a_638_19518.t33 VSS 0.07629f
C2468 a_638_19518.n41 VSS 0.20508f
C2469 a_638_19518.t64 VSS 0.07629f
C2470 a_638_19518.n42 VSS 0.20508f
C2471 a_638_19518.t37 VSS 0.07629f
C2472 a_638_19518.n43 VSS 0.2351f
C2473 a_638_19518.t48 VSS 0.07629f
C2474 a_638_19518.n44 VSS 0.2351f
C2475 a_638_19518.t50 VSS 0.07629f
C2476 a_638_19518.n45 VSS 0.20508f
C2477 a_638_19518.t55 VSS 0.07629f
C2478 a_638_19518.n46 VSS 0.20508f
C2479 a_638_19518.t28 VSS 0.07629f
C2480 a_638_19518.n47 VSS 0.20508f
C2481 a_638_19518.t5 VSS 0.07629f
C2482 a_638_19518.n48 VSS 0.20508f
C2483 a_638_19518.t13 VSS 0.07629f
C2484 a_638_19518.n49 VSS 0.20508f
C2485 a_638_19518.t20 VSS 0.07629f
C2486 a_638_19518.n50 VSS 0.20508f
C2487 a_638_19518.t42 VSS 0.07629f
C2488 a_638_19518.n51 VSS 0.2351f
C2489 a_638_19518.t10 VSS 0.07629f
C2490 a_638_19518.n52 VSS 0.2351f
C2491 a_638_19518.t67 VSS 0.07629f
C2492 a_638_19518.n53 VSS 0.20508f
C2493 a_638_19518.t31 VSS 0.07629f
C2494 a_638_19518.n54 VSS 0.20508f
C2495 a_638_19518.t4 VSS 0.07629f
C2496 a_638_19518.n55 VSS 0.20508f
C2497 a_638_19518.t22 VSS 0.07629f
C2498 a_638_19518.n56 VSS 0.20508f
C2499 a_638_19518.t32 VSS 0.07629f
C2500 a_638_19518.n57 VSS 0.20508f
C2501 a_638_19518.t46 VSS 0.07629f
C2502 a_638_19518.n58 VSS 0.20508f
C2503 a_638_19518.t7 VSS 0.07629f
C2504 a_638_19518.n59 VSS 0.2351f
C2505 a_638_19518.t30 VSS 0.07629f
C2506 a_638_19518.n60 VSS 0.2351f
C2507 a_638_19518.t3 VSS 0.07629f
C2508 a_638_19518.n61 VSS 0.20508f
C2509 a_638_19518.t27 VSS 0.07629f
C2510 a_638_19518.n62 VSS 0.20508f
C2511 a_638_19518.t2 VSS 0.07629f
C2512 a_638_19518.n63 VSS 0.20508f
C2513 a_638_19518.t53 VSS 0.07629f
C2514 a_638_19518.n64 VSS 0.20508f
C2515 a_638_19518.t62 VSS 0.07629f
C2516 a_638_19518.n65 VSS 0.20508f
C2517 a_638_19518.t14 VSS 0.07629f
C2518 a_638_19518.n66 VSS 0.20508f
C2519 a_638_19518.t49 VSS 0.07629f
C2520 a_638_19518.n67 VSS 0.19068f
C2521 a_638_19518.t11 VSS 0.07629f
C2522 a_638_19518.t59 VSS 0.21301f
C2523 a_638_19518.t57 VSS 0.21301f
C2524 a_638_19518.n68 VSS 0.42602f
C2525 a_638_19518.n69 VSS -0.52759f
C2526 a_638_19518.n70 VSS 0.15155f
C2527 a_638_19518.n71 VSS 0.13888f
C2528 a_638_19518.t58 VSS 0.50628f
C2529 a_638_19518.n72 VSS 0.82359f
C2530 a_7830_29923.t0 VSS 2.33483f
C2531 a_7830_29923.t1 VSS 3.66517f
C2532 a_14320_12904.t0 VSS 1.69351f
C2533 a_14320_12904.t1 VSS 4.30649f
C2534 BIT_SEL[34].t2 VSS 4.05315f
C2535 BIT_SEL[34].n0 VSS 6.86345f
C2536 BIT_SEL[34].t0 VSS 4.05315f
C2537 BIT_SEL[34].n1 VSS 6.86345f
C2538 BIT_SEL[34].t6 VSS 4.05315f
C2539 BIT_SEL[34].n2 VSS 6.86345f
C2540 BIT_SEL[34].t3 VSS 4.05315f
C2541 BIT_SEL[34].n3 VSS 6.86345f
C2542 BIT_SEL[34].t4 VSS 4.05315f
C2543 BIT_SEL[34].n4 VSS 6.86345f
C2544 BIT_SEL[34].t5 VSS 4.05315f
C2545 BIT_SEL[34].n5 VSS 6.86345f
C2546 BIT_SEL[34].t7 VSS 4.05315f
C2547 BIT_SEL[34].n6 VSS 6.86345f
C2548 BIT_SEL[34].t1 VSS 4.12109f
C2549 a_14320_40906.t0 VSS 4.20807f
C2550 a_14320_40906.t1 VSS 1.79193f
C2551 a_20810_58293.t0 VSS 4.60993f
C2552 a_20810_58293.t1 VSS 1.39007f
C2553 a_14228_4081.t0 VSS 1.47655f
C2554 a_14228_4081.t1 VSS 4.52345f
C2555 a_20810_57556.t0 VSS 1.6826f
C2556 a_20810_57556.t1 VSS 4.3174f
C2557 a_20810_21149.t0 VSS 4.27849f
C2558 a_20810_21149.t1 VSS 1.72151f
C2559 a_7830_44780.t0 VSS 4.27849f
C2560 a_7830_44780.t1 VSS 1.72151f
C2561 BIT_SEL[20].t6 VSS 4.02347f
C2562 BIT_SEL[20].n0 VSS 6.87043f
C2563 BIT_SEL[20].t5 VSS 4.02347f
C2564 BIT_SEL[20].n1 VSS 6.87043f
C2565 BIT_SEL[20].t3 VSS 4.02347f
C2566 BIT_SEL[20].n2 VSS 6.87043f
C2567 BIT_SEL[20].t7 VSS 4.02347f
C2568 BIT_SEL[20].n3 VSS 6.87043f
C2569 BIT_SEL[20].t1 VSS 4.02347f
C2570 BIT_SEL[20].n4 VSS 6.87043f
C2571 BIT_SEL[20].t0 VSS 4.02347f
C2572 BIT_SEL[20].n5 VSS 6.87043f
C2573 BIT_SEL[20].t2 VSS 4.02347f
C2574 BIT_SEL[20].n6 VSS 6.87043f
C2575 BIT_SEL[20].t4 VSS 4.11755f
C2576 a_7830_29555.t0 VSS 1.745f
C2577 a_7830_29555.t1 VSS 4.255f
C2578 BIT_SEL[22].t7 VSS 4.07324f
C2579 BIT_SEL[22].n0 VSS 7.01202f
C2580 BIT_SEL[22].t2 VSS 4.07324f
C2581 BIT_SEL[22].n1 VSS 7.01202f
C2582 BIT_SEL[22].t4 VSS 4.07324f
C2583 BIT_SEL[22].n2 VSS 7.01202f
C2584 BIT_SEL[22].t0 VSS 4.07324f
C2585 BIT_SEL[22].n3 VSS 7.01202f
C2586 BIT_SEL[22].t1 VSS 4.07324f
C2587 BIT_SEL[22].n4 VSS 7.01202f
C2588 BIT_SEL[22].t3 VSS 4.07324f
C2589 BIT_SEL[22].n5 VSS 7.01202f
C2590 BIT_SEL[22].t5 VSS 4.07324f
C2591 BIT_SEL[22].n6 VSS 7.01202f
C2592 BIT_SEL[22].t6 VSS 4.21129f
C2593 a_14320_61431.t0 VSS 2.33483f
C2594 a_14320_61431.t1 VSS 3.66517f
C2595 a_7830_14169.t0 VSS 2.33483f
C2596 a_7830_14169.t1 VSS 3.66517f
C2597 a_14320_25152.t0 VSS 4.20807f
C2598 a_14320_25152.t1 VSS 1.79193f
C2599 a_20810_42539.t0 VSS 1.39007f
C2600 a_20810_42539.t1 VSS 4.60993f
C2601 a_1340_23887.t0 VSS 3.68292f
C2602 a_1340_23887.t1 VSS 2.41708f
C2603 BIT_SEL[15].t2 VSS 3.1518f
C2604 BIT_SEL[15].n0 VSS 5.61038f
C2605 BIT_SEL[15].t0 VSS 3.1518f
C2606 BIT_SEL[15].n1 VSS 5.61038f
C2607 BIT_SEL[15].t3 VSS 3.1518f
C2608 BIT_SEL[15].n2 VSS 5.61038f
C2609 BIT_SEL[15].t6 VSS 3.1518f
C2610 BIT_SEL[15].n3 VSS 5.61038f
C2611 BIT_SEL[15].t7 VSS 3.1518f
C2612 BIT_SEL[15].n4 VSS 5.61038f
C2613 BIT_SEL[15].t1 VSS 3.1518f
C2614 BIT_SEL[15].n5 VSS 5.61038f
C2615 BIT_SEL[15].t4 VSS 3.1518f
C2616 BIT_SEL[15].n6 VSS 5.61038f
C2617 BIT_SEL[15].t5 VSS 3.38636f
C2618 COL_PROG_N[0].t3 VSS 1.10931f
C2619 COL_PROG_N[0].n0 VSS 0.38563f
C2620 COL_PROG_N[0].t0 VSS 1.10931f
C2621 COL_PROG_N[0].n1 VSS 0.39369f
C2622 COL_PROG_N[0].t1 VSS 1.10931f
C2623 COL_PROG_N[0].n2 VSS 0.77937f
C2624 COL_PROG_N[0].t2 VSS 1.10971f
C2625 a_20718_19835.t0 VSS 1.47655f
C2626 a_20718_19835.t1 VSS 4.52345f
C2627 BIT_SEL[48].t1 VSS 3.45483f
C2628 BIT_SEL[48].n0 VSS 5.80298f
C2629 BIT_SEL[48].t6 VSS 3.45483f
C2630 BIT_SEL[48].n1 VSS 5.80298f
C2631 BIT_SEL[48].t0 VSS 3.45483f
C2632 BIT_SEL[48].n2 VSS 5.80298f
C2633 BIT_SEL[48].t3 VSS 3.45483f
C2634 BIT_SEL[48].n3 VSS 5.80298f
C2635 BIT_SEL[48].t4 VSS 3.45483f
C2636 BIT_SEL[48].n4 VSS 5.80298f
C2637 BIT_SEL[48].t7 VSS 3.45483f
C2638 BIT_SEL[48].n5 VSS 5.80298f
C2639 BIT_SEL[48].t5 VSS 3.45483f
C2640 BIT_SEL[48].n6 VSS 5.80298f
C2641 BIT_SEL[48].t2 VSS 3.49229f
C2642 a_14320_45677.t0 VSS 3.66536f
C2643 a_14320_45677.t1 VSS 2.33464f
C2644 BIT_SEL[40].t6 VSS 4.14071f
C2645 BIT_SEL[40].n0 VSS 7.18434f
C2646 BIT_SEL[40].t2 VSS 4.14071f
C2647 BIT_SEL[40].n1 VSS 7.18434f
C2648 BIT_SEL[40].t4 VSS 4.14071f
C2649 BIT_SEL[40].n2 VSS 7.18434f
C2650 BIT_SEL[40].t5 VSS 4.14071f
C2651 BIT_SEL[40].n3 VSS 7.18434f
C2652 BIT_SEL[40].t7 VSS 4.14071f
C2653 BIT_SEL[40].n4 VSS 7.18434f
C2654 BIT_SEL[40].t0 VSS 4.14071f
C2655 BIT_SEL[40].n5 VSS 7.18434f
C2656 BIT_SEL[40].t3 VSS 4.14071f
C2657 BIT_SEL[40].n6 VSS 7.18434f
C2658 BIT_SEL[40].t1 VSS 4.31483f
C2659 a_1340_55395.t0 VSS 2.41699f
C2660 a_1340_55395.t1 VSS 3.68301f
C2661 a_14320_1521.t0 VSS 4.20807f
C2662 a_14320_1521.t1 VSS 1.79193f
C2663 a_20810_26785.t0 VSS 1.39007f
C2664 a_20810_26785.t1 VSS 4.60993f
C2665 a_638_51026.t0 VSS 0.07629f
C2666 a_638_51026.n0 VSS 0.20508f
C2667 a_638_51026.n1 VSS 0.07801f
C2668 a_638_51026.n2 VSS 0.2494f
C2669 a_638_51026.t59 VSS 0.07629f
C2670 a_638_51026.n3 VSS 0.20508f
C2671 a_638_51026.t3 VSS 0.07629f
C2672 a_638_51026.n4 VSS 0.20508f
C2673 a_638_51026.t5 VSS 0.07629f
C2674 a_638_51026.n5 VSS 0.20508f
C2675 a_638_51026.t58 VSS 0.07629f
C2676 a_638_51026.n6 VSS 0.20508f
C2677 a_638_51026.t22 VSS 0.07629f
C2678 a_638_51026.n7 VSS 0.20508f
C2679 a_638_51026.t10 VSS 0.07629f
C2680 a_638_51026.n8 VSS 0.20508f
C2681 a_638_51026.t20 VSS 0.07629f
C2682 a_638_51026.n9 VSS 0.2351f
C2683 a_638_51026.t27 VSS 0.07629f
C2684 a_638_51026.n10 VSS 0.2351f
C2685 a_638_51026.t40 VSS 0.07629f
C2686 a_638_51026.n11 VSS 0.20508f
C2687 a_638_51026.t55 VSS 0.07629f
C2688 a_638_51026.n12 VSS 0.20508f
C2689 a_638_51026.t52 VSS 0.07629f
C2690 a_638_51026.n13 VSS 0.20508f
C2691 a_638_51026.t42 VSS 0.07629f
C2692 a_638_51026.n14 VSS 0.20508f
C2693 a_638_51026.t6 VSS 0.07629f
C2694 a_638_51026.n15 VSS 0.20508f
C2695 a_638_51026.t66 VSS 0.07629f
C2696 a_638_51026.n16 VSS 0.20508f
C2697 a_638_51026.t67 VSS 0.07629f
C2698 a_638_51026.n17 VSS 0.2351f
C2699 a_638_51026.t32 VSS 0.07629f
C2700 a_638_51026.n18 VSS 0.2351f
C2701 a_638_51026.t36 VSS 0.07629f
C2702 a_638_51026.n19 VSS 0.20508f
C2703 a_638_51026.t56 VSS 0.07629f
C2704 a_638_51026.n20 VSS 0.20508f
C2705 a_638_51026.t2 VSS 0.07629f
C2706 a_638_51026.n21 VSS 0.20508f
C2707 a_638_51026.t28 VSS 0.07629f
C2708 a_638_51026.n22 VSS 0.20508f
C2709 a_638_51026.t45 VSS 0.07629f
C2710 a_638_51026.n23 VSS 0.20508f
C2711 a_638_51026.t65 VSS 0.07629f
C2712 a_638_51026.n24 VSS 0.2351f
C2713 a_638_51026.t26 VSS 0.07629f
C2714 a_638_51026.n25 VSS 0.2351f
C2715 a_638_51026.t50 VSS 0.07629f
C2716 a_638_51026.n26 VSS 0.20508f
C2717 a_638_51026.t54 VSS 0.07629f
C2718 a_638_51026.n27 VSS 0.20508f
C2719 a_638_51026.t29 VSS 0.07629f
C2720 a_638_51026.n28 VSS 0.20508f
C2721 a_638_51026.t57 VSS 0.07629f
C2722 a_638_51026.n29 VSS 0.20508f
C2723 a_638_51026.t46 VSS 0.07629f
C2724 a_638_51026.n30 VSS 0.20508f
C2725 a_638_51026.t41 VSS 0.07629f
C2726 a_638_51026.n31 VSS 0.20508f
C2727 a_638_51026.t39 VSS 0.07629f
C2728 a_638_51026.n32 VSS 0.19068f
C2729 a_638_51026.t64 VSS 0.07629f
C2730 a_638_51026.n33 VSS 0.13888f
C2731 a_638_51026.n34 VSS 0.22837f
C2732 a_638_51026.t31 VSS 0.01725f
C2733 a_638_51026.n35 VSS 0.20832f
C2734 a_638_51026.t43 VSS 0.07629f
C2735 a_638_51026.n36 VSS 0.1989f
C2736 a_638_51026.t1 VSS 0.07629f
C2737 a_638_51026.n37 VSS 0.1989f
C2738 a_638_51026.t44 VSS 0.07629f
C2739 a_638_51026.n38 VSS 0.1989f
C2740 a_638_51026.t34 VSS 0.07629f
C2741 a_638_51026.n39 VSS 0.1989f
C2742 a_638_51026.t9 VSS 0.07629f
C2743 a_638_51026.n40 VSS 0.1989f
C2744 a_638_51026.t68 VSS 0.07629f
C2745 a_638_51026.n41 VSS 0.1989f
C2746 a_638_51026.t12 VSS 0.07629f
C2747 a_638_51026.n42 VSS 0.22891f
C2748 a_638_51026.t53 VSS 0.07629f
C2749 a_638_51026.n43 VSS 0.22891f
C2750 a_638_51026.t21 VSS 0.07629f
C2751 a_638_51026.n44 VSS 0.1989f
C2752 a_638_51026.t18 VSS 0.07629f
C2753 a_638_51026.n45 VSS 0.1989f
C2754 a_638_51026.t15 VSS 0.07629f
C2755 a_638_51026.n46 VSS 0.1989f
C2756 a_638_51026.t30 VSS 0.07629f
C2757 a_638_51026.n47 VSS 0.1989f
C2758 a_638_51026.t48 VSS 0.07629f
C2759 a_638_51026.n48 VSS 0.1989f
C2760 a_638_51026.t49 VSS 0.07629f
C2761 a_638_51026.n49 VSS 0.1989f
C2762 a_638_51026.t7 VSS 0.07629f
C2763 a_638_51026.n50 VSS 0.22891f
C2764 a_638_51026.t25 VSS 0.07629f
C2765 a_638_51026.n51 VSS 0.22891f
C2766 a_638_51026.t33 VSS 0.07629f
C2767 a_638_51026.n52 VSS 0.1989f
C2768 a_638_51026.t17 VSS 0.07629f
C2769 a_638_51026.n53 VSS 0.1989f
C2770 a_638_51026.t47 VSS 0.07629f
C2771 a_638_51026.n54 VSS 0.1989f
C2772 a_638_51026.t14 VSS 0.07629f
C2773 a_638_51026.n55 VSS 0.1989f
C2774 a_638_51026.t16 VSS 0.07629f
C2775 a_638_51026.n56 VSS 0.1989f
C2776 a_638_51026.t4 VSS 0.07629f
C2777 a_638_51026.n57 VSS 0.1989f
C2778 a_638_51026.t51 VSS 0.07629f
C2779 a_638_51026.n58 VSS 0.22891f
C2780 a_638_51026.t24 VSS 0.07629f
C2781 a_638_51026.n59 VSS 0.22891f
C2782 a_638_51026.t23 VSS 0.07629f
C2783 a_638_51026.n60 VSS 0.1989f
C2784 a_638_51026.t8 VSS 0.07629f
C2785 a_638_51026.n61 VSS 0.1989f
C2786 a_638_51026.t37 VSS 0.07629f
C2787 a_638_51026.n62 VSS 0.1989f
C2788 a_638_51026.t19 VSS 0.07629f
C2789 a_638_51026.n63 VSS 0.1989f
C2790 a_638_51026.t38 VSS 0.07629f
C2791 a_638_51026.n64 VSS 0.1989f
C2792 a_638_51026.t13 VSS 0.07629f
C2793 a_638_51026.n65 VSS 0.1989f
C2794 a_638_51026.t35 VSS 0.07629f
C2795 a_638_51026.n66 VSS 0.21781f
C2796 a_638_51026.t11 VSS 0.07629f
C2797 a_638_51026.t61 VSS 0.50628f
C2798 a_638_51026.n67 VSS 0.82359f
C2799 a_638_51026.n68 VSS 0.15155f
C2800 a_638_51026.t62 VSS 0.21301f
C2801 a_638_51026.t63 VSS 0.21301f
C2802 a_638_51026.n69 VSS 0.42602f
C2803 a_638_51026.n70 VSS -0.52759f
C2804 a_638_51026.n71 VSS 0.10989f
C2805 a_638_51026.t60 VSS 0.50628f
C2806 a_638_51026.n72 VSS -0.31292f
C2807 a_7830_52657.t0 VSS 4.27849f
C2808 a_7830_52657.t1 VSS 1.72151f
C2809 a_1340_23311.t0 VSS 3.74618f
C2810 a_1340_23311.t1 VSS 2.35382f
C2811 BIT_SEL[14].t6 VSS 4.1517f
C2812 BIT_SEL[14].n0 VSS 7.36453f
C2813 BIT_SEL[14].t0 VSS 4.1517f
C2814 BIT_SEL[14].n1 VSS 7.36453f
C2815 BIT_SEL[14].t2 VSS 4.1517f
C2816 BIT_SEL[14].n2 VSS 7.36453f
C2817 BIT_SEL[14].t5 VSS 4.1517f
C2818 BIT_SEL[14].n3 VSS 7.36453f
C2819 BIT_SEL[14].t7 VSS 4.1517f
C2820 BIT_SEL[14].n4 VSS 7.36453f
C2821 BIT_SEL[14].t4 VSS 4.1517f
C2822 BIT_SEL[14].n5 VSS 7.36453f
C2823 BIT_SEL[14].t1 VSS 4.45988f
C2824 BIT_SEL[14].t3 VSS 4.1517f
C2825 BIT_SEL[14].n6 VSS 7.36453f
C2826 a_14320_9398.t0 VSS 1.79192f
C2827 a_14320_9398.t1 VSS 4.20808f
C2828 a_1340_57028.t0 VSS 1.69725f
C2829 a_1340_57028.t1 VSS 4.30275f
C2830 BIT_SEL[62].t0 VSS 4.1517f
C2831 BIT_SEL[62].n0 VSS 7.36453f
C2832 BIT_SEL[62].t3 VSS 4.1517f
C2833 BIT_SEL[62].n1 VSS 7.36453f
C2834 BIT_SEL[62].t5 VSS 4.1517f
C2835 BIT_SEL[62].n2 VSS 7.36453f
C2836 BIT_SEL[62].t7 VSS 4.1517f
C2837 BIT_SEL[62].n3 VSS 7.36453f
C2838 BIT_SEL[62].t2 VSS 4.1517f
C2839 BIT_SEL[62].n4 VSS 7.36453f
C2840 BIT_SEL[62].t4 VSS 4.1517f
C2841 BIT_SEL[62].n5 VSS 7.36453f
C2842 BIT_SEL[62].t1 VSS 4.1517f
C2843 BIT_SEL[62].n6 VSS 7.36453f
C2844 BIT_SEL[62].t6 VSS 4.45988f
C2845 a_1340_42539.t0 VSS 1.39007f
C2846 a_1340_42539.t1 VSS 4.60993f
C2847 a_14320_45309.t0 VSS 4.25498f
C2848 a_14320_45309.t1 VSS 1.74502f
C2849 a_20810_26417.t0 VSS 4.34773f
C2850 a_20810_26417.t1 VSS 1.65227f
C2851 BIT_SEL[51].t2 VSS 4.04507f
C2852 BIT_SEL[51].n0 VSS 6.87869f
C2853 BIT_SEL[51].t6 VSS 4.04507f
C2854 BIT_SEL[51].n1 VSS 6.87869f
C2855 BIT_SEL[51].t0 VSS 4.04507f
C2856 BIT_SEL[51].n2 VSS 6.87869f
C2857 BIT_SEL[51].t1 VSS 4.04507f
C2858 BIT_SEL[51].n3 VSS 6.87869f
C2859 BIT_SEL[51].t3 VSS 4.04507f
C2860 BIT_SEL[51].n4 VSS 6.87869f
C2861 BIT_SEL[51].t4 VSS 4.04507f
C2862 BIT_SEL[51].n5 VSS 6.87869f
C2863 BIT_SEL[51].t5 VSS 4.04507f
C2864 BIT_SEL[51].n6 VSS 6.87869f
C2865 BIT_SEL[51].t7 VSS 4.1133f
C2866 a_1340_1889.t0 VSS 4.30261f
C2867 a_1340_1889.t1 VSS 1.69739f
C2868 BIT_SEL[7].t7 VSS 4.06977f
C2869 BIT_SEL[7].n0 VSS 7.03381f
C2870 BIT_SEL[7].t2 VSS 4.06977f
C2871 BIT_SEL[7].n1 VSS 7.03381f
C2872 BIT_SEL[7].t4 VSS 4.06977f
C2873 BIT_SEL[7].n2 VSS 7.03381f
C2874 BIT_SEL[7].t5 VSS 4.06977f
C2875 BIT_SEL[7].n3 VSS 7.03381f
C2876 BIT_SEL[7].t6 VSS 4.06977f
C2877 BIT_SEL[7].n4 VSS 7.03381f
C2878 BIT_SEL[7].t3 VSS 4.06977f
C2879 BIT_SEL[7].n5 VSS 7.03381f
C2880 BIT_SEL[7].t1 VSS 4.06977f
C2881 BIT_SEL[7].n6 VSS 7.03381f
C2882 BIT_SEL[7].t0 VSS 4.20835f
C2883 a_20810_38168.t0 VSS 4.08932f
C2884 a_20810_38168.t1 VSS 1.91068f
C2885 BIT_SEL[58].t1 VSS 4.02969f
C2886 BIT_SEL[58].n0 VSS 7.04511f
C2887 BIT_SEL[58].t3 VSS 4.02969f
C2888 BIT_SEL[58].n1 VSS 7.04511f
C2889 BIT_SEL[58].t6 VSS 4.02969f
C2890 BIT_SEL[58].n2 VSS 7.04511f
C2891 BIT_SEL[58].t0 VSS 4.02969f
C2892 BIT_SEL[58].n3 VSS 7.04511f
C2893 BIT_SEL[58].t2 VSS 4.02969f
C2894 BIT_SEL[58].n4 VSS 7.04511f
C2895 BIT_SEL[58].t4 VSS 4.02969f
C2896 BIT_SEL[58].n5 VSS 7.04511f
C2897 BIT_SEL[58].t5 VSS 4.2344f
C2898 BIT_SEL[58].t7 VSS 4.02969f
C2899 BIT_SEL[58].n6 VSS 7.04511f
C2900 a_20810_55763.t0 VSS 3.86539f
C2901 a_20810_55763.t1 VSS 2.23461f
C2902 a_20810_7189.t0 VSS 2.2362f
C2903 a_20810_7189.t1 VSS 4.0638f
C2904 BIT_SEL[60].t6 VSS 4.12331f
C2905 BIT_SEL[60].n0 VSS 7.26213f
C2906 BIT_SEL[60].t7 VSS 4.12331f
C2907 BIT_SEL[60].n1 VSS 7.26213f
C2908 BIT_SEL[60].t3 VSS 4.12331f
C2909 BIT_SEL[60].n2 VSS 7.26213f
C2910 BIT_SEL[60].t1 VSS 4.12331f
C2911 BIT_SEL[60].n3 VSS 7.26213f
C2912 BIT_SEL[60].t4 VSS 4.12331f
C2913 BIT_SEL[60].n4 VSS 7.26213f
C2914 BIT_SEL[60].t2 VSS 4.12331f
C2915 BIT_SEL[60].n5 VSS 7.26213f
C2916 BIT_SEL[60].t5 VSS 4.3879f
C2917 BIT_SEL[60].t0 VSS 4.12331f
C2918 BIT_SEL[60].n6 VSS 7.26213f
C2919 BIT_SEL[57].t4 VSS 4.14534f
C2920 BIT_SEL[57].n0 VSS 7.22001f
C2921 BIT_SEL[57].t7 VSS 4.14534f
C2922 BIT_SEL[57].n1 VSS 7.22001f
C2923 BIT_SEL[57].t2 VSS 4.14534f
C2924 BIT_SEL[57].n2 VSS 7.22001f
C2925 BIT_SEL[57].t0 VSS 4.14534f
C2926 BIT_SEL[57].n3 VSS 7.22001f
C2927 BIT_SEL[57].t3 VSS 4.14534f
C2928 BIT_SEL[57].n4 VSS 7.22001f
C2929 BIT_SEL[57].t6 VSS 4.14534f
C2930 BIT_SEL[57].n5 VSS 7.22001f
C2931 BIT_SEL[57].t1 VSS 4.14534f
C2932 BIT_SEL[57].n6 VSS 7.22001f
C2933 BIT_SEL[57].t5 VSS 4.32038f
C2934 a_20810_40906.t0 VSS 1.79192f
C2935 a_20810_40906.t1 VSS 4.20808f
C2936 a_1340_7557.t0 VSS 2.354f
C2937 a_1340_7557.t1 VSS 3.746f
C2938 a_1340_26785.t0 VSS 4.60993f
C2939 a_1340_26785.t1 VSS 1.39007f
C2940 a_1248_59220.t0 VSS 4.52345f
C2941 a_1248_59220.t1 VSS 1.47655f
C2942 a_20810_52657.t0 VSS 1.7215f
C2943 a_20810_52657.t1 VSS 4.2785f
C2944 a_20810_37432.t0 VSS 4.25498f
C2945 a_20810_37432.t1 VSS 1.74502f
C2946 BIT_SEL[54].t1 VSS 4.07324f
C2947 BIT_SEL[54].n0 VSS 7.01202f
C2948 BIT_SEL[54].t3 VSS 4.07324f
C2949 BIT_SEL[54].n1 VSS 7.01202f
C2950 BIT_SEL[54].t7 VSS 4.07324f
C2951 BIT_SEL[54].n2 VSS 7.01202f
C2952 BIT_SEL[54].t0 VSS 4.07324f
C2953 BIT_SEL[54].n3 VSS 7.01202f
C2954 BIT_SEL[54].t2 VSS 4.07324f
C2955 BIT_SEL[54].n4 VSS 7.01202f
C2956 BIT_SEL[54].t4 VSS 4.07324f
C2957 BIT_SEL[54].n5 VSS 7.01202f
C2958 BIT_SEL[54].t5 VSS 4.21129f
C2959 BIT_SEL[54].t6 VSS 4.07324f
C2960 BIT_SEL[54].n6 VSS 7.01202f
C2961 a_14320_62328.t0 VSS 4.06398f
C2962 a_14320_62328.t1 VSS 2.23602f
C2963 a_638_3764.t0 VSS 0.07629f
C2964 a_638_3764.n0 VSS 0.22891f
C2965 a_638_3764.n1 VSS 0.20832f
C2966 a_638_3764.t64 VSS 0.07629f
C2967 a_638_3764.n2 VSS 0.1989f
C2968 a_638_3764.t32 VSS 0.07629f
C2969 a_638_3764.n3 VSS 0.1989f
C2970 a_638_3764.t23 VSS 0.07629f
C2971 a_638_3764.n4 VSS 0.1989f
C2972 a_638_3764.t19 VSS 0.07629f
C2973 a_638_3764.n5 VSS 0.1989f
C2974 a_638_3764.t38 VSS 0.07629f
C2975 a_638_3764.n6 VSS 0.1989f
C2976 a_638_3764.t42 VSS 0.07629f
C2977 a_638_3764.n7 VSS 0.1989f
C2978 a_638_3764.t55 VSS 0.07629f
C2979 a_638_3764.n8 VSS 0.22891f
C2980 a_638_3764.t28 VSS 0.07629f
C2981 a_638_3764.n9 VSS 0.22891f
C2982 a_638_3764.t61 VSS 0.07629f
C2983 a_638_3764.n10 VSS 0.1989f
C2984 a_638_3764.t35 VSS 0.07629f
C2985 a_638_3764.n11 VSS 0.1989f
C2986 a_638_3764.t26 VSS 0.07629f
C2987 a_638_3764.n12 VSS 0.1989f
C2988 a_638_3764.t41 VSS 0.07629f
C2989 a_638_3764.n13 VSS 0.1989f
C2990 a_638_3764.t16 VSS 0.07629f
C2991 a_638_3764.n14 VSS 0.1989f
C2992 a_638_3764.t11 VSS 0.07629f
C2993 a_638_3764.n15 VSS 0.1989f
C2994 a_638_3764.t68 VSS 0.07629f
C2995 a_638_3764.n16 VSS 0.22891f
C2996 a_638_3764.t15 VSS 0.07629f
C2997 a_638_3764.n17 VSS 0.1989f
C2998 a_638_3764.t53 VSS 0.07629f
C2999 a_638_3764.n18 VSS 0.1989f
C3000 a_638_3764.t62 VSS 0.07629f
C3001 a_638_3764.n19 VSS 0.1989f
C3002 a_638_3764.t18 VSS 0.07629f
C3003 a_638_3764.n20 VSS 0.1989f
C3004 a_638_3764.t51 VSS 0.07629f
C3005 a_638_3764.n21 VSS 0.1989f
C3006 a_638_3764.t31 VSS 0.07629f
C3007 a_638_3764.n22 VSS 0.1989f
C3008 a_638_3764.t58 VSS 0.07629f
C3009 a_638_3764.n23 VSS 0.22891f
C3010 a_638_3764.t2 VSS 0.07629f
C3011 a_638_3764.n24 VSS 0.22891f
C3012 a_638_3764.t54 VSS 0.07629f
C3013 a_638_3764.n25 VSS 0.1989f
C3014 a_638_3764.t30 VSS 0.07629f
C3015 a_638_3764.n26 VSS 0.1989f
C3016 a_638_3764.t59 VSS 0.07629f
C3017 a_638_3764.n27 VSS 0.1989f
C3018 a_638_3764.t1 VSS 0.07629f
C3019 a_638_3764.n28 VSS 0.1989f
C3020 a_638_3764.t52 VSS 0.07629f
C3021 a_638_3764.n29 VSS 0.1989f
C3022 a_638_3764.t14 VSS 0.07629f
C3023 a_638_3764.n30 VSS 0.1989f
C3024 a_638_3764.t4 VSS 0.07629f
C3025 a_638_3764.n31 VSS 0.21781f
C3026 a_638_3764.t57 VSS 0.07629f
C3027 a_638_3764.n32 VSS 0.22837f
C3028 a_638_3764.t33 VSS 0.01725f
C3029 a_638_3764.t5 VSS 0.50628f
C3030 a_638_3764.n33 VSS -0.31292f
C3031 a_638_3764.n34 VSS 0.10989f
C3032 a_638_3764.n35 VSS 0.07801f
C3033 a_638_3764.n36 VSS 0.2494f
C3034 a_638_3764.t40 VSS 0.07629f
C3035 a_638_3764.n37 VSS 0.20508f
C3036 a_638_3764.t13 VSS 0.07629f
C3037 a_638_3764.n38 VSS 0.20508f
C3038 a_638_3764.t12 VSS 0.07629f
C3039 a_638_3764.n39 VSS 0.20508f
C3040 a_638_3764.t9 VSS 0.07629f
C3041 a_638_3764.n40 VSS 0.20508f
C3042 a_638_3764.t48 VSS 0.07629f
C3043 a_638_3764.n41 VSS 0.20508f
C3044 a_638_3764.t60 VSS 0.07629f
C3045 a_638_3764.n42 VSS 0.20508f
C3046 a_638_3764.t10 VSS 0.07629f
C3047 a_638_3764.n43 VSS 0.2351f
C3048 a_638_3764.t36 VSS 0.07629f
C3049 a_638_3764.n44 VSS 0.2351f
C3050 a_638_3764.t49 VSS 0.07629f
C3051 a_638_3764.n45 VSS 0.20508f
C3052 a_638_3764.t25 VSS 0.07629f
C3053 a_638_3764.n46 VSS 0.20508f
C3054 a_638_3764.t50 VSS 0.07629f
C3055 a_638_3764.n47 VSS 0.20508f
C3056 a_638_3764.t44 VSS 0.07629f
C3057 a_638_3764.n48 VSS 0.20508f
C3058 a_638_3764.t17 VSS 0.07629f
C3059 a_638_3764.n49 VSS 0.20508f
C3060 a_638_3764.t66 VSS 0.07629f
C3061 a_638_3764.n50 VSS 0.20508f
C3062 a_638_3764.t22 VSS 0.07629f
C3063 a_638_3764.n51 VSS 0.2351f
C3064 a_638_3764.t8 VSS 0.07629f
C3065 a_638_3764.n52 VSS 0.2351f
C3066 a_638_3764.t43 VSS 0.07629f
C3067 a_638_3764.n53 VSS 0.20508f
C3068 a_638_3764.t63 VSS 0.07629f
C3069 a_638_3764.n54 VSS 0.20508f
C3070 a_638_3764.t34 VSS 0.07629f
C3071 a_638_3764.n55 VSS 0.20508f
C3072 a_638_3764.t24 VSS 0.07629f
C3073 a_638_3764.n56 VSS 0.20508f
C3074 a_638_3764.t56 VSS 0.07629f
C3075 a_638_3764.n57 VSS 0.20508f
C3076 a_638_3764.t46 VSS 0.07629f
C3077 a_638_3764.n58 VSS 0.20508f
C3078 a_638_3764.t3 VSS 0.07629f
C3079 a_638_3764.n59 VSS 0.2351f
C3080 a_638_3764.t21 VSS 0.07629f
C3081 a_638_3764.n60 VSS 0.2351f
C3082 a_638_3764.t45 VSS 0.07629f
C3083 a_638_3764.n61 VSS 0.20508f
C3084 a_638_3764.t65 VSS 0.07629f
C3085 a_638_3764.n62 VSS 0.20508f
C3086 a_638_3764.t47 VSS 0.07629f
C3087 a_638_3764.n63 VSS 0.20508f
C3088 a_638_3764.t39 VSS 0.07629f
C3089 a_638_3764.n64 VSS 0.20508f
C3090 a_638_3764.t67 VSS 0.07629f
C3091 a_638_3764.n65 VSS 0.20508f
C3092 a_638_3764.t37 VSS 0.07629f
C3093 a_638_3764.n66 VSS 0.20508f
C3094 a_638_3764.t20 VSS 0.07629f
C3095 a_638_3764.n67 VSS 0.19068f
C3096 a_638_3764.t27 VSS 0.07629f
C3097 a_638_3764.t7 VSS 0.21301f
C3098 a_638_3764.t29 VSS 0.21301f
C3099 a_638_3764.n68 VSS 0.42602f
C3100 a_638_3764.n69 VSS -0.52759f
C3101 a_638_3764.n70 VSS 0.15155f
C3102 a_638_3764.n71 VSS 0.13888f
C3103 a_638_3764.t6 VSS 0.50628f
C3104 a_638_3764.n72 VSS 0.82359f
C3105 a_20810_7557.t0 VSS 3.74618f
C3106 a_20810_7557.t1 VSS 2.35382f
C3107 a_7830_25520.t0 VSS 4.30261f
C3108 a_7830_25520.t1 VSS 1.69739f
C3109 BIT_SEL[23].t6 VSS 4.06977f
C3110 BIT_SEL[23].n0 VSS 7.03381f
C3111 BIT_SEL[23].t0 VSS 4.06977f
C3112 BIT_SEL[23].n1 VSS 7.03381f
C3113 BIT_SEL[23].t1 VSS 4.06977f
C3114 BIT_SEL[23].n2 VSS 7.03381f
C3115 BIT_SEL[23].t3 VSS 4.06977f
C3116 BIT_SEL[23].n3 VSS 7.03381f
C3117 BIT_SEL[23].t7 VSS 4.06977f
C3118 BIT_SEL[23].n4 VSS 7.03381f
C3119 BIT_SEL[23].t5 VSS 4.06977f
C3120 BIT_SEL[23].n5 VSS 7.03381f
C3121 BIT_SEL[23].t2 VSS 4.06977f
C3122 BIT_SEL[23].n6 VSS 7.03381f
C3123 BIT_SEL[23].t4 VSS 4.20835f
C3124 a_20810_25152.t0 VSS 1.79192f
C3125 a_20810_25152.t1 VSS 4.20808f
C3126 a_14320_13801.t0 VSS 4.25498f
C3127 a_14320_13801.t1 VSS 1.74502f
C3128 BIT_SEL[38].t5 VSS 4.07324f
C3129 BIT_SEL[38].n0 VSS 7.01202f
C3130 BIT_SEL[38].t0 VSS 4.07324f
C3131 BIT_SEL[38].n1 VSS 7.01202f
C3132 BIT_SEL[38].t2 VSS 4.07324f
C3133 BIT_SEL[38].n2 VSS 7.01202f
C3134 BIT_SEL[38].t6 VSS 4.07324f
C3135 BIT_SEL[38].n3 VSS 7.01202f
C3136 BIT_SEL[38].t7 VSS 4.07324f
C3137 BIT_SEL[38].n4 VSS 7.01202f
C3138 BIT_SEL[38].t1 VSS 4.07324f
C3139 BIT_SEL[38].n5 VSS 7.01202f
C3140 BIT_SEL[38].t3 VSS 4.07324f
C3141 BIT_SEL[38].n6 VSS 7.01202f
C3142 BIT_SEL[38].t4 VSS 4.21129f
C3143 a_20810_52289.t0 VSS 4.30649f
C3144 a_20810_52289.t1 VSS 1.69351f
C3145 a_1340_11031.t0 VSS 4.60993f
C3146 a_1340_11031.t1 VSS 1.39007f
C3147 a_20810_36903.t0 VSS 1.7215f
C3148 a_20810_36903.t1 VSS 4.2785f
C3149 BIT_SEL[52].t6 VSS 4.02347f
C3150 BIT_SEL[52].n0 VSS 6.87043f
C3151 BIT_SEL[52].t4 VSS 4.02347f
C3152 BIT_SEL[52].n1 VSS 6.87043f
C3153 BIT_SEL[52].t2 VSS 4.02347f
C3154 BIT_SEL[52].n2 VSS 6.87043f
C3155 BIT_SEL[52].t5 VSS 4.02347f
C3156 BIT_SEL[52].n3 VSS 6.87043f
C3157 BIT_SEL[52].t0 VSS 4.02347f
C3158 BIT_SEL[52].n4 VSS 6.87043f
C3159 BIT_SEL[52].t7 VSS 4.02347f
C3160 BIT_SEL[52].n5 VSS 6.87043f
C3161 BIT_SEL[52].t1 VSS 4.02347f
C3162 BIT_SEL[52].n6 VSS 6.87043f
C3163 BIT_SEL[52].t3 VSS 4.11755f
C3164 a_7738_43466.t0 VSS 4.52345f
C3165 a_7738_43466.t1 VSS 1.47655f
C3166 a_7830_25152.t0 VSS 4.20807f
C3167 a_7830_25152.t1 VSS 1.79193f
C3168 BIT_SEL[25].t6 VSS 4.14534f
C3169 BIT_SEL[25].n0 VSS 7.22001f
C3170 BIT_SEL[25].t0 VSS 4.14534f
C3171 BIT_SEL[25].n1 VSS 7.22001f
C3172 BIT_SEL[25].t4 VSS 4.14534f
C3173 BIT_SEL[25].n2 VSS 7.22001f
C3174 BIT_SEL[25].t2 VSS 4.14534f
C3175 BIT_SEL[25].n3 VSS 7.22001f
C3176 BIT_SEL[25].t5 VSS 4.14534f
C3177 BIT_SEL[25].n4 VSS 7.22001f
C3178 BIT_SEL[25].t7 VSS 4.14534f
C3179 BIT_SEL[25].n5 VSS 7.22001f
C3180 BIT_SEL[25].t1 VSS 4.14534f
C3181 BIT_SEL[25].n6 VSS 7.22001f
C3182 BIT_SEL[25].t3 VSS 4.32038f
C3183 a_20810_9398.t0 VSS 4.20807f
C3184 a_20810_9398.t1 VSS 1.79193f
C3185 a_638_11641.t0 VSS 0.07629f
C3186 a_638_11641.n0 VSS 0.20508f
C3187 a_638_11641.n1 VSS 0.07801f
C3188 a_638_11641.n2 VSS 0.2494f
C3189 a_638_11641.t29 VSS 0.07629f
C3190 a_638_11641.n3 VSS 0.20508f
C3191 a_638_11641.t25 VSS 0.07629f
C3192 a_638_11641.n4 VSS 0.20508f
C3193 a_638_11641.t50 VSS 0.07629f
C3194 a_638_11641.n5 VSS 0.20508f
C3195 a_638_11641.t13 VSS 0.07629f
C3196 a_638_11641.n6 VSS 0.20508f
C3197 a_638_11641.t37 VSS 0.07629f
C3198 a_638_11641.n7 VSS 0.20508f
C3199 a_638_11641.t16 VSS 0.07629f
C3200 a_638_11641.n8 VSS 0.2351f
C3201 a_638_11641.t52 VSS 0.07629f
C3202 a_638_11641.n9 VSS 0.2351f
C3203 a_638_11641.t64 VSS 0.07629f
C3204 a_638_11641.n10 VSS 0.20508f
C3205 a_638_11641.t56 VSS 0.07629f
C3206 a_638_11641.n11 VSS 0.20508f
C3207 a_638_11641.t35 VSS 0.07629f
C3208 a_638_11641.n12 VSS 0.20508f
C3209 a_638_11641.t28 VSS 0.07629f
C3210 a_638_11641.n13 VSS 0.20508f
C3211 a_638_11641.t24 VSS 0.07629f
C3212 a_638_11641.n14 VSS 0.20508f
C3213 a_638_11641.t33 VSS 0.07629f
C3214 a_638_11641.n15 VSS 0.20508f
C3215 a_638_11641.t22 VSS 0.07629f
C3216 a_638_11641.n16 VSS 0.2351f
C3217 a_638_11641.t57 VSS 0.07629f
C3218 a_638_11641.n17 VSS 0.2351f
C3219 a_638_11641.t10 VSS 0.07629f
C3220 a_638_11641.n18 VSS 0.20508f
C3221 a_638_11641.t27 VSS 0.07629f
C3222 a_638_11641.n19 VSS 0.20508f
C3223 a_638_11641.t11 VSS 0.07629f
C3224 a_638_11641.n20 VSS 0.20508f
C3225 a_638_11641.t7 VSS 0.07629f
C3226 a_638_11641.n21 VSS 0.20508f
C3227 a_638_11641.t2 VSS 0.07629f
C3228 a_638_11641.n22 VSS 0.20508f
C3229 a_638_11641.t44 VSS 0.07629f
C3230 a_638_11641.n23 VSS 0.20508f
C3231 a_638_11641.t54 VSS 0.07629f
C3232 a_638_11641.n24 VSS 0.2351f
C3233 a_638_11641.t59 VSS 0.07629f
C3234 a_638_11641.n25 VSS 0.2351f
C3235 a_638_11641.t18 VSS 0.07629f
C3236 a_638_11641.n26 VSS 0.20508f
C3237 a_638_11641.t12 VSS 0.07629f
C3238 a_638_11641.n27 VSS 0.20508f
C3239 a_638_11641.t17 VSS 0.07629f
C3240 a_638_11641.n28 VSS 0.20508f
C3241 a_638_11641.t51 VSS 0.07629f
C3242 a_638_11641.n29 VSS 0.20508f
C3243 a_638_11641.t66 VSS 0.07629f
C3244 a_638_11641.n30 VSS 0.20508f
C3245 a_638_11641.t48 VSS 0.07629f
C3246 a_638_11641.n31 VSS 0.20508f
C3247 a_638_11641.t8 VSS 0.07629f
C3248 a_638_11641.n32 VSS 0.19068f
C3249 a_638_11641.t41 VSS 0.07629f
C3250 a_638_11641.n33 VSS 0.13888f
C3251 a_638_11641.n34 VSS 0.22837f
C3252 a_638_11641.t26 VSS 0.01725f
C3253 a_638_11641.n35 VSS 0.20832f
C3254 a_638_11641.t1 VSS 0.07629f
C3255 a_638_11641.n36 VSS 0.1989f
C3256 a_638_11641.t42 VSS 0.07629f
C3257 a_638_11641.n37 VSS 0.1989f
C3258 a_638_11641.t23 VSS 0.07629f
C3259 a_638_11641.n38 VSS 0.1989f
C3260 a_638_11641.t63 VSS 0.07629f
C3261 a_638_11641.n39 VSS 0.1989f
C3262 a_638_11641.t65 VSS 0.07629f
C3263 a_638_11641.n40 VSS 0.1989f
C3264 a_638_11641.t53 VSS 0.07629f
C3265 a_638_11641.n41 VSS 0.1989f
C3266 a_638_11641.t55 VSS 0.07629f
C3267 a_638_11641.n42 VSS 0.22891f
C3268 a_638_11641.t30 VSS 0.07629f
C3269 a_638_11641.n43 VSS 0.22891f
C3270 a_638_11641.t40 VSS 0.07629f
C3271 a_638_11641.n44 VSS 0.1989f
C3272 a_638_11641.t19 VSS 0.07629f
C3273 a_638_11641.n45 VSS 0.1989f
C3274 a_638_11641.t36 VSS 0.07629f
C3275 a_638_11641.n46 VSS 0.1989f
C3276 a_638_11641.t9 VSS 0.07629f
C3277 a_638_11641.n47 VSS 0.1989f
C3278 a_638_11641.t5 VSS 0.07629f
C3279 a_638_11641.n48 VSS 0.1989f
C3280 a_638_11641.t4 VSS 0.07629f
C3281 a_638_11641.n49 VSS 0.1989f
C3282 a_638_11641.t46 VSS 0.07629f
C3283 a_638_11641.n50 VSS 0.22891f
C3284 a_638_11641.t14 VSS 0.07629f
C3285 a_638_11641.n51 VSS 0.22891f
C3286 a_638_11641.t39 VSS 0.07629f
C3287 a_638_11641.n52 VSS 0.1989f
C3288 a_638_11641.t3 VSS 0.07629f
C3289 a_638_11641.n53 VSS 0.1989f
C3290 a_638_11641.t58 VSS 0.07629f
C3291 a_638_11641.n54 VSS 0.1989f
C3292 a_638_11641.t60 VSS 0.07629f
C3293 a_638_11641.n55 VSS 0.1989f
C3294 a_638_11641.t45 VSS 0.07629f
C3295 a_638_11641.n56 VSS 0.1989f
C3296 a_638_11641.t43 VSS 0.07629f
C3297 a_638_11641.n57 VSS 0.1989f
C3298 a_638_11641.t6 VSS 0.07629f
C3299 a_638_11641.n58 VSS 0.22891f
C3300 a_638_11641.t31 VSS 0.07629f
C3301 a_638_11641.n59 VSS 0.22891f
C3302 a_638_11641.t47 VSS 0.07629f
C3303 a_638_11641.n60 VSS 0.1989f
C3304 a_638_11641.t38 VSS 0.07629f
C3305 a_638_11641.n61 VSS 0.1989f
C3306 a_638_11641.t32 VSS 0.07629f
C3307 a_638_11641.n62 VSS 0.1989f
C3308 a_638_11641.t62 VSS 0.07629f
C3309 a_638_11641.n63 VSS 0.1989f
C3310 a_638_11641.t15 VSS 0.07629f
C3311 a_638_11641.n64 VSS 0.1989f
C3312 a_638_11641.t61 VSS 0.07629f
C3313 a_638_11641.n65 VSS 0.1989f
C3314 a_638_11641.t49 VSS 0.07629f
C3315 a_638_11641.n66 VSS 0.21781f
C3316 a_638_11641.t34 VSS 0.07629f
C3317 a_638_11641.t67 VSS 0.50628f
C3318 a_638_11641.n67 VSS 0.82359f
C3319 a_638_11641.n68 VSS 0.15155f
C3320 a_638_11641.t68 VSS 0.21301f
C3321 a_638_11641.t21 VSS 0.21301f
C3322 a_638_11641.n69 VSS 0.42602f
C3323 a_638_11641.n70 VSS -0.52759f
C3324 a_638_11641.n71 VSS 0.10989f
C3325 a_638_11641.t20 VSS 0.50628f
C3326 a_638_11641.n72 VSS -0.31292f
C3327 a_1340_9029.t0 VSS 1.98079f
C3328 a_1340_9029.t1 VSS 4.01921f
C3329 BIT_SEL[11].t3 VSS 4.11768f
C3330 BIT_SEL[11].n0 VSS 7.22573f
C3331 BIT_SEL[11].t5 VSS 4.11768f
C3332 BIT_SEL[11].n1 VSS 7.22573f
C3333 BIT_SEL[11].t1 VSS 4.11768f
C3334 BIT_SEL[11].n2 VSS 7.22573f
C3335 BIT_SEL[11].t6 VSS 4.11768f
C3336 BIT_SEL[11].n3 VSS 7.22573f
C3337 BIT_SEL[11].t4 VSS 4.11768f
C3338 BIT_SEL[11].n4 VSS 7.22573f
C3339 BIT_SEL[11].t7 VSS 4.11768f
C3340 BIT_SEL[11].n5 VSS 7.22573f
C3341 BIT_SEL[11].t0 VSS 4.11768f
C3342 BIT_SEL[11].n6 VSS 7.22573f
C3343 BIT_SEL[11].t2 VSS 4.3277f
C3344 a_7738_27712.t0 VSS 4.52345f
C3345 a_7738_27712.t1 VSS 1.47655f
C3346 a_1340_40906.t0 VSS 1.79192f
C3347 a_1340_40906.t1 VSS 4.20808f
C3348 a_638_43149.t0 VSS 0.07629f
C3349 a_638_43149.n0 VSS 0.1989f
C3350 a_638_43149.n1 VSS 0.20832f
C3351 a_638_43149.t6 VSS 0.07629f
C3352 a_638_43149.n2 VSS 0.1989f
C3353 a_638_43149.t20 VSS 0.07629f
C3354 a_638_43149.n3 VSS 0.1989f
C3355 a_638_43149.t10 VSS 0.07629f
C3356 a_638_43149.n4 VSS 0.1989f
C3357 a_638_43149.t60 VSS 0.07629f
C3358 a_638_43149.n5 VSS 0.1989f
C3359 a_638_43149.t9 VSS 0.07629f
C3360 a_638_43149.n6 VSS 0.1989f
C3361 a_638_43149.t26 VSS 0.07629f
C3362 a_638_43149.n7 VSS 0.1989f
C3363 a_638_43149.t54 VSS 0.07629f
C3364 a_638_43149.n8 VSS 0.22891f
C3365 a_638_43149.t1 VSS 0.07629f
C3366 a_638_43149.n9 VSS 0.22891f
C3367 a_638_43149.t59 VSS 0.07629f
C3368 a_638_43149.n10 VSS 0.1989f
C3369 a_638_43149.t62 VSS 0.07629f
C3370 a_638_43149.n11 VSS 0.1989f
C3371 a_638_43149.t66 VSS 0.07629f
C3372 a_638_43149.n12 VSS 0.1989f
C3373 a_638_43149.t63 VSS 0.07629f
C3374 a_638_43149.n13 VSS 0.1989f
C3375 a_638_43149.t18 VSS 0.07629f
C3376 a_638_43149.n14 VSS 0.1989f
C3377 a_638_43149.t65 VSS 0.07629f
C3378 a_638_43149.n15 VSS 0.1989f
C3379 a_638_43149.t38 VSS 0.07629f
C3380 a_638_43149.n16 VSS 0.22891f
C3381 a_638_43149.t15 VSS 0.07629f
C3382 a_638_43149.n17 VSS 0.22891f
C3383 a_638_43149.t67 VSS 0.07629f
C3384 a_638_43149.n18 VSS 0.1989f
C3385 a_638_43149.t61 VSS 0.07629f
C3386 a_638_43149.n19 VSS 0.1989f
C3387 a_638_43149.t53 VSS 0.07629f
C3388 a_638_43149.n20 VSS 0.1989f
C3389 a_638_43149.t22 VSS 0.07629f
C3390 a_638_43149.n21 VSS 0.1989f
C3391 a_638_43149.t45 VSS 0.07629f
C3392 a_638_43149.n22 VSS 0.1989f
C3393 a_638_43149.t46 VSS 0.07629f
C3394 a_638_43149.n23 VSS 0.22891f
C3395 a_638_43149.t19 VSS 0.07629f
C3396 a_638_43149.n24 VSS 0.22891f
C3397 a_638_43149.t34 VSS 0.07629f
C3398 a_638_43149.n25 VSS 0.1989f
C3399 a_638_43149.t56 VSS 0.07629f
C3400 a_638_43149.n26 VSS 0.1989f
C3401 a_638_43149.t44 VSS 0.07629f
C3402 a_638_43149.n27 VSS 0.1989f
C3403 a_638_43149.t23 VSS 0.07629f
C3404 a_638_43149.n28 VSS 0.1989f
C3405 a_638_43149.t21 VSS 0.07629f
C3406 a_638_43149.n29 VSS 0.1989f
C3407 a_638_43149.t36 VSS 0.07629f
C3408 a_638_43149.n30 VSS 0.1989f
C3409 a_638_43149.t57 VSS 0.07629f
C3410 a_638_43149.n31 VSS 0.21781f
C3411 a_638_43149.t47 VSS 0.07629f
C3412 a_638_43149.n32 VSS 0.22837f
C3413 a_638_43149.t30 VSS 0.01725f
C3414 a_638_43149.t28 VSS 0.50628f
C3415 a_638_43149.n33 VSS -0.31292f
C3416 a_638_43149.n34 VSS 0.10989f
C3417 a_638_43149.n35 VSS 0.07801f
C3418 a_638_43149.n36 VSS 0.2494f
C3419 a_638_43149.t4 VSS 0.07629f
C3420 a_638_43149.n37 VSS 0.20508f
C3421 a_638_43149.t51 VSS 0.07629f
C3422 a_638_43149.n38 VSS 0.20508f
C3423 a_638_43149.t39 VSS 0.07629f
C3424 a_638_43149.n39 VSS 0.20508f
C3425 a_638_43149.t14 VSS 0.07629f
C3426 a_638_43149.n40 VSS 0.20508f
C3427 a_638_43149.t5 VSS 0.07629f
C3428 a_638_43149.n41 VSS 0.20508f
C3429 a_638_43149.t50 VSS 0.07629f
C3430 a_638_43149.n42 VSS 0.20508f
C3431 a_638_43149.t12 VSS 0.07629f
C3432 a_638_43149.n43 VSS 0.2351f
C3433 a_638_43149.t13 VSS 0.07629f
C3434 a_638_43149.n44 VSS 0.2351f
C3435 a_638_43149.t16 VSS 0.07629f
C3436 a_638_43149.n45 VSS 0.20508f
C3437 a_638_43149.t49 VSS 0.07629f
C3438 a_638_43149.n46 VSS 0.20508f
C3439 a_638_43149.t40 VSS 0.07629f
C3440 a_638_43149.n47 VSS 0.20508f
C3441 a_638_43149.t3 VSS 0.07629f
C3442 a_638_43149.n48 VSS 0.20508f
C3443 a_638_43149.t31 VSS 0.07629f
C3444 a_638_43149.n49 VSS 0.20508f
C3445 a_638_43149.t27 VSS 0.07629f
C3446 a_638_43149.n50 VSS 0.20508f
C3447 a_638_43149.t41 VSS 0.07629f
C3448 a_638_43149.n51 VSS 0.2351f
C3449 a_638_43149.t11 VSS 0.07629f
C3450 a_638_43149.n52 VSS 0.2351f
C3451 a_638_43149.t52 VSS 0.07629f
C3452 a_638_43149.n53 VSS 0.20508f
C3453 a_638_43149.t55 VSS 0.07629f
C3454 a_638_43149.n54 VSS 0.20508f
C3455 a_638_43149.t8 VSS 0.07629f
C3456 a_638_43149.n55 VSS 0.20508f
C3457 a_638_43149.t43 VSS 0.07629f
C3458 a_638_43149.n56 VSS 0.20508f
C3459 a_638_43149.t29 VSS 0.07629f
C3460 a_638_43149.n57 VSS 0.20508f
C3461 a_638_43149.t25 VSS 0.07629f
C3462 a_638_43149.n58 VSS 0.20508f
C3463 a_638_43149.t48 VSS 0.07629f
C3464 a_638_43149.n59 VSS 0.2351f
C3465 a_638_43149.t64 VSS 0.07629f
C3466 a_638_43149.n60 VSS 0.2351f
C3467 a_638_43149.t7 VSS 0.07629f
C3468 a_638_43149.n61 VSS 0.20508f
C3469 a_638_43149.t42 VSS 0.07629f
C3470 a_638_43149.n62 VSS 0.20508f
C3471 a_638_43149.t2 VSS 0.07629f
C3472 a_638_43149.n63 VSS 0.20508f
C3473 a_638_43149.t33 VSS 0.07629f
C3474 a_638_43149.n64 VSS 0.20508f
C3475 a_638_43149.t17 VSS 0.07629f
C3476 a_638_43149.n65 VSS 0.20508f
C3477 a_638_43149.t37 VSS 0.07629f
C3478 a_638_43149.n66 VSS 0.20508f
C3479 a_638_43149.t58 VSS 0.07629f
C3480 a_638_43149.n67 VSS 0.19068f
C3481 a_638_43149.t68 VSS 0.07629f
C3482 a_638_43149.t24 VSS 0.21301f
C3483 a_638_43149.t35 VSS 0.21301f
C3484 a_638_43149.n68 VSS 0.42602f
C3485 a_638_43149.n69 VSS -0.52759f
C3486 a_638_43149.n70 VSS 0.15155f
C3487 a_638_43149.n71 VSS 0.13888f
C3488 a_638_43149.t32 VSS 0.50628f
C3489 a_638_43149.n72 VSS 0.82359f
C3490 a_14320_41274.t0 VSS 4.30261f
C3491 a_14320_41274.t1 VSS 1.69739f
C3492 BIT_SEL[39].t7 VSS 4.06977f
C3493 BIT_SEL[39].n0 VSS 7.03381f
C3494 BIT_SEL[39].t3 VSS 4.06977f
C3495 BIT_SEL[39].n1 VSS 7.03381f
C3496 BIT_SEL[39].t5 VSS 4.06977f
C3497 BIT_SEL[39].n2 VSS 7.03381f
C3498 BIT_SEL[39].t6 VSS 4.06977f
C3499 BIT_SEL[39].n3 VSS 7.03381f
C3500 BIT_SEL[39].t0 VSS 4.06977f
C3501 BIT_SEL[39].n4 VSS 7.03381f
C3502 BIT_SEL[39].t4 VSS 4.06977f
C3503 BIT_SEL[39].n5 VSS 7.03381f
C3504 BIT_SEL[39].t2 VSS 4.06977f
C3505 BIT_SEL[39].n6 VSS 7.03381f
C3506 BIT_SEL[39].t1 VSS 4.20835f
C3507 a_1340_32660.t0 VSS 1.98079f
C3508 a_1340_32660.t1 VSS 4.01921f
C3509 a_638_35272.t0 VSS 0.07629f
C3510 a_638_35272.n0 VSS 0.22891f
C3511 a_638_35272.n1 VSS 0.20832f
C3512 a_638_35272.t68 VSS 0.07629f
C3513 a_638_35272.n2 VSS 0.1989f
C3514 a_638_35272.t56 VSS 0.07629f
C3515 a_638_35272.n3 VSS 0.1989f
C3516 a_638_35272.t63 VSS 0.07629f
C3517 a_638_35272.n4 VSS 0.1989f
C3518 a_638_35272.t38 VSS 0.07629f
C3519 a_638_35272.n5 VSS 0.1989f
C3520 a_638_35272.t60 VSS 0.07629f
C3521 a_638_35272.n6 VSS 0.1989f
C3522 a_638_35272.t14 VSS 0.07629f
C3523 a_638_35272.n7 VSS 0.1989f
C3524 a_638_35272.t52 VSS 0.07629f
C3525 a_638_35272.n8 VSS 0.22891f
C3526 a_638_35272.t34 VSS 0.07629f
C3527 a_638_35272.n9 VSS 0.22891f
C3528 a_638_35272.t33 VSS 0.07629f
C3529 a_638_35272.n10 VSS 0.1989f
C3530 a_638_35272.t15 VSS 0.07629f
C3531 a_638_35272.n11 VSS 0.1989f
C3532 a_638_35272.t47 VSS 0.07629f
C3533 a_638_35272.n12 VSS 0.1989f
C3534 a_638_35272.t6 VSS 0.07629f
C3535 a_638_35272.n13 VSS 0.1989f
C3536 a_638_35272.t24 VSS 0.07629f
C3537 a_638_35272.n14 VSS 0.1989f
C3538 a_638_35272.t1 VSS 0.07629f
C3539 a_638_35272.n15 VSS 0.1989f
C3540 a_638_35272.t62 VSS 0.07629f
C3541 a_638_35272.n16 VSS 0.22891f
C3542 a_638_35272.t30 VSS 0.07629f
C3543 a_638_35272.n17 VSS 0.1989f
C3544 a_638_35272.t8 VSS 0.07629f
C3545 a_638_35272.n18 VSS 0.1989f
C3546 a_638_35272.t11 VSS 0.07629f
C3547 a_638_35272.n19 VSS 0.1989f
C3548 a_638_35272.t43 VSS 0.07629f
C3549 a_638_35272.n20 VSS 0.1989f
C3550 a_638_35272.t37 VSS 0.07629f
C3551 a_638_35272.n21 VSS 0.1989f
C3552 a_638_35272.t49 VSS 0.07629f
C3553 a_638_35272.n22 VSS 0.1989f
C3554 a_638_35272.t39 VSS 0.07629f
C3555 a_638_35272.n23 VSS 0.22891f
C3556 a_638_35272.t46 VSS 0.07629f
C3557 a_638_35272.n24 VSS 0.22891f
C3558 a_638_35272.t50 VSS 0.07629f
C3559 a_638_35272.n25 VSS 0.1989f
C3560 a_638_35272.t48 VSS 0.07629f
C3561 a_638_35272.n26 VSS 0.1989f
C3562 a_638_35272.t5 VSS 0.07629f
C3563 a_638_35272.n27 VSS 0.1989f
C3564 a_638_35272.t67 VSS 0.07629f
C3565 a_638_35272.n28 VSS 0.1989f
C3566 a_638_35272.t57 VSS 0.07629f
C3567 a_638_35272.n29 VSS 0.1989f
C3568 a_638_35272.t40 VSS 0.07629f
C3569 a_638_35272.n30 VSS 0.1989f
C3570 a_638_35272.t12 VSS 0.07629f
C3571 a_638_35272.n31 VSS 0.21781f
C3572 a_638_35272.t29 VSS 0.07629f
C3573 a_638_35272.n32 VSS 0.22837f
C3574 a_638_35272.t32 VSS 0.01725f
C3575 a_638_35272.t3 VSS 0.50628f
C3576 a_638_35272.n33 VSS -0.31292f
C3577 a_638_35272.n34 VSS 0.10989f
C3578 a_638_35272.n35 VSS 0.07801f
C3579 a_638_35272.n36 VSS 0.2494f
C3580 a_638_35272.t19 VSS 0.07629f
C3581 a_638_35272.n37 VSS 0.20508f
C3582 a_638_35272.t54 VSS 0.07629f
C3583 a_638_35272.n38 VSS 0.20508f
C3584 a_638_35272.t26 VSS 0.07629f
C3585 a_638_35272.n39 VSS 0.20508f
C3586 a_638_35272.t18 VSS 0.07629f
C3587 a_638_35272.n40 VSS 0.20508f
C3588 a_638_35272.t31 VSS 0.07629f
C3589 a_638_35272.n41 VSS 0.20508f
C3590 a_638_35272.t13 VSS 0.07629f
C3591 a_638_35272.n42 VSS 0.20508f
C3592 a_638_35272.t45 VSS 0.07629f
C3593 a_638_35272.n43 VSS 0.2351f
C3594 a_638_35272.t35 VSS 0.07629f
C3595 a_638_35272.n44 VSS 0.2351f
C3596 a_638_35272.t61 VSS 0.07629f
C3597 a_638_35272.n45 VSS 0.20508f
C3598 a_638_35272.t36 VSS 0.07629f
C3599 a_638_35272.n46 VSS 0.20508f
C3600 a_638_35272.t55 VSS 0.07629f
C3601 a_638_35272.n47 VSS 0.20508f
C3602 a_638_35272.t17 VSS 0.07629f
C3603 a_638_35272.n48 VSS 0.20508f
C3604 a_638_35272.t64 VSS 0.07629f
C3605 a_638_35272.n49 VSS 0.20508f
C3606 a_638_35272.t65 VSS 0.07629f
C3607 a_638_35272.n50 VSS 0.20508f
C3608 a_638_35272.t41 VSS 0.07629f
C3609 a_638_35272.n51 VSS 0.2351f
C3610 a_638_35272.t7 VSS 0.07629f
C3611 a_638_35272.n52 VSS 0.2351f
C3612 a_638_35272.t22 VSS 0.07629f
C3613 a_638_35272.n53 VSS 0.20508f
C3614 a_638_35272.t25 VSS 0.07629f
C3615 a_638_35272.n54 VSS 0.20508f
C3616 a_638_35272.t42 VSS 0.07629f
C3617 a_638_35272.n55 VSS 0.20508f
C3618 a_638_35272.t53 VSS 0.07629f
C3619 a_638_35272.n56 VSS 0.20508f
C3620 a_638_35272.t20 VSS 0.07629f
C3621 a_638_35272.n57 VSS 0.20508f
C3622 a_638_35272.t4 VSS 0.07629f
C3623 a_638_35272.n58 VSS 0.20508f
C3624 a_638_35272.t66 VSS 0.07629f
C3625 a_638_35272.n59 VSS 0.2351f
C3626 a_638_35272.t44 VSS 0.07629f
C3627 a_638_35272.n60 VSS 0.2351f
C3628 a_638_35272.t9 VSS 0.07629f
C3629 a_638_35272.n61 VSS 0.20508f
C3630 a_638_35272.t51 VSS 0.07629f
C3631 a_638_35272.n62 VSS 0.20508f
C3632 a_638_35272.t27 VSS 0.07629f
C3633 a_638_35272.n63 VSS 0.20508f
C3634 a_638_35272.t21 VSS 0.07629f
C3635 a_638_35272.n64 VSS 0.20508f
C3636 a_638_35272.t28 VSS 0.07629f
C3637 a_638_35272.n65 VSS 0.20508f
C3638 a_638_35272.t16 VSS 0.07629f
C3639 a_638_35272.n66 VSS 0.20508f
C3640 a_638_35272.t10 VSS 0.07629f
C3641 a_638_35272.n67 VSS 0.19068f
C3642 a_638_35272.t23 VSS 0.07629f
C3643 a_638_35272.t58 VSS 0.21301f
C3644 a_638_35272.t59 VSS 0.21301f
C3645 a_638_35272.n68 VSS 0.42602f
C3646 a_638_35272.n69 VSS -0.52759f
C3647 a_638_35272.n70 VSS 0.15155f
C3648 a_638_35272.n71 VSS 0.13888f
C3649 a_638_35272.t2 VSS 0.50628f
C3650 a_638_35272.n72 VSS 0.82359f
C3651 VDD.n0 VSS 1.13271f
C3652 VDD.n1 VSS 0.72948f
C3653 VDD.n2 VSS 0.72948f
C3654 VDD.n3 VSS 0.72948f
C3655 VDD.n4 VSS 0.72948f
C3656 VDD.n5 VSS 0.69303f
C3657 VDD.n6 VSS 0.76593f
C3658 VDD.n7 VSS 0.72948f
C3659 VDD.n8 VSS 0.72948f
C3660 VDD.n9 VSS 0.72948f
C3661 VDD.n10 VSS 0.03962f
C3662 VDD.n11 VSS 0.06962f
C3663 VDD.n12 VSS 0.06962f
C3664 VDD.n13 VSS 0.07284f
C3665 VDD.t88 VSS 0.27515f
C3666 VDD.t90 VSS 0.27515f
C3667 VDD.n14 VSS 0.5503f
C3668 VDD.n15 VSS 0.06133f
C3669 VDD.n16 VSS 0.06649f
C3670 VDD.n17 VSS 0.06962f
C3671 VDD.n18 VSS 0.06962f
C3672 VDD.n19 VSS 0.06962f
C3673 VDD.n20 VSS 0.08585f
C3674 VDD.n21 VSS 1.4977f
C3675 VDD.n22 VSS 0.03962f
C3676 VDD.n23 VSS 0.06962f
C3677 VDD.n24 VSS 0.06962f
C3678 VDD.n25 VSS 0.07284f
C3679 VDD.t87 VSS 0.27515f
C3680 VDD.t89 VSS 0.27515f
C3681 VDD.n26 VSS 0.5503f
C3682 VDD.n27 VSS 0.06133f
C3683 VDD.n28 VSS 0.06649f
C3684 VDD.n29 VSS 0.06962f
C3685 VDD.n30 VSS 0.06962f
C3686 VDD.n31 VSS 0.06962f
C3687 VDD.n32 VSS 0.08585f
C3688 VDD.n33 VSS 1.13271f
C3689 VDD.n34 VSS 0.72948f
C3690 VDD.n35 VSS 0.72948f
C3691 VDD.n36 VSS 0.72948f
C3692 VDD.n37 VSS 0.72948f
C3693 VDD.n38 VSS 0.69303f
C3694 VDD.n39 VSS 0.76593f
C3695 VDD.n40 VSS 0.72948f
C3696 VDD.n41 VSS 0.72948f
C3697 VDD.n42 VSS 0.72948f
C3698 VDD.n43 VSS 0.03962f
C3699 VDD.n44 VSS 0.06962f
C3700 VDD.n45 VSS 0.06962f
C3701 VDD.n46 VSS 0.07284f
C3702 VDD.t246 VSS 0.27515f
C3703 VDD.t253 VSS 0.27515f
C3704 VDD.n47 VSS 0.5503f
C3705 VDD.n48 VSS 0.06133f
C3706 VDD.n49 VSS 0.06649f
C3707 VDD.n50 VSS 0.06962f
C3708 VDD.n51 VSS 0.06962f
C3709 VDD.n52 VSS 0.06962f
C3710 VDD.n53 VSS 0.08585f
C3711 VDD.n54 VSS 1.13024f
C3712 VDD.n55 VSS 0.03962f
C3713 VDD.n56 VSS 0.06962f
C3714 VDD.n57 VSS 0.06962f
C3715 VDD.n58 VSS 0.07284f
C3716 VDD.t254 VSS 0.27515f
C3717 VDD.t252 VSS 0.27515f
C3718 VDD.n59 VSS 0.5503f
C3719 VDD.n60 VSS 0.06133f
C3720 VDD.n61 VSS 0.06649f
C3721 VDD.n62 VSS 0.06962f
C3722 VDD.n63 VSS 0.06962f
C3723 VDD.n64 VSS 0.06962f
C3724 VDD.n65 VSS 0.08585f
C3725 VDD.n66 VSS 1.13271f
C3726 VDD.n67 VSS 0.72948f
C3727 VDD.n68 VSS 0.72948f
C3728 VDD.n69 VSS 0.72948f
C3729 VDD.n70 VSS 0.72948f
C3730 VDD.n71 VSS 0.69303f
C3731 VDD.n72 VSS 0.76593f
C3732 VDD.n73 VSS 0.72948f
C3733 VDD.n74 VSS 0.72948f
C3734 VDD.n75 VSS 0.72948f
C3735 VDD.n76 VSS 0.03962f
C3736 VDD.n77 VSS 0.06962f
C3737 VDD.n78 VSS 0.06962f
C3738 VDD.n79 VSS 0.07284f
C3739 VDD.t123 VSS 0.27515f
C3740 VDD.t122 VSS 0.27515f
C3741 VDD.n80 VSS 0.5503f
C3742 VDD.n81 VSS 0.06133f
C3743 VDD.n82 VSS 0.06649f
C3744 VDD.n83 VSS 0.06962f
C3745 VDD.n84 VSS 0.06962f
C3746 VDD.n85 VSS 0.06962f
C3747 VDD.n86 VSS 0.08585f
C3748 VDD.n87 VSS 1.13024f
C3749 VDD.n88 VSS 0.03962f
C3750 VDD.n89 VSS 0.06962f
C3751 VDD.n90 VSS 0.06962f
C3752 VDD.n91 VSS 0.07284f
C3753 VDD.t166 VSS 0.27515f
C3754 VDD.t141 VSS 0.27515f
C3755 VDD.n92 VSS 0.5503f
C3756 VDD.n93 VSS 0.06133f
C3757 VDD.n94 VSS 0.06649f
C3758 VDD.n95 VSS 0.06962f
C3759 VDD.n96 VSS 0.06962f
C3760 VDD.n97 VSS 0.06962f
C3761 VDD.n98 VSS 0.08585f
C3762 VDD.n99 VSS 1.13271f
C3763 VDD.n100 VSS 0.72948f
C3764 VDD.n101 VSS 0.72948f
C3765 VDD.n102 VSS 0.72948f
C3766 VDD.n103 VSS 0.72948f
C3767 VDD.n104 VSS 0.69303f
C3768 VDD.n105 VSS 0.76593f
C3769 VDD.n106 VSS 0.72948f
C3770 VDD.n107 VSS 0.72948f
C3771 VDD.n108 VSS 0.72948f
C3772 VDD.n109 VSS 0.03962f
C3773 VDD.n110 VSS 0.06962f
C3774 VDD.n111 VSS 0.06962f
C3775 VDD.n112 VSS 0.07284f
C3776 VDD.t7 VSS 0.27515f
C3777 VDD.t208 VSS 0.27515f
C3778 VDD.n113 VSS 0.5503f
C3779 VDD.n114 VSS 0.06133f
C3780 VDD.n115 VSS 0.06649f
C3781 VDD.n116 VSS 0.06962f
C3782 VDD.n117 VSS 0.06962f
C3783 VDD.n118 VSS 0.06962f
C3784 VDD.n119 VSS 0.08585f
C3785 VDD.n120 VSS 1.13024f
C3786 VDD.n121 VSS 0.03962f
C3787 VDD.n122 VSS 0.06962f
C3788 VDD.n123 VSS 0.06962f
C3789 VDD.n124 VSS 0.07284f
C3790 VDD.t209 VSS 0.27515f
C3791 VDD.t3 VSS 0.27515f
C3792 VDD.n125 VSS 0.5503f
C3793 VDD.n126 VSS 0.06133f
C3794 VDD.n127 VSS 0.06649f
C3795 VDD.n128 VSS 0.06962f
C3796 VDD.n129 VSS 0.06962f
C3797 VDD.n130 VSS 0.06962f
C3798 VDD.n131 VSS 0.08585f
C3799 VDD.n132 VSS 1.13271f
C3800 VDD.n133 VSS 0.72948f
C3801 VDD.n134 VSS 0.72948f
C3802 VDD.n135 VSS 0.72948f
C3803 VDD.n136 VSS 0.72948f
C3804 VDD.n137 VSS 0.69303f
C3805 VDD.n138 VSS 0.76593f
C3806 VDD.n139 VSS 0.72948f
C3807 VDD.n140 VSS 0.72948f
C3808 VDD.n141 VSS 0.72948f
C3809 VDD.n142 VSS 0.03962f
C3810 VDD.n143 VSS 0.06962f
C3811 VDD.n144 VSS 0.06962f
C3812 VDD.n145 VSS 0.07284f
C3813 VDD.t167 VSS 0.27515f
C3814 VDD.t124 VSS 0.27515f
C3815 VDD.n146 VSS 0.5503f
C3816 VDD.n147 VSS 0.06133f
C3817 VDD.n148 VSS 0.06649f
C3818 VDD.n149 VSS 0.06962f
C3819 VDD.n150 VSS 0.06962f
C3820 VDD.n151 VSS 0.06962f
C3821 VDD.n152 VSS 0.08585f
C3822 VDD.n153 VSS 1.13024f
C3823 VDD.n154 VSS 0.03962f
C3824 VDD.n155 VSS 0.06962f
C3825 VDD.n156 VSS 0.06962f
C3826 VDD.n157 VSS 0.07284f
C3827 VDD.t140 VSS 0.27515f
C3828 VDD.t125 VSS 0.27515f
C3829 VDD.n158 VSS 0.5503f
C3830 VDD.n159 VSS 0.06133f
C3831 VDD.n160 VSS 0.06649f
C3832 VDD.n161 VSS 0.06962f
C3833 VDD.n162 VSS 0.06962f
C3834 VDD.n163 VSS 0.06962f
C3835 VDD.n164 VSS 0.08585f
C3836 VDD.n165 VSS 1.13271f
C3837 VDD.n166 VSS 0.72948f
C3838 VDD.n167 VSS 0.72948f
C3839 VDD.n168 VSS 0.72948f
C3840 VDD.n169 VSS 0.72948f
C3841 VDD.n170 VSS 0.69303f
C3842 VDD.n171 VSS 0.76593f
C3843 VDD.n172 VSS 0.72948f
C3844 VDD.n173 VSS 0.72948f
C3845 VDD.n174 VSS 0.72948f
C3846 VDD.n175 VSS 0.03962f
C3847 VDD.n176 VSS 0.06962f
C3848 VDD.n177 VSS 0.06962f
C3849 VDD.n178 VSS 0.07284f
C3850 VDD.t247 VSS 0.27515f
C3851 VDD.t263 VSS 0.27515f
C3852 VDD.n179 VSS 0.5503f
C3853 VDD.n180 VSS 0.06133f
C3854 VDD.n181 VSS 0.06649f
C3855 VDD.n182 VSS 0.06962f
C3856 VDD.n183 VSS 0.06962f
C3857 VDD.n184 VSS 0.06962f
C3858 VDD.n185 VSS 0.08585f
C3859 VDD.n186 VSS 1.13024f
C3860 VDD.n187 VSS 0.03962f
C3861 VDD.n188 VSS 0.06962f
C3862 VDD.n189 VSS 0.06962f
C3863 VDD.n190 VSS 0.07284f
C3864 VDD.t261 VSS 0.27515f
C3865 VDD.t262 VSS 0.27515f
C3866 VDD.n191 VSS 0.5503f
C3867 VDD.n192 VSS 0.06133f
C3868 VDD.n193 VSS 0.06649f
C3869 VDD.n194 VSS 0.06962f
C3870 VDD.n195 VSS 0.06962f
C3871 VDD.n196 VSS 0.06962f
C3872 VDD.n197 VSS 0.08585f
C3873 VDD.n198 VSS 1.13271f
C3874 VDD.n199 VSS 0.72948f
C3875 VDD.n200 VSS 0.72948f
C3876 VDD.n201 VSS 0.72948f
C3877 VDD.n202 VSS 0.72948f
C3878 VDD.n203 VSS 0.69303f
C3879 VDD.n204 VSS 0.76593f
C3880 VDD.n205 VSS 0.72948f
C3881 VDD.n206 VSS 0.72948f
C3882 VDD.n207 VSS 0.72948f
C3883 VDD.n208 VSS 0.03962f
C3884 VDD.n209 VSS 0.06962f
C3885 VDD.n210 VSS 0.06962f
C3886 VDD.n211 VSS 0.07284f
C3887 VDD.t120 VSS 0.27515f
C3888 VDD.t289 VSS 0.27515f
C3889 VDD.n212 VSS 0.5503f
C3890 VDD.n213 VSS 0.06133f
C3891 VDD.n214 VSS 0.06649f
C3892 VDD.n215 VSS 0.06962f
C3893 VDD.n216 VSS 0.06962f
C3894 VDD.n217 VSS 0.06962f
C3895 VDD.n218 VSS 0.08585f
C3896 VDD.n219 VSS 1.13024f
C3897 VDD.n220 VSS 0.03962f
C3898 VDD.n221 VSS 0.06962f
C3899 VDD.n222 VSS 0.06962f
C3900 VDD.n223 VSS 0.07284f
C3901 VDD.t121 VSS 0.27515f
C3902 VDD.t282 VSS 0.27515f
C3903 VDD.n224 VSS 0.5503f
C3904 VDD.n225 VSS 0.06133f
C3905 VDD.n226 VSS 0.06649f
C3906 VDD.n227 VSS 0.06962f
C3907 VDD.n228 VSS 0.06962f
C3908 VDD.n229 VSS 0.06962f
C3909 VDD.n230 VSS 0.08585f
C3910 VDD.n231 VSS 0.94046f
C3911 VDD.n232 VSS 0.72948f
C3912 VDD.n233 VSS 0.72948f
C3913 VDD.n234 VSS 0.72948f
C3914 VDD.n235 VSS 0.72948f
C3915 VDD.n236 VSS 0.69303f
C3916 VDD.n237 VSS 0.76593f
C3917 VDD.n238 VSS 0.72948f
C3918 VDD.n239 VSS 0.72948f
C3919 VDD.n240 VSS 0.72948f
C3920 VDD.n241 VSS 0.03962f
C3921 VDD.n242 VSS 0.06962f
C3922 VDD.n243 VSS 0.06962f
C3923 VDD.n244 VSS 0.07284f
C3924 VDD.t46 VSS 0.27515f
C3925 VDD.t77 VSS 0.27515f
C3926 VDD.n245 VSS 0.5503f
C3927 VDD.n246 VSS 0.06133f
C3928 VDD.n247 VSS 0.06649f
C3929 VDD.n248 VSS 0.06962f
C3930 VDD.n249 VSS 0.06962f
C3931 VDD.n250 VSS 0.06962f
C3932 VDD.n251 VSS 0.08585f
C3933 VDD.n252 VSS 1.13024f
C3934 VDD.n253 VSS 0.03962f
C3935 VDD.n254 VSS 0.06962f
C3936 VDD.n255 VSS 0.06962f
C3937 VDD.n256 VSS 0.07284f
C3938 VDD.t111 VSS 0.27515f
C3939 VDD.t75 VSS 0.27515f
C3940 VDD.n257 VSS 0.5503f
C3941 VDD.n258 VSS 0.06133f
C3942 VDD.n259 VSS 0.06649f
C3943 VDD.n260 VSS 0.06962f
C3944 VDD.n261 VSS 0.06962f
C3945 VDD.n262 VSS 0.06962f
C3946 VDD.n263 VSS 0.08585f
C3947 VDD.n264 VSS 0.01739f
C3948 VDD.n265 VSS 13.9747f
C3949 VDD.n266 VSS 0.01285f
C3950 VDD.n267 VSS 0.22521f
C3951 VDD.n268 VSS 0.08103f
C3952 VDD.n269 VSS 0.08103f
C3953 VDD.n270 VSS 0.07726f
C3954 VDD.n271 VSS 0.0848f
C3955 VDD.n272 VSS 0.08103f
C3956 VDD.n273 VSS 0.2761f
C3957 VDD.n274 VSS 0.01739f
C3958 VDD.n275 VSS -0.39259f
C3959 VDD.n276 VSS 0.01285f
C3960 VDD.n277 VSS 0.22521f
C3961 VDD.n278 VSS 0.08103f
C3962 VDD.n279 VSS 0.08103f
C3963 VDD.n280 VSS 0.07726f
C3964 VDD.n281 VSS 0.0848f
C3965 VDD.n282 VSS 0.08103f
C3966 VDD.n283 VSS 0.2761f
C3967 VDD.n284 VSS 0.01739f
C3968 VDD.n285 VSS -0.39259f
C3969 VDD.n286 VSS 0.01285f
C3970 VDD.n287 VSS 0.22521f
C3971 VDD.n288 VSS 0.08103f
C3972 VDD.n289 VSS 0.08103f
C3973 VDD.n290 VSS 0.07726f
C3974 VDD.n291 VSS 0.0848f
C3975 VDD.n292 VSS 0.08103f
C3976 VDD.n293 VSS 0.2761f
C3977 VDD.n294 VSS 0.01739f
C3978 VDD.n295 VSS -0.39259f
C3979 VDD.n296 VSS 0.01285f
C3980 VDD.n297 VSS 0.22521f
C3981 VDD.n298 VSS 0.08103f
C3982 VDD.n299 VSS 0.08103f
C3983 VDD.n300 VSS 0.07726f
C3984 VDD.n301 VSS 0.0848f
C3985 VDD.n302 VSS 0.08103f
C3986 VDD.n303 VSS 0.2761f
C3987 VDD.n304 VSS 0.01739f
C3988 VDD.n305 VSS -0.39259f
C3989 VDD.n306 VSS 0.01285f
C3990 VDD.n307 VSS 0.22521f
C3991 VDD.n308 VSS 0.08103f
C3992 VDD.n309 VSS 0.08103f
C3993 VDD.n310 VSS 0.07726f
C3994 VDD.n311 VSS 0.0848f
C3995 VDD.n312 VSS 0.08103f
C3996 VDD.n313 VSS 0.2761f
C3997 VDD.n314 VSS 0.01739f
C3998 VDD.n315 VSS -0.39259f
C3999 VDD.n316 VSS 0.01285f
C4000 VDD.n317 VSS 0.22521f
C4001 VDD.n318 VSS 0.08103f
C4002 VDD.n319 VSS 0.08103f
C4003 VDD.n320 VSS 0.07726f
C4004 VDD.n321 VSS 0.0848f
C4005 VDD.n322 VSS 0.08103f
C4006 VDD.n323 VSS 0.2761f
C4007 VDD.n324 VSS 0.01739f
C4008 VDD.n325 VSS -0.39259f
C4009 VDD.n326 VSS 0.01285f
C4010 VDD.n327 VSS 0.22521f
C4011 VDD.n328 VSS 0.08103f
C4012 VDD.n329 VSS 0.08103f
C4013 VDD.n330 VSS 0.07726f
C4014 VDD.n331 VSS 0.0848f
C4015 VDD.n332 VSS 0.08103f
C4016 VDD.n333 VSS 0.2761f
C4017 VDD.n334 VSS 0.01739f
C4018 VDD.n335 VSS -0.39259f
C4019 VDD.t6 VSS 31.3888f
C4020 VDD.t76 VSS 17.787f
C4021 VDD.t86 VSS 17.787f
C4022 VDD.t2 VSS 19.9668f
C4023 VDD.n336 VSS -0.39259f
C4024 VDD.n337 VSS 0.01285f
C4025 VDD.n338 VSS 0.22521f
C4026 VDD.n339 VSS 0.08103f
C4027 VDD.n340 VSS 0.08103f
C4028 VDD.n341 VSS 0.07726f
C4029 VDD.n342 VSS 0.0848f
C4030 VDD.n343 VSS 0.08103f
C4031 VDD.n344 VSS 0.2761f
C4032 a_1340_25152.t0 VSS 4.20807f
C4033 a_1340_25152.t1 VSS 1.79193f
C4034 a_638_27395.t0 VSS 0.07629f
C4035 a_638_27395.n0 VSS 0.20508f
C4036 a_638_27395.n1 VSS 0.07801f
C4037 a_638_27395.n2 VSS 0.2494f
C4038 a_638_27395.t9 VSS 0.07629f
C4039 a_638_27395.n3 VSS 0.20508f
C4040 a_638_27395.t13 VSS 0.07629f
C4041 a_638_27395.n4 VSS 0.20508f
C4042 a_638_27395.t51 VSS 0.07629f
C4043 a_638_27395.n5 VSS 0.20508f
C4044 a_638_27395.t56 VSS 0.07629f
C4045 a_638_27395.n6 VSS 0.20508f
C4046 a_638_27395.t36 VSS 0.07629f
C4047 a_638_27395.n7 VSS 0.20508f
C4048 a_638_27395.t55 VSS 0.07629f
C4049 a_638_27395.n8 VSS 0.20508f
C4050 a_638_27395.t38 VSS 0.07629f
C4051 a_638_27395.n9 VSS 0.2351f
C4052 a_638_27395.t12 VSS 0.07629f
C4053 a_638_27395.n10 VSS 0.2351f
C4054 a_638_27395.t15 VSS 0.07629f
C4055 a_638_27395.n11 VSS 0.20508f
C4056 a_638_27395.t41 VSS 0.07629f
C4057 a_638_27395.n12 VSS 0.20508f
C4058 a_638_27395.t61 VSS 0.07629f
C4059 a_638_27395.n13 VSS 0.20508f
C4060 a_638_27395.t67 VSS 0.07629f
C4061 a_638_27395.n14 VSS 0.20508f
C4062 a_638_27395.t33 VSS 0.07629f
C4063 a_638_27395.n15 VSS 0.20508f
C4064 a_638_27395.t47 VSS 0.07629f
C4065 a_638_27395.n16 VSS 0.20508f
C4066 a_638_27395.t27 VSS 0.07629f
C4067 a_638_27395.n17 VSS 0.2351f
C4068 a_638_27395.t11 VSS 0.07629f
C4069 a_638_27395.n18 VSS 0.2351f
C4070 a_638_27395.t48 VSS 0.07629f
C4071 a_638_27395.n19 VSS 0.20508f
C4072 a_638_27395.t45 VSS 0.07629f
C4073 a_638_27395.n20 VSS 0.20508f
C4074 a_638_27395.t37 VSS 0.07629f
C4075 a_638_27395.n21 VSS 0.20508f
C4076 a_638_27395.t66 VSS 0.07629f
C4077 a_638_27395.n22 VSS 0.20508f
C4078 a_638_27395.t53 VSS 0.07629f
C4079 a_638_27395.n23 VSS 0.20508f
C4080 a_638_27395.t3 VSS 0.07629f
C4081 a_638_27395.n24 VSS 0.2351f
C4082 a_638_27395.t26 VSS 0.07629f
C4083 a_638_27395.n25 VSS 0.2351f
C4084 a_638_27395.t8 VSS 0.07629f
C4085 a_638_27395.n26 VSS 0.20508f
C4086 a_638_27395.t31 VSS 0.07629f
C4087 a_638_27395.n27 VSS 0.20508f
C4088 a_638_27395.t58 VSS 0.07629f
C4089 a_638_27395.n28 VSS 0.20508f
C4090 a_638_27395.t21 VSS 0.07629f
C4091 a_638_27395.n29 VSS 0.20508f
C4092 a_638_27395.t1 VSS 0.07629f
C4093 a_638_27395.n30 VSS 0.20508f
C4094 a_638_27395.t18 VSS 0.07629f
C4095 a_638_27395.n31 VSS 0.20508f
C4096 a_638_27395.t16 VSS 0.07629f
C4097 a_638_27395.n32 VSS 0.19068f
C4098 a_638_27395.t17 VSS 0.07629f
C4099 a_638_27395.n33 VSS 0.13888f
C4100 a_638_27395.n34 VSS 0.22837f
C4101 a_638_27395.t23 VSS 0.01725f
C4102 a_638_27395.n35 VSS 0.20832f
C4103 a_638_27395.t5 VSS 0.07629f
C4104 a_638_27395.n36 VSS 0.1989f
C4105 a_638_27395.t39 VSS 0.07629f
C4106 a_638_27395.n37 VSS 0.1989f
C4107 a_638_27395.t4 VSS 0.07629f
C4108 a_638_27395.n38 VSS 0.1989f
C4109 a_638_27395.t42 VSS 0.07629f
C4110 a_638_27395.n39 VSS 0.1989f
C4111 a_638_27395.t57 VSS 0.07629f
C4112 a_638_27395.n40 VSS 0.1989f
C4113 a_638_27395.t44 VSS 0.07629f
C4114 a_638_27395.n41 VSS 0.1989f
C4115 a_638_27395.t65 VSS 0.07629f
C4116 a_638_27395.n42 VSS 0.22891f
C4117 a_638_27395.t60 VSS 0.07629f
C4118 a_638_27395.n43 VSS 0.22891f
C4119 a_638_27395.t52 VSS 0.07629f
C4120 a_638_27395.n44 VSS 0.1989f
C4121 a_638_27395.t46 VSS 0.07629f
C4122 a_638_27395.n45 VSS 0.1989f
C4123 a_638_27395.t50 VSS 0.07629f
C4124 a_638_27395.n46 VSS 0.1989f
C4125 a_638_27395.t7 VSS 0.07629f
C4126 a_638_27395.n47 VSS 0.1989f
C4127 a_638_27395.t2 VSS 0.07629f
C4128 a_638_27395.n48 VSS 0.1989f
C4129 a_638_27395.t6 VSS 0.07629f
C4130 a_638_27395.n49 VSS 0.1989f
C4131 a_638_27395.t32 VSS 0.07629f
C4132 a_638_27395.n50 VSS 0.22891f
C4133 a_638_27395.t30 VSS 0.07629f
C4134 a_638_27395.n51 VSS 0.22891f
C4135 a_638_27395.t35 VSS 0.07629f
C4136 a_638_27395.n52 VSS 0.1989f
C4137 a_638_27395.t10 VSS 0.07629f
C4138 a_638_27395.n53 VSS 0.1989f
C4139 a_638_27395.t63 VSS 0.07629f
C4140 a_638_27395.n54 VSS 0.1989f
C4141 a_638_27395.t64 VSS 0.07629f
C4142 a_638_27395.n55 VSS 0.1989f
C4143 a_638_27395.t24 VSS 0.07629f
C4144 a_638_27395.n56 VSS 0.1989f
C4145 a_638_27395.t62 VSS 0.07629f
C4146 a_638_27395.n57 VSS 0.1989f
C4147 a_638_27395.t68 VSS 0.07629f
C4148 a_638_27395.n58 VSS 0.22891f
C4149 a_638_27395.t14 VSS 0.07629f
C4150 a_638_27395.n59 VSS 0.22891f
C4151 a_638_27395.t43 VSS 0.07629f
C4152 a_638_27395.n60 VSS 0.1989f
C4153 a_638_27395.t22 VSS 0.07629f
C4154 a_638_27395.n61 VSS 0.1989f
C4155 a_638_27395.t34 VSS 0.07629f
C4156 a_638_27395.n62 VSS 0.1989f
C4157 a_638_27395.t40 VSS 0.07629f
C4158 a_638_27395.n63 VSS 0.1989f
C4159 a_638_27395.t54 VSS 0.07629f
C4160 a_638_27395.n64 VSS 0.1989f
C4161 a_638_27395.t49 VSS 0.07629f
C4162 a_638_27395.n65 VSS 0.1989f
C4163 a_638_27395.t59 VSS 0.07629f
C4164 a_638_27395.n66 VSS 0.21781f
C4165 a_638_27395.t28 VSS 0.07629f
C4166 a_638_27395.t20 VSS 0.50628f
C4167 a_638_27395.n67 VSS 0.82359f
C4168 a_638_27395.n68 VSS 0.15155f
C4169 a_638_27395.t19 VSS 0.21301f
C4170 a_638_27395.t25 VSS 0.21301f
C4171 a_638_27395.n69 VSS 0.42602f
C4172 a_638_27395.n70 VSS -0.52759f
C4173 a_638_27395.n71 VSS 0.10989f
C4174 a_638_27395.t29 VSS 0.50628f
C4175 a_638_27395.n72 VSS -0.31292f
C4176 a_20810_3154.t0 VSS 4.60993f
C4177 a_20810_3154.t1 VSS 1.39007f
C4178 BIT_SEL[49].t5 VSS 4.07792f
C4179 BIT_SEL[49].n0 VSS 6.88058f
C4180 BIT_SEL[49].t7 VSS 4.07792f
C4181 BIT_SEL[49].n1 VSS 6.88058f
C4182 BIT_SEL[49].t1 VSS 4.07792f
C4183 BIT_SEL[49].n2 VSS 6.88058f
C4184 BIT_SEL[49].t4 VSS 4.07792f
C4185 BIT_SEL[49].n3 VSS 6.88058f
C4186 BIT_SEL[49].t2 VSS 4.07792f
C4187 BIT_SEL[49].n4 VSS 6.88058f
C4188 BIT_SEL[49].t6 VSS 4.07792f
C4189 BIT_SEL[49].n5 VSS 6.88058f
C4190 BIT_SEL[49].t3 VSS 4.07792f
C4191 BIT_SEL[49].n6 VSS 6.88058f
C4192 BIT_SEL[49].t0 VSS 4.12246f
C4193 a_20810_20781.t0 VSS 4.30649f
C4194 a_20810_20781.t1 VSS 1.69351f
C4195 BIT_SEL[50].t4 VSS 4.05315f
C4196 BIT_SEL[50].n0 VSS 6.86345f
C4197 BIT_SEL[50].t2 VSS 4.05315f
C4198 BIT_SEL[50].n1 VSS 6.86345f
C4199 BIT_SEL[50].t0 VSS 4.05315f
C4200 BIT_SEL[50].n2 VSS 6.86345f
C4201 BIT_SEL[50].t5 VSS 4.05315f
C4202 BIT_SEL[50].n3 VSS 6.86345f
C4203 BIT_SEL[50].t6 VSS 4.05315f
C4204 BIT_SEL[50].n4 VSS 6.86345f
C4205 BIT_SEL[50].t7 VSS 4.05315f
C4206 BIT_SEL[50].n5 VSS 6.86345f
C4207 BIT_SEL[50].t1 VSS 4.05315f
C4208 BIT_SEL[50].n6 VSS 6.86345f
C4209 BIT_SEL[50].t3 VSS 4.12109f
C4210 a_7830_61063.t0 VSS 4.25498f
C4211 a_7830_61063.t1 VSS 1.74502f
C4212 a_638_58903.t0 VSS 0.07629f
C4213 a_638_58903.n0 VSS 0.1989f
C4214 a_638_58903.n1 VSS 0.20832f
C4215 a_638_58903.t18 VSS 0.07629f
C4216 a_638_58903.n2 VSS 0.1989f
C4217 a_638_58903.t57 VSS 0.07629f
C4218 a_638_58903.n3 VSS 0.1989f
C4219 a_638_58903.t27 VSS 0.07629f
C4220 a_638_58903.n4 VSS 0.1989f
C4221 a_638_58903.t59 VSS 0.07629f
C4222 a_638_58903.n5 VSS 0.1989f
C4223 a_638_58903.t29 VSS 0.07629f
C4224 a_638_58903.n6 VSS 0.1989f
C4225 a_638_58903.t24 VSS 0.07629f
C4226 a_638_58903.n7 VSS 0.1989f
C4227 a_638_58903.t60 VSS 0.07629f
C4228 a_638_58903.n8 VSS 0.22891f
C4229 a_638_58903.t16 VSS 0.07629f
C4230 a_638_58903.n9 VSS 0.22891f
C4231 a_638_58903.t63 VSS 0.07629f
C4232 a_638_58903.n10 VSS 0.1989f
C4233 a_638_58903.t45 VSS 0.07629f
C4234 a_638_58903.n11 VSS 0.1989f
C4235 a_638_58903.t11 VSS 0.07629f
C4236 a_638_58903.n12 VSS 0.1989f
C4237 a_638_58903.t56 VSS 0.07629f
C4238 a_638_58903.n13 VSS 0.1989f
C4239 a_638_58903.t66 VSS 0.07629f
C4240 a_638_58903.n14 VSS 0.1989f
C4241 a_638_58903.t48 VSS 0.07629f
C4242 a_638_58903.n15 VSS 0.22891f
C4243 a_638_58903.t25 VSS 0.07629f
C4244 a_638_58903.n16 VSS 0.22891f
C4245 a_638_58903.t55 VSS 0.07629f
C4246 a_638_58903.n17 VSS 0.1989f
C4247 a_638_58903.t34 VSS 0.07629f
C4248 a_638_58903.n18 VSS 0.1989f
C4249 a_638_58903.t68 VSS 0.07629f
C4250 a_638_58903.n19 VSS 0.1989f
C4251 a_638_58903.t43 VSS 0.07629f
C4252 a_638_58903.n20 VSS 0.1989f
C4253 a_638_58903.t12 VSS 0.07629f
C4254 a_638_58903.n21 VSS 0.1989f
C4255 a_638_58903.t33 VSS 0.07629f
C4256 a_638_58903.n22 VSS 0.1989f
C4257 a_638_58903.t61 VSS 0.07629f
C4258 a_638_58903.n23 VSS 0.22891f
C4259 a_638_58903.t41 VSS 0.07629f
C4260 a_638_58903.n24 VSS 0.22891f
C4261 a_638_58903.t49 VSS 0.07629f
C4262 a_638_58903.n25 VSS 0.1989f
C4263 a_638_58903.t22 VSS 0.07629f
C4264 a_638_58903.n26 VSS 0.1989f
C4265 a_638_58903.t3 VSS 0.07629f
C4266 a_638_58903.n27 VSS 0.1989f
C4267 a_638_58903.t67 VSS 0.07629f
C4268 a_638_58903.n28 VSS 0.1989f
C4269 a_638_58903.t62 VSS 0.07629f
C4270 a_638_58903.n29 VSS 0.1989f
C4271 a_638_58903.t40 VSS 0.07629f
C4272 a_638_58903.n30 VSS 0.1989f
C4273 a_638_58903.t14 VSS 0.07629f
C4274 a_638_58903.n31 VSS 0.21781f
C4275 a_638_58903.t35 VSS 0.07629f
C4276 a_638_58903.n32 VSS 0.22837f
C4277 a_638_58903.t30 VSS 0.01725f
C4278 a_638_58903.t8 VSS 0.50628f
C4279 a_638_58903.n33 VSS -0.31292f
C4280 a_638_58903.n34 VSS 0.10989f
C4281 a_638_58903.n35 VSS 0.07801f
C4282 a_638_58903.n36 VSS 0.2494f
C4283 a_638_58903.t53 VSS 0.07629f
C4284 a_638_58903.n37 VSS 0.20508f
C4285 a_638_58903.t19 VSS 0.07629f
C4286 a_638_58903.n38 VSS 0.20508f
C4287 a_638_58903.t37 VSS 0.07629f
C4288 a_638_58903.n39 VSS 0.20508f
C4289 a_638_58903.t1 VSS 0.07629f
C4290 a_638_58903.n40 VSS 0.20508f
C4291 a_638_58903.t52 VSS 0.07629f
C4292 a_638_58903.n41 VSS 0.20508f
C4293 a_638_58903.t64 VSS 0.07629f
C4294 a_638_58903.n42 VSS 0.20508f
C4295 a_638_58903.t26 VSS 0.07629f
C4296 a_638_58903.n43 VSS 0.2351f
C4297 a_638_58903.t13 VSS 0.07629f
C4298 a_638_58903.n44 VSS 0.2351f
C4299 a_638_58903.t17 VSS 0.07629f
C4300 a_638_58903.n45 VSS 0.20508f
C4301 a_638_58903.t44 VSS 0.07629f
C4302 a_638_58903.n46 VSS 0.20508f
C4303 a_638_58903.t15 VSS 0.07629f
C4304 a_638_58903.n47 VSS 0.20508f
C4305 a_638_58903.t51 VSS 0.07629f
C4306 a_638_58903.n48 VSS 0.20508f
C4307 a_638_58903.t2 VSS 0.07629f
C4308 a_638_58903.n49 VSS 0.20508f
C4309 a_638_58903.t42 VSS 0.07629f
C4310 a_638_58903.n50 VSS 0.20508f
C4311 a_638_58903.t6 VSS 0.07629f
C4312 a_638_58903.n51 VSS 0.2351f
C4313 a_638_58903.t54 VSS 0.07629f
C4314 a_638_58903.n52 VSS 0.2351f
C4315 a_638_58903.t31 VSS 0.07629f
C4316 a_638_58903.n53 VSS 0.20508f
C4317 a_638_58903.t28 VSS 0.07629f
C4318 a_638_58903.n54 VSS 0.20508f
C4319 a_638_58903.t50 VSS 0.07629f
C4320 a_638_58903.n55 VSS 0.20508f
C4321 a_638_58903.t65 VSS 0.07629f
C4322 a_638_58903.n56 VSS 0.20508f
C4323 a_638_58903.t46 VSS 0.07629f
C4324 a_638_58903.n57 VSS 0.20508f
C4325 a_638_58903.t21 VSS 0.07629f
C4326 a_638_58903.n58 VSS 0.20508f
C4327 a_638_58903.t47 VSS 0.07629f
C4328 a_638_58903.n59 VSS 0.2351f
C4329 a_638_58903.t20 VSS 0.07629f
C4330 a_638_58903.n60 VSS 0.2351f
C4331 a_638_58903.t36 VSS 0.07629f
C4332 a_638_58903.n61 VSS 0.20508f
C4333 a_638_58903.t38 VSS 0.07629f
C4334 a_638_58903.n62 VSS 0.20508f
C4335 a_638_58903.t4 VSS 0.07629f
C4336 a_638_58903.n63 VSS 0.20508f
C4337 a_638_58903.t39 VSS 0.07629f
C4338 a_638_58903.n64 VSS 0.20508f
C4339 a_638_58903.t23 VSS 0.07629f
C4340 a_638_58903.n65 VSS 0.20508f
C4341 a_638_58903.t5 VSS 0.07629f
C4342 a_638_58903.n66 VSS 0.20508f
C4343 a_638_58903.t32 VSS 0.07629f
C4344 a_638_58903.n67 VSS 0.19068f
C4345 a_638_58903.t58 VSS 0.07629f
C4346 a_638_58903.t10 VSS 0.21301f
C4347 a_638_58903.t7 VSS 0.21301f
C4348 a_638_58903.n68 VSS 0.42602f
C4349 a_638_58903.n69 VSS -0.52759f
C4350 a_638_58903.n70 VSS 0.15155f
C4351 a_638_58903.n71 VSS 0.13888f
C4352 a_638_58903.t9 VSS 0.50628f
C4353 a_638_58903.n72 VSS 0.82359f
C4354 a_1340_61431.t0 VSS 3.66536f
C4355 a_1340_61431.t1 VSS 2.33464f
.ends

