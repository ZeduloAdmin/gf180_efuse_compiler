* eFuse array netlist with word_width=8, nwords=64
    
.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
X0 ZN I VSS VPW nfet_06v0 W=8.2e-07 L=6e-07  
X1 ZN I VDD VNW pfet_06v0 W=1.22e-06 L=5e-07
.ENDS

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
X00 ZN I VSS VPW nfet_06v0 W=8.2e-07 L=6e-07
X01 VSS I ZN VPW nfet_06v0 W=8.2e-07 L=6e-07
X10 ZN I VDD VNW pfet_06v0 W=1.22e-06 L=5e-07
X11 VDD I ZN VNW pfet_06v0 W=1.22e-06 L=5e-07
.ENDS

.subckt efuse_bitcell VSS VDD SELECT ANODE PARAMS: NUM=-1
X0 ANODE CATHODE efuse NUM={NUM}
X1 CATHODE SELECT VSS VSS nfet_06v0 L=0.60u W=30.5u

.ends

.subckt efuse_senseamp VSS VDD PRESET_N OUT SENSE FUSE
X2 net1 PRESET_N VDD VDD pfet_06v0 L=0.5u W=2.44u nf=2
X1 net2 OUT VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X2 net1 net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X3 net2 net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X1 net1 SENSE FUSE VSS nfet_06v0 L=0.60u W=0.82u
.ends


.subckt efuse_bitline VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63] COL_PROG_N OUT PARAMS: LNUM=0
X0 VSS VDD BIT_SEL[0] bitline efuse_bitcell NUM={LNUM*1000+0}
X1 VSS VDD BIT_SEL[1] bitline efuse_bitcell NUM={LNUM*1000+1}
X2 VSS VDD BIT_SEL[2] bitline efuse_bitcell NUM={LNUM*1000+2}
X3 VSS VDD BIT_SEL[3] bitline efuse_bitcell NUM={LNUM*1000+3}
X4 VSS VDD BIT_SEL[4] bitline efuse_bitcell NUM={LNUM*1000+4}
X5 VSS VDD BIT_SEL[5] bitline efuse_bitcell NUM={LNUM*1000+5}
X6 VSS VDD BIT_SEL[6] bitline efuse_bitcell NUM={LNUM*1000+6}
X7 VSS VDD BIT_SEL[7] bitline efuse_bitcell NUM={LNUM*1000+7}
X8 VSS VDD BIT_SEL[8] bitline efuse_bitcell NUM={LNUM*1000+8}
X9 VSS VDD BIT_SEL[9] bitline efuse_bitcell NUM={LNUM*1000+9}
X10 VSS VDD BIT_SEL[10] bitline efuse_bitcell NUM={LNUM*1000+10}
X11 VSS VDD BIT_SEL[11] bitline efuse_bitcell NUM={LNUM*1000+11}
X12 VSS VDD BIT_SEL[12] bitline efuse_bitcell NUM={LNUM*1000+12}
X13 VSS VDD BIT_SEL[13] bitline efuse_bitcell NUM={LNUM*1000+13}
X14 VSS VDD BIT_SEL[14] bitline efuse_bitcell NUM={LNUM*1000+14}
X15 VSS VDD BIT_SEL[15] bitline efuse_bitcell NUM={LNUM*1000+15}
X16 VSS VDD BIT_SEL[16] bitline efuse_bitcell NUM={LNUM*1000+16}
X17 VSS VDD BIT_SEL[17] bitline efuse_bitcell NUM={LNUM*1000+17}
X18 VSS VDD BIT_SEL[18] bitline efuse_bitcell NUM={LNUM*1000+18}
X19 VSS VDD BIT_SEL[19] bitline efuse_bitcell NUM={LNUM*1000+19}
X20 VSS VDD BIT_SEL[20] bitline efuse_bitcell NUM={LNUM*1000+20}
X21 VSS VDD BIT_SEL[21] bitline efuse_bitcell NUM={LNUM*1000+21}
X22 VSS VDD BIT_SEL[22] bitline efuse_bitcell NUM={LNUM*1000+22}
X23 VSS VDD BIT_SEL[23] bitline efuse_bitcell NUM={LNUM*1000+23}
X24 VSS VDD BIT_SEL[24] bitline efuse_bitcell NUM={LNUM*1000+24}
X25 VSS VDD BIT_SEL[25] bitline efuse_bitcell NUM={LNUM*1000+25}
X26 VSS VDD BIT_SEL[26] bitline efuse_bitcell NUM={LNUM*1000+26}
X27 VSS VDD BIT_SEL[27] bitline efuse_bitcell NUM={LNUM*1000+27}
X28 VSS VDD BIT_SEL[28] bitline efuse_bitcell NUM={LNUM*1000+28}
X29 VSS VDD BIT_SEL[29] bitline efuse_bitcell NUM={LNUM*1000+29}
X30 VSS VDD BIT_SEL[30] bitline efuse_bitcell NUM={LNUM*1000+30}
X31 VSS VDD BIT_SEL[31] bitline efuse_bitcell NUM={LNUM*1000+31}
X32 VSS VDD BIT_SEL[32] bitline efuse_bitcell NUM={LNUM*1000+32}
X33 VSS VDD BIT_SEL[33] bitline efuse_bitcell NUM={LNUM*1000+33}
X34 VSS VDD BIT_SEL[34] bitline efuse_bitcell NUM={LNUM*1000+34}
X35 VSS VDD BIT_SEL[35] bitline efuse_bitcell NUM={LNUM*1000+35}
X36 VSS VDD BIT_SEL[36] bitline efuse_bitcell NUM={LNUM*1000+36}
X37 VSS VDD BIT_SEL[37] bitline efuse_bitcell NUM={LNUM*1000+37}
X38 VSS VDD BIT_SEL[38] bitline efuse_bitcell NUM={LNUM*1000+38}
X39 VSS VDD BIT_SEL[39] bitline efuse_bitcell NUM={LNUM*1000+39}
X40 VSS VDD BIT_SEL[40] bitline efuse_bitcell NUM={LNUM*1000+40}
X41 VSS VDD BIT_SEL[41] bitline efuse_bitcell NUM={LNUM*1000+41}
X42 VSS VDD BIT_SEL[42] bitline efuse_bitcell NUM={LNUM*1000+42}
X43 VSS VDD BIT_SEL[43] bitline efuse_bitcell NUM={LNUM*1000+43}
X44 VSS VDD BIT_SEL[44] bitline efuse_bitcell NUM={LNUM*1000+44}
X45 VSS VDD BIT_SEL[45] bitline efuse_bitcell NUM={LNUM*1000+45}
X46 VSS VDD BIT_SEL[46] bitline efuse_bitcell NUM={LNUM*1000+46}
X47 VSS VDD BIT_SEL[47] bitline efuse_bitcell NUM={LNUM*1000+47}
X48 VSS VDD BIT_SEL[48] bitline efuse_bitcell NUM={LNUM*1000+48}
X49 VSS VDD BIT_SEL[49] bitline efuse_bitcell NUM={LNUM*1000+49}
X50 VSS VDD BIT_SEL[50] bitline efuse_bitcell NUM={LNUM*1000+50}
X51 VSS VDD BIT_SEL[51] bitline efuse_bitcell NUM={LNUM*1000+51}
X52 VSS VDD BIT_SEL[52] bitline efuse_bitcell NUM={LNUM*1000+52}
X53 VSS VDD BIT_SEL[53] bitline efuse_bitcell NUM={LNUM*1000+53}
X54 VSS VDD BIT_SEL[54] bitline efuse_bitcell NUM={LNUM*1000+54}
X55 VSS VDD BIT_SEL[55] bitline efuse_bitcell NUM={LNUM*1000+55}
X56 VSS VDD BIT_SEL[56] bitline efuse_bitcell NUM={LNUM*1000+56}
X57 VSS VDD BIT_SEL[57] bitline efuse_bitcell NUM={LNUM*1000+57}
X58 VSS VDD BIT_SEL[58] bitline efuse_bitcell NUM={LNUM*1000+58}
X59 VSS VDD BIT_SEL[59] bitline efuse_bitcell NUM={LNUM*1000+59}
X60 VSS VDD BIT_SEL[60] bitline efuse_bitcell NUM={LNUM*1000+60}
X61 VSS VDD BIT_SEL[61] bitline efuse_bitcell NUM={LNUM*1000+61}
X62 VSS VDD BIT_SEL[62] bitline efuse_bitcell NUM={LNUM*1000+62}
X63 VSS VDD BIT_SEL[63] bitline efuse_bitcell NUM={LNUM*1000+63}
X0 bitline COL_PROG_N VDD VDD pfet_06v0 L=0.50u W=76.5u nf=2
X1 bitline COL_PROG_N VDD VDD pfet_06v0 L=0.50u W=76.5u nf=2
Xsense VSS VDD PRESET_N OUT SENSE bitline efuse_senseamp
.ends
    

.subckt efuse_array_64x8 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63] COL_PROG_N[0] OUT[0] COL_PROG_N[1] OUT[1] COL_PROG_N[2] OUT[2] COL_PROG_N[3] OUT[3] COL_PROG_N[4] OUT[4] COL_PROG_N[5] OUT[5] COL_PROG_N[6] OUT[6] COL_PROG_N[7] OUT[7]  
X0 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[0] OUT[0]  efuse_bitline LNUM=0
X1 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[1] OUT[1]  efuse_bitline LNUM=1
X2 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[2] OUT[2]  efuse_bitline LNUM=2
X3 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[3] OUT[3]  efuse_bitline LNUM=3
X4 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[4] OUT[4]  efuse_bitline LNUM=4
X5 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[5] OUT[5]  efuse_bitline LNUM=5
X6 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[6] OUT[6]  efuse_bitline LNUM=6
X7 VSS VDD SENSE PRESET_N BIT_SEL[0] BIT_SEL[1] BIT_SEL[2] BIT_SEL[3] BIT_SEL[4] BIT_SEL[5] BIT_SEL[6] BIT_SEL[7] BIT_SEL[8] BIT_SEL[9] BIT_SEL[10] BIT_SEL[11] BIT_SEL[12] BIT_SEL[13] BIT_SEL[14] BIT_SEL[15] BIT_SEL[16] BIT_SEL[17] BIT_SEL[18] BIT_SEL[19] BIT_SEL[20] BIT_SEL[21] BIT_SEL[22] BIT_SEL[23] BIT_SEL[24] BIT_SEL[25] BIT_SEL[26] BIT_SEL[27] BIT_SEL[28] BIT_SEL[29] BIT_SEL[30] BIT_SEL[31] BIT_SEL[32] BIT_SEL[33] BIT_SEL[34] BIT_SEL[35] BIT_SEL[36] BIT_SEL[37] BIT_SEL[38] BIT_SEL[39] BIT_SEL[40] BIT_SEL[41] BIT_SEL[42] BIT_SEL[43] BIT_SEL[44] BIT_SEL[45] BIT_SEL[46] BIT_SEL[47] BIT_SEL[48] BIT_SEL[49] BIT_SEL[50] BIT_SEL[51] BIT_SEL[52] BIT_SEL[53] BIT_SEL[54] BIT_SEL[55] BIT_SEL[56] BIT_SEL[57] BIT_SEL[58] BIT_SEL[59] BIT_SEL[60] BIT_SEL[61] BIT_SEL[62] BIT_SEL[63]  COL_PROG_N[7] OUT[7]  efuse_bitline LNUM=7

.ends
    
.end
    